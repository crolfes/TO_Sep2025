** Cell name: SARADC_FILL1_NOPOWER
.SUBCKT SARADC_FILL1_NOPOWER dummy
.ENDS
