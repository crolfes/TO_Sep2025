module ac_controller_soc_top (clk_pad,
    gpio_1_pad,
    gpio_2_pad,
    pwm_out_pad,
    resetn_pad,
    ser_rx_pad,
    ser_tx_pad,
    spi_flash_clk_pad,
    spi_flash_cs_n_pad,
    spi_flash_io0_pad,
    spi_flash_io1_pad,
    spi_flash_io2_pad,
    spi_flash_io3_pad,
    spi_sensor_clk_pad,
    spi_sensor_cs_n_pad,
    spi_sensor_miso_pad,
    spi_sensor_mosi_pad);
 input clk_pad;
 inout gpio_1_pad;
 inout gpio_2_pad;
 output pwm_out_pad;
 input resetn_pad;
 input ser_rx_pad;
 output ser_tx_pad;
 output spi_flash_clk_pad;
 output spi_flash_cs_n_pad;
 inout spi_flash_io0_pad;
 inout spi_flash_io1_pad;
 inout spi_flash_io2_pad;
 inout spi_flash_io3_pad;
 output spi_sensor_clk_pad;
 output spi_sensor_cs_n_pad;
 input spi_sensor_miso_pad;
 output spi_sensor_mosi_pad;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire clknet_leaf_470_clk;
 wire clknet_leaf_465_clk;
 wire clknet_leaf_463_clk;
 wire clknet_leaf_461_clk;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire clknet_leaf_0_clk;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire net10887;
 wire net10782;
 wire net10871;
 wire net10868;
 wire net11001;
 wire net11010;
 wire net10785;
 wire net10775;
 wire net10960;
 wire net10735;
 wire net10847;
 wire net10770;
 wire net10907;
 wire net10865;
 wire net10961;
 wire net10963;
 wire net10772;
 wire net10771;
 wire net10765;
 wire net10792;
 wire net10905;
 wire net10795;
 wire net10959;
 wire net10967;
 wire net10857;
 wire net10862;
 wire net10766;
 wire net10767;
 wire net10783;
 wire net10794;
 wire net10860;
 wire net10760;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire net10296;
 wire net10291;
 wire _02178_;
 wire _02179_;
 wire net10290;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire clknet_leaf_284_clk;
 wire net10326;
 wire net10286;
 wire clknet_leaf_281_clk;
 wire _02191_;
 wire _02192_;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_278_clk;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire clknet_leaf_285_clk;
 wire net10294;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire net10289;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire net10285;
 wire net10284;
 wire _02218_;
 wire net10282;
 wire _02220_;
 wire _02221_;
 wire net10276;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire clknet_leaf_288_clk;
 wire net10288;
 wire net10287;
 wire net10315;
 wire _02232_;
 wire net10281;
 wire net10275;
 wire _02235_;
 wire net10273;
 wire net10272;
 wire net10267;
 wire net10261;
 wire _02240_;
 wire clknet_leaf_293_clk;
 wire net10274;
 wire _02243_;
 wire net10260;
 wire _02245_;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_289_clk;
 wire _02248_;
 wire net10283;
 wire clknet_leaf_299_clk;
 wire _02251_;
 wire clknet_leaf_295_clk;
 wire net10259;
 wire net10271;
 wire net10270;
 wire _02256_;
 wire net10277;
 wire clknet_leaf_315_clk;
 wire _02259_;
 wire clknet_leaf_304_clk;
 wire net10279;
 wire net10351;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire net10349;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire clknet_leaf_301_clk;
 wire _02279_;
 wire _02280_;
 wire net10258;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire net10269;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire net10265;
 wire clknet_leaf_314_clk;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_311_clk;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire clknet_leaf_308_clk;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire clknet_leaf_306_clk;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire net10266;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire net10332;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire net10346;
 wire net10762;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire net10257;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire net10347;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire net10340;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire net10268;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire net10256;
 wire net10263;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire net10262;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire net10264;
 wire net10327;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire net10429;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire net10253;
 wire _02493_;
 wire net10391;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire net10278;
 wire net10328;
 wire _02508_;
 wire _02509_;
 wire net10251;
 wire net10378;
 wire _02512_;
 wire _02513_;
 wire net10246;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire net10236;
 wire clknet_leaf_318_clk;
 wire _02526_;
 wire _02527_;
 wire net10233;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire clknet_leaf_317_clk;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire net10379;
 wire net10235;
 wire _02583_;
 wire _02584_;
 wire net10393;
 wire net10234;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire net10237;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire clknet_leaf_316_clk;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire net10415;
 wire net10398;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire net10231;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire net10331;
 wire net10341;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire net10353;
 wire net10227;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire net10232;
 wire _02692_;
 wire net10307;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire net10333;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire net10342;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire net10304;
 wire _02777_;
 wire net10390;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire net10255;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire net10218;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire net10226;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire net10239;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire net10215;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire net10198;
 wire net10197;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire net10254;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire net10196;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire net10230;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire net10228;
 wire net10195;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire net10352;
 wire _03278_;
 wire _03279_;
 wire net10428;
 wire net10280;
 wire net10377;
 wire net10224;
 wire net10250;
 wire net10194;
 wire _03286_;
 wire _03287_;
 wire net10238;
 wire clknet_leaf_320_clk;
 wire _03290_;
 wire clknet_leaf_319_clk;
 wire net10221;
 wire _03293_;
 wire net10208;
 wire net10220;
 wire clknet_leaf_321_clk;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire net10201;
 wire net10214;
 wire _03302_;
 wire net10192;
 wire net10213;
 wire _03305_;
 wire _03306_;
 wire net10219;
 wire _03308_;
 wire _03309_;
 wire net10187;
 wire net10193;
 wire _03312_;
 wire net10199;
 wire net10200;
 wire clknet_leaf_322_clk;
 wire net10188;
 wire net10191;
 wire _03318_;
 wire net10242;
 wire net10189;
 wire _03321_;
 wire net10190;
 wire net10183;
 wire net10186;
 wire net10181;
 wire _03326_;
 wire net10180;
 wire net10177;
 wire _03329_;
 wire clknet_leaf_331_clk;
 wire clknet_leaf_330_clk;
 wire _03332_;
 wire clknet_leaf_329_clk;
 wire net10182;
 wire _03335_;
 wire net10175;
 wire net10172;
 wire _03338_;
 wire clknet_leaf_328_clk;
 wire net10185;
 wire _03341_;
 wire net10184;
 wire clknet_leaf_325_clk;
 wire _03344_;
 wire clknet_leaf_323_clk;
 wire net10173;
 wire _03347_;
 wire net10168;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire net10768;
 wire _03354_;
 wire _03355_;
 wire net10179;
 wire net10225;
 wire _03358_;
 wire _03359_;
 wire net10769;
 wire net10249;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire net10339;
 wire net10223;
 wire _03367_;
 wire net10222;
 wire net10241;
 wire _03370_;
 wire net10229;
 wire net10248;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire net10252;
 wire net10247;
 wire net10174;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire net10163;
 wire net10240;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire net10207;
 wire net10209;
 wire _03462_;
 wire net10212;
 wire net10211;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire net10167;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire net10205;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire net10243;
 wire net10216;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire clknet_leaf_334_clk;
 wire net10161;
 wire _03730_;
 wire net10149;
 wire _03732_;
 wire net10150;
 wire net10153;
 wire _03735_;
 wire clknet_leaf_333_clk;
 wire clknet_leaf_332_clk;
 wire net10176;
 wire net10210;
 wire net10178;
 wire clknet_leaf_335_clk;
 wire _03742_;
 wire net10171;
 wire net10162;
 wire _03745_;
 wire _03746_;
 wire net10144;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire net10157;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire net10202;
 wire net10146;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire net10170;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire net10206;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire net10145;
 wire _03812_;
 wire clknet_leaf_337_clk;
 wire clknet_leaf_336_clk;
 wire net10137;
 wire _03816_;
 wire net10136;
 wire net10135;
 wire _03819_;
 wire net10421;
 wire _03821_;
 wire _03822_;
 wire net10165;
 wire net10152;
 wire net10134;
 wire _03826_;
 wire net10151;
 wire net10169;
 wire _03829_;
 wire _03830_;
 wire clknet_leaf_340_clk;
 wire clknet_leaf_338_clk;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire net10133;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire net10132;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire net10148;
 wire net10131;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire net10138;
 wire net10155;
 wire net10154;
 wire net10156;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire net10130;
 wire clknet_leaf_342_clk;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire clknet_leaf_341_clk;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire net10139;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire net10147;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire net10128;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire net10126;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire net10143;
 wire net10142;
 wire net10141;
 wire _04046_;
 wire net10127;
 wire net10140;
 wire _04049_;
 wire clknet_leaf_344_clk;
 wire _04051_;
 wire clknet_leaf_343_clk;
 wire _04053_;
 wire net10118;
 wire _04055_;
 wire net10119;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire net10117;
 wire _04061_;
 wire net10125;
 wire _04063_;
 wire net10121;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire net10124;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire net10120;
 wire net10122;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire net10123;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire net10116;
 wire _04094_;
 wire net10109;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire net10164;
 wire net10114;
 wire _04107_;
 wire net10113;
 wire net10112;
 wire _04110_;
 wire _04111_;
 wire net10108;
 wire _04113_;
 wire _04114_;
 wire net10110;
 wire net10107;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire net10115;
 wire clknet_leaf_346_clk;
 wire _04124_;
 wire net10104;
 wire net10106;
 wire _04127_;
 wire net10105;
 wire net10103;
 wire _04130_;
 wire net10099;
 wire net10098;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire net10101;
 wire net10100;
 wire _04138_;
 wire net10102;
 wire clknet_leaf_348_clk;
 wire _04141_;
 wire _04142_;
 wire net10203;
 wire net10093;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire net10096;
 wire net10095;
 wire _04150_;
 wire net10088;
 wire _04152_;
 wire net10092;
 wire net10091;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire net10204;
 wire net10094;
 wire _04162_;
 wire _04163_;
 wire net10082;
 wire net10158;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire net10244;
 wire net10080;
 wire _04171_;
 wire net10087;
 wire net10081;
 wire _04174_;
 wire net10086;
 wire net10079;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire net10085;
 wire net10083;
 wire _04225_;
 wire net10071;
 wire _04227_;
 wire net10077;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire net10166;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire net10076;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire net10070;
 wire _04251_;
 wire net10073;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire net10072;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire net10074;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire net10075;
 wire net10069;
 wire net10063;
 wire net10065;
 wire net10061;
 wire net10962;
 wire _04302_;
 wire net10068;
 wire _04304_;
 wire _04305_;
 wire net10798;
 wire net10062;
 wire net10064;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire net10067;
 wire _04321_;
 wire net10060;
 wire _04323_;
 wire net10066;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire clknet_leaf_349_clk;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire net10053;
 wire net10089;
 wire _04334_;
 wire net10052;
 wire net10059;
 wire _04337_;
 wire net10058;
 wire net10056;
 wire _04340_;
 wire _04341_;
 wire net10051;
 wire net10055;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire net10054;
 wire net10057;
 wire _04349_;
 wire net10048;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire net10050;
 wire net10880;
 wire _04356_;
 wire net10045;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire net10049;
 wire net10043;
 wire _04367_;
 wire _04368_;
 wire net10042;
 wire _04370_;
 wire net10044;
 wire net10046;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire net10047;
 wire net10037;
 wire _04379_;
 wire net10041;
 wire net10035;
 wire _04382_;
 wire net10034;
 wire net10090;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire net10036;
 wire net10028;
 wire _04390_;
 wire net10040;
 wire net10039;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire net10078;
 wire net10031;
 wire _04401_;
 wire net10016;
 wire net10021;
 wire _04404_;
 wire clknet_leaf_352_clk;
 wire clknet_leaf_350_clk;
 wire _04407_;
 wire _04408_;
 wire net10024;
 wire net10004;
 wire _04411_;
 wire net10038;
 wire net10015;
 wire _04414_;
 wire clknet_leaf_355_clk;
 wire clknet_leaf_353_clk;
 wire _04417_;
 wire _04418_;
 wire net9997;
 wire net10013;
 wire _04421_;
 wire _04422_;
 wire net10008;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire net10014;
 wire clknet_leaf_356_clk;
 wire _04432_;
 wire net10006;
 wire net9990;
 wire _04435_;
 wire net9998;
 wire net10005;
 wire _04438_;
 wire clknet_leaf_365_clk;
 wire net9995;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire net9996;
 wire _04445_;
 wire net9989;
 wire net9987;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire clknet_leaf_362_clk;
 wire clknet_leaf_360_clk;
 wire _04453_;
 wire clknet_leaf_357_clk;
 wire clknet_leaf_359_clk;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire clknet_leaf_358_clk;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire clknet_leaf_366_clk;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire net9992;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire net10029;
 wire _04527_;
 wire net9991;
 wire net9986;
 wire net10027;
 wire _04531_;
 wire net10012;
 wire net10030;
 wire _04534_;
 wire _04535_;
 wire net10020;
 wire _04537_;
 wire net9988;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire clknet_leaf_367_clk;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire net10007;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire net9994;
 wire _04556_;
 wire net9983;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire net10018;
 wire _04565_;
 wire _04566_;
 wire net10019;
 wire _04568_;
 wire net9982;
 wire _04570_;
 wire net10017;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire net9985;
 wire _04583_;
 wire net9984;
 wire _04585_;
 wire _04586_;
 wire clknet_leaf_369_clk;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire clknet_leaf_368_clk;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire net9980;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire net10032;
 wire net9978;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire net10010;
 wire _04614_;
 wire net10009;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire net9993;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire net9979;
 wire _04639_;
 wire net10011;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire net9981;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire clknet_leaf_371_clk;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire clknet_leaf_370_clk;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire net9974;
 wire net10084;
 wire net9999;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire net9977;
 wire net10003;
 wire net9976;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire net10000;
 wire _04720_;
 wire net9975;
 wire _04722_;
 wire net10002;
 wire _04724_;
 wire clknet_leaf_372_clk;
 wire net9968;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire net9969;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire net9967;
 wire net9971;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire net9973;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire net9972;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire net9965;
 wire _04806_;
 wire _04807_;
 wire net9970;
 wire _04809_;
 wire net9966;
 wire _04811_;
 wire clknet_leaf_374_clk;
 wire _04813_;
 wire net9957;
 wire net10026;
 wire net9955;
 wire _04817_;
 wire net9963;
 wire _04819_;
 wire _04820_;
 wire net9962;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire net9959;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire net9961;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire net9956;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire net9958;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire net9960;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire clknet_leaf_375_clk;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire net9951;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire net9950;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire net10023;
 wire net9947;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire net9946;
 wire _04926_;
 wire net9953;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire net10217;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire net9945;
 wire net9949;
 wire net9948;
 wire _04959_;
 wire net9940;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire net9939;
 wire _04966_;
 wire _04967_;
 wire net10033;
 wire _04969_;
 wire net9944;
 wire _04971_;
 wire net9952;
 wire net9964;
 wire _04974_;
 wire net9942;
 wire net9954;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire net9943;
 wire _04981_;
 wire net9941;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire clknet_leaf_376_clk;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire net9927;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire net9926;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire net9938;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire net9933;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire net9929;
 wire _05013_;
 wire net9932;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire net9928;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire net9930;
 wire _05023_;
 wire net9931;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire clknet_leaf_377_clk;
 wire _05029_;
 wire net9924;
 wire net9918;
 wire net9922;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire net9921;
 wire _05037_;
 wire net9937;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire net9917;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire net9916;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire net9923;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire net9919;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire net9913;
 wire _05068_;
 wire net9907;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire net10888;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire net9915;
 wire _05078_;
 wire net9911;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire net9909;
 wire _05084_;
 wire net9912;
 wire net9914;
 wire net9908;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire net9910;
 wire _05092_;
 wire net9906;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire net9920;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire net9903;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire net9901;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire net9905;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire net9900;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire net9898;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire net9899;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire net9902;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire net9904;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire clknet_leaf_378_clk;
 wire _05143_;
 wire net9891;
 wire net10946;
 wire net9895;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire net9897;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire net9896;
 wire net9892;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire net9894;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire net9890;
 wire net9889;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire net9893;
 wire clknet_leaf_379_clk;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire net9883;
 wire net9881;
 wire net10939;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire net9886;
 wire net9925;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire net9885;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire net9884;
 wire net9888;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire net9887;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire net9882;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire net9880;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire net10001;
 wire net9875;
 wire _05429_;
 wire net9872;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire net9879;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire net9877;
 wire net9876;
 wire _05441_;
 wire _05442_;
 wire net9874;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire net9878;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire net9873;
 wire _05459_;
 wire _05460_;
 wire net9936;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire net9869;
 wire _05469_;
 wire _05470_;
 wire net10025;
 wire _05472_;
 wire _05473_;
 wire net9868;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire net9867;
 wire net9864;
 wire _05485_;
 wire net9866;
 wire net9853;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire net10376;
 wire net9861;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire net9858;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire net9844;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire net9850;
 wire net9849;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire net9855;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire net9848;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire net9862;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire net9865;
 wire net9835;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire net9860;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire net9837;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire net9870;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire net9843;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire net9857;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire net9854;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire net9826;
 wire net9859;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire net9836;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire net9829;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire net9828;
 wire net9827;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire net9825;
 wire _05745_;
 wire net9824;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire net9823;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire net9839;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire clknet_leaf_380_clk;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire net9831;
 wire net9814;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire net9820;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire net9817;
 wire clknet_leaf_391_clk;
 wire clknet_leaf_389_clk;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire clknet_leaf_386_clk;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire net9830;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire net9806;
 wire clknet_leaf_385_clk;
 wire _05836_;
 wire net9813;
 wire clknet_leaf_384_clk;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire clknet_leaf_382_clk;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire net9812;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire clknet_leaf_388_clk;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire clknet_leaf_387_clk;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire clknet_leaf_394_clk;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire clknet_leaf_393_clk;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire net9822;
 wire net9808;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire net9809;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire net10940;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire net9821;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire net9863;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire net9818;
 wire _05968_;
 wire net9805;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire net9807;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire clknet_leaf_395_clk;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire net9816;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire net9802;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire net9819;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire net9846;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire net9800;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire net9845;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire net9840;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire net9801;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire net9803;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire clknet_leaf_396_clk;
 wire _06093_;
 wire _06094_;
 wire net9815;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire net10329;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire net9799;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire net9841;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire net9842;
 wire net10330;
 wire net9838;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire net9796;
 wire _06149_;
 wire net9795;
 wire _06151_;
 wire _06152_;
 wire net9804;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire net9791;
 wire net9832;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire net9792;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire net9810;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire net9794;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire net9789;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire net9793;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire net9779;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire net9788;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire net9787;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire net9834;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire net9770;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire net9775;
 wire _06300_;
 wire _06301_;
 wire net9777;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire net9778;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire net10736;
 wire _06321_;
 wire net9762;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire net9755;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire net9833;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire net9763;
 wire net9761;
 wire net9754;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire net9753;
 wire _06397_;
 wire _06398_;
 wire net9752;
 wire _06400_;
 wire net9750;
 wire _06402_;
 wire net9756;
 wire _06404_;
 wire _06405_;
 wire net9748;
 wire _06407_;
 wire _06408_;
 wire net9751;
 wire _06410_;
 wire _06411_;
 wire net9747;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire net9785;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire net9784;
 wire _06421_;
 wire net9745;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire net9764;
 wire _06434_;
 wire net9744;
 wire _06436_;
 wire _06437_;
 wire net9746;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire net9743;
 wire _06446_;
 wire net9811;
 wire _06448_;
 wire _06449_;
 wire net9735;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire net9742;
 wire _06457_;
 wire _06458_;
 wire net9741;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire net9739;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire clknet_leaf_397_clk;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire net9737;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire net9736;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire net9734;
 wire _06489_;
 wire net9738;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire net9733;
 wire _06517_;
 wire net9731;
 wire net9730;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire net9732;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire net9726;
 wire _06535_;
 wire _06536_;
 wire net9727;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire net9729;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire net9740;
 wire _06556_;
 wire _06557_;
 wire clknet_leaf_398_clk;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire net9721;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire net9728;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire net9769;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire net9724;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire net9776;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire net9723;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire net9722;
 wire net9718;
 wire _06637_;
 wire _06638_;
 wire net9871;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire net9717;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire net9720;
 wire net9719;
 wire net9749;
 wire _06669_;
 wire clknet_leaf_399_clk;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire net9712;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire net9715;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire net9714;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire net9711;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire net9716;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire clknet_leaf_400_clk;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire net9700;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire net9710;
 wire _06727_;
 wire net9709;
 wire _06729_;
 wire _06730_;
 wire net9713;
 wire _06732_;
 wire net9780;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire net9702;
 wire _06739_;
 wire clknet_leaf_401_clk;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire net9701;
 wire _06745_;
 wire net9706;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire net9693;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire net9705;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire net9699;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire net9704;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire net9697;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire net9698;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire net9707;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire clknet_leaf_410_clk;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire net9786;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire net9684;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire net9696;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire net9695;
 wire clknet_leaf_409_clk;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire clknet_leaf_408_clk;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire clknet_leaf_407_clk;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire net9694;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire clknet_leaf_406_clk;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire clknet_leaf_404_clk;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire clknet_leaf_403_clk;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire net9683;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire net10945;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire net10896;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire net10882;
 wire _07056_;
 wire clknet_leaf_411_clk;
 wire _07058_;
 wire net9692;
 wire _07060_;
 wire _07061_;
 wire net9774;
 wire _07063_;
 wire _07064_;
 wire net9685;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire net9690;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire net9687;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire net9689;
 wire net9783;
 wire _07148_;
 wire net9782;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire net10881;
 wire net10732;
 wire net9772;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire net9773;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire net9680;
 wire _07171_;
 wire net9765;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire net9790;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire net9681;
 wire net9768;
 wire net9676;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire net9767;
 wire net9766;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire net9781;
 wire _07223_;
 wire _07224_;
 wire net9677;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire net9672;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire net9675;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire net9674;
 wire net9686;
 wire _07260_;
 wire _07261_;
 wire net9682;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire net9671;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire net9669;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire net9663;
 wire _07342_;
 wire _07343_;
 wire net9654;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire clknet_leaf_412_clk;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire net9655;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire net9653;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire net9657;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire net9656;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire clknet_leaf_416_clk;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire clknet_leaf_414_clk;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire net9652;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire net9651;
 wire _07540_;
 wire net9650;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire net9649;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire clknet_leaf_832_clk;
 wire _07697_;
 wire clknet_leaf_831_clk;
 wire _07699_;
 wire clknet_leaf_829_clk;
 wire _07701_;
 wire clknet_leaf_828_clk;
 wire clknet_leaf_824_clk;
 wire clknet_leaf_823_clk;
 wire _07705_;
 wire clknet_leaf_821_clk;
 wire _07707_;
 wire clknet_leaf_820_clk;
 wire clknet_leaf_817_clk;
 wire _07710_;
 wire clknet_leaf_816_clk;
 wire clknet_leaf_815_clk;
 wire clknet_leaf_814_clk;
 wire _07714_;
 wire clknet_leaf_813_clk;
 wire clknet_leaf_811_clk;
 wire clknet_leaf_810_clk;
 wire _07718_;
 wire clknet_leaf_808_clk;
 wire _07720_;
 wire clknet_leaf_807_clk;
 wire clknet_leaf_806_clk;
 wire clknet_leaf_803_clk;
 wire _07724_;
 wire clknet_leaf_801_clk;
 wire clknet_leaf_800_clk;
 wire _07727_;
 wire clknet_leaf_799_clk;
 wire _07729_;
 wire clknet_leaf_798_clk;
 wire clknet_leaf_797_clk;
 wire _07732_;
 wire _07733_;
 wire clknet_leaf_795_clk;
 wire _07735_;
 wire clknet_leaf_794_clk;
 wire _07737_;
 wire clknet_leaf_793_clk;
 wire _07739_;
 wire clknet_leaf_792_clk;
 wire _07741_;
 wire _07742_;
 wire clknet_leaf_791_clk;
 wire _07744_;
 wire clknet_leaf_790_clk;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire clknet_leaf_789_clk;
 wire clknet_leaf_788_clk;
 wire _07754_;
 wire clknet_leaf_787_clk;
 wire clknet_leaf_786_clk;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire clknet_leaf_781_clk;
 wire clknet_leaf_780_clk;
 wire clknet_leaf_778_clk;
 wire clknet_leaf_777_clk;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire clknet_leaf_776_clk;
 wire _07776_;
 wire _07777_;
 wire clknet_leaf_775_clk;
 wire _07779_;
 wire _07780_;
 wire clknet_leaf_774_clk;
 wire clknet_leaf_773_clk;
 wire clknet_leaf_772_clk;
 wire clknet_leaf_771_clk;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire clknet_leaf_770_clk;
 wire clknet_leaf_769_clk;
 wire clknet_leaf_768_clk;
 wire clknet_leaf_767_clk;
 wire clknet_leaf_765_clk;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire clknet_leaf_759_clk;
 wire clknet_leaf_758_clk;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire clknet_leaf_757_clk;
 wire clknet_leaf_755_clk;
 wire clknet_leaf_754_clk;
 wire clknet_leaf_753_clk;
 wire clknet_leaf_752_clk;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire clknet_leaf_750_clk;
 wire clknet_leaf_749_clk;
 wire _07830_;
 wire clknet_leaf_748_clk;
 wire clknet_leaf_747_clk;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire clknet_leaf_744_clk;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire clknet_leaf_743_clk;
 wire clknet_leaf_742_clk;
 wire clknet_leaf_740_clk;
 wire clknet_leaf_739_clk;
 wire _07846_;
 wire _07847_;
 wire clknet_leaf_738_clk;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire clknet_leaf_736_clk;
 wire clknet_leaf_734_clk;
 wire clknet_leaf_733_clk;
 wire clknet_leaf_731_clk;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire clknet_leaf_730_clk;
 wire _07874_;
 wire clknet_leaf_728_clk;
 wire _07876_;
 wire clknet_leaf_727_clk;
 wire _07878_;
 wire clknet_leaf_726_clk;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire clknet_leaf_725_clk;
 wire _07889_;
 wire _07890_;
 wire clknet_leaf_724_clk;
 wire _07892_;
 wire clknet_leaf_723_clk;
 wire _07894_;
 wire _07895_;
 wire clknet_leaf_722_clk;
 wire _07897_;
 wire clknet_leaf_721_clk;
 wire _07899_;
 wire clknet_leaf_718_clk;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire clknet_leaf_717_clk;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire clknet_leaf_714_clk;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire clknet_leaf_712_clk;
 wire _07926_;
 wire _07927_;
 wire clknet_leaf_711_clk;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire clknet_leaf_708_clk;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire clknet_leaf_707_clk;
 wire _07938_;
 wire clknet_leaf_706_clk;
 wire _07940_;
 wire clknet_leaf_705_clk;
 wire _07942_;
 wire clknet_leaf_704_clk;
 wire clknet_leaf_703_clk;
 wire clknet_leaf_701_clk;
 wire _07946_;
 wire _07947_;
 wire clknet_leaf_700_clk;
 wire _07949_;
 wire clknet_leaf_699_clk;
 wire _07951_;
 wire clknet_leaf_698_clk;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire clknet_leaf_697_clk;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire clknet_leaf_696_clk;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire clknet_leaf_695_clk;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire clknet_leaf_694_clk;
 wire clknet_leaf_693_clk;
 wire _07977_;
 wire clknet_leaf_692_clk;
 wire _07979_;
 wire clknet_leaf_690_clk;
 wire clknet_leaf_689_clk;
 wire _07982_;
 wire clknet_leaf_688_clk;
 wire clknet_leaf_687_clk;
 wire clknet_leaf_685_clk;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire clknet_leaf_684_clk;
 wire _07992_;
 wire clknet_leaf_682_clk;
 wire _07994_;
 wire clknet_leaf_681_clk;
 wire _07996_;
 wire clknet_leaf_680_clk;
 wire _07998_;
 wire clknet_leaf_679_clk;
 wire _08000_;
 wire clknet_leaf_678_clk;
 wire _08002_;
 wire clknet_leaf_677_clk;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire clknet_leaf_676_clk;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire clknet_leaf_672_clk;
 wire _08033_;
 wire clknet_leaf_671_clk;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire clknet_leaf_669_clk;
 wire _08066_;
 wire clknet_leaf_668_clk;
 wire _08068_;
 wire clknet_leaf_667_clk;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire clknet_leaf_666_clk;
 wire clknet_leaf_660_clk;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire clknet_leaf_658_clk;
 wire _08118_;
 wire clknet_leaf_657_clk;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire clknet_leaf_656_clk;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire clknet_leaf_654_clk;
 wire clknet_leaf_653_clk;
 wire clknet_leaf_652_clk;
 wire clknet_leaf_650_clk;
 wire clknet_leaf_648_clk;
 wire clknet_leaf_647_clk;
 wire _08158_;
 wire _08159_;
 wire clknet_leaf_646_clk;
 wire clknet_leaf_645_clk;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire clknet_leaf_644_clk;
 wire clknet_leaf_641_clk;
 wire _08167_;
 wire _08168_;
 wire clknet_leaf_640_clk;
 wire clknet_leaf_636_clk;
 wire _08171_;
 wire clknet_leaf_634_clk;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire clknet_leaf_633_clk;
 wire _08180_;
 wire clknet_leaf_631_clk;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire clknet_leaf_627_clk;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire clknet_leaf_625_clk;
 wire _08199_;
 wire _08200_;
 wire clknet_leaf_624_clk;
 wire clknet_leaf_622_clk;
 wire clknet_leaf_621_clk;
 wire _08204_;
 wire clknet_leaf_620_clk;
 wire _08206_;
 wire _08207_;
 wire clknet_leaf_618_clk;
 wire _08209_;
 wire clknet_leaf_615_clk;
 wire clknet_leaf_613_clk;
 wire _08212_;
 wire _08213_;
 wire clknet_leaf_611_clk;
 wire _08215_;
 wire clknet_leaf_609_clk;
 wire _08217_;
 wire clknet_leaf_608_clk;
 wire clknet_leaf_607_clk;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire clknet_leaf_606_clk;
 wire clknet_leaf_605_clk;
 wire clknet_leaf_604_clk;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire clknet_leaf_603_clk;
 wire clknet_leaf_602_clk;
 wire _08231_;
 wire clknet_leaf_601_clk;
 wire _08233_;
 wire clknet_leaf_599_clk;
 wire clknet_leaf_596_clk;
 wire clknet_leaf_594_clk;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire clknet_leaf_593_clk;
 wire _08243_;
 wire _08244_;
 wire clknet_leaf_592_clk;
 wire _08246_;
 wire clknet_leaf_591_clk;
 wire _08248_;
 wire clknet_leaf_590_clk;
 wire _08250_;
 wire clknet_leaf_587_clk;
 wire _08252_;
 wire clknet_leaf_586_clk;
 wire _08254_;
 wire _08255_;
 wire clknet_leaf_585_clk;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire clknet_leaf_584_clk;
 wire _08261_;
 wire _08262_;
 wire clknet_leaf_583_clk;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire clknet_leaf_582_clk;
 wire clknet_leaf_581_clk;
 wire clknet_leaf_580_clk;
 wire clknet_leaf_579_clk;
 wire _08281_;
 wire clknet_leaf_578_clk;
 wire clknet_leaf_574_clk;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire clknet_leaf_572_clk;
 wire _08289_;
 wire clknet_leaf_571_clk;
 wire clknet_leaf_570_clk;
 wire _08292_;
 wire clknet_leaf_569_clk;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire clknet_leaf_567_clk;
 wire clknet_leaf_566_clk;
 wire clknet_leaf_565_clk;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire clknet_leaf_564_clk;
 wire _08306_;
 wire clknet_leaf_559_clk;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire clknet_leaf_558_clk;
 wire _08312_;
 wire clknet_leaf_557_clk;
 wire _08314_;
 wire clknet_leaf_556_clk;
 wire _08316_;
 wire clknet_leaf_555_clk;
 wire clknet_leaf_554_clk;
 wire clknet_leaf_553_clk;
 wire _08320_;
 wire clknet_leaf_552_clk;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire clknet_leaf_550_clk;
 wire _08328_;
 wire clknet_leaf_547_clk;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire clknet_leaf_546_clk;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire clknet_leaf_543_clk;
 wire clknet_leaf_541_clk;
 wire _08339_;
 wire clknet_leaf_540_clk;
 wire _08341_;
 wire clknet_leaf_539_clk;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire clknet_leaf_538_clk;
 wire clknet_leaf_537_clk;
 wire _08348_;
 wire clknet_leaf_535_clk;
 wire _08350_;
 wire _08351_;
 wire clknet_leaf_534_clk;
 wire _08353_;
 wire clknet_leaf_533_clk;
 wire clknet_leaf_532_clk;
 wire clknet_leaf_530_clk;
 wire clknet_leaf_529_clk;
 wire clknet_leaf_528_clk;
 wire clknet_leaf_526_clk;
 wire clknet_leaf_525_clk;
 wire clknet_leaf_523_clk;
 wire clknet_leaf_519_clk;
 wire _08363_;
 wire clknet_leaf_518_clk;
 wire _08365_;
 wire clknet_leaf_517_clk;
 wire _08367_;
 wire _08368_;
 wire clknet_leaf_513_clk;
 wire _08370_;
 wire clknet_leaf_512_clk;
 wire clknet_leaf_511_clk;
 wire clknet_leaf_509_clk;
 wire _08374_;
 wire _08375_;
 wire clknet_leaf_508_clk;
 wire clknet_leaf_507_clk;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire clknet_leaf_506_clk;
 wire clknet_leaf_505_clk;
 wire clknet_leaf_502_clk;
 wire _08384_;
 wire clknet_leaf_501_clk;
 wire clknet_leaf_498_clk;
 wire _08387_;
 wire clknet_leaf_497_clk;
 wire clknet_leaf_496_clk;
 wire _08390_;
 wire clknet_leaf_495_clk;
 wire clknet_leaf_493_clk;
 wire clknet_leaf_492_clk;
 wire _08394_;
 wire _08395_;
 wire clknet_leaf_491_clk;
 wire _08397_;
 wire clknet_leaf_490_clk;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire clknet_leaf_489_clk;
 wire clknet_leaf_488_clk;
 wire clknet_leaf_487_clk;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire clknet_leaf_486_clk;
 wire _08410_;
 wire clknet_leaf_485_clk;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire clknet_leaf_482_clk;
 wire _08417_;
 wire clknet_leaf_481_clk;
 wire clknet_leaf_478_clk;
 wire _08420_;
 wire clknet_leaf_477_clk;
 wire _08422_;
 wire clknet_leaf_475_clk;
 wire _08424_;
 wire _08425_;
 wire clknet_leaf_474_clk;
 wire _08427_;
 wire _08428_;
 wire clknet_leaf_473_clk;
 wire clknet_leaf_472_clk;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire clknet_leaf_469_clk;
 wire clknet_leaf_467_clk;
 wire _08444_;
 wire clknet_leaf_466_clk;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire clknet_leaf_464_clk;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire clknet_leaf_457_clk;
 wire clknet_leaf_456_clk;
 wire _08463_;
 wire _08464_;
 wire clknet_leaf_455_clk;
 wire clknet_leaf_453_clk;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire clknet_leaf_450_clk;
 wire clknet_leaf_447_clk;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire clknet_leaf_445_clk;
 wire clknet_leaf_444_clk;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire clknet_leaf_442_clk;
 wire clknet_leaf_440_clk;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire clknet_leaf_439_clk;
 wire clknet_leaf_438_clk;
 wire clknet_leaf_437_clk;
 wire _08494_;
 wire _08495_;
 wire clknet_leaf_436_clk;
 wire clknet_leaf_435_clk;
 wire _08498_;
 wire clknet_leaf_434_clk;
 wire _08500_;
 wire clknet_leaf_433_clk;
 wire clknet_leaf_432_clk;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire clknet_leaf_430_clk;
 wire clknet_leaf_429_clk;
 wire _08509_;
 wire _08510_;
 wire clknet_leaf_428_clk;
 wire _08512_;
 wire clknet_leaf_427_clk;
 wire _08514_;
 wire _08515_;
 wire clknet_leaf_426_clk;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire clknet_leaf_425_clk;
 wire clknet_leaf_424_clk;
 wire _08525_;
 wire clknet_leaf_422_clk;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire clknet_leaf_421_clk;
 wire clknet_leaf_420_clk;
 wire _08534_;
 wire clknet_leaf_419_clk;
 wire _08536_;
 wire _08537_;
 wire clknet_leaf_417_clk;
 wire net9645;
 wire _08540_;
 wire net9648;
 wire _08542_;
 wire _08543_;
 wire net9679;
 wire net9646;
 wire _08546_;
 wire net9670;
 wire _08548_;
 wire _08549_;
 wire net9636;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire net10827;
 wire net10845;
 wire net9644;
 wire _08557_;
 wire net9642;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire net9643;
 wire _08566_;
 wire _08567_;
 wire net9641;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire clknet_leaf_45_clk;
 wire net9934;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire net9725;
 wire net11054;
 wire _08584_;
 wire net10944;
 wire _08586_;
 wire net9708;
 wire net9771;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire net9703;
 wire _08593_;
 wire net10937;
 wire net10938;
 wire net10943;
 wire _08597_;
 wire net10936;
 wire net10974;
 wire _08600_;
 wire _08601_;
 wire net10957;
 wire net10891;
 wire net10955;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire net10942;
 wire _08610_;
 wire _08611_;
 wire net10879;
 wire net10966;
 wire _08614_;
 wire _08615_;
 wire net10878;
 wire net10890;
 wire clknet_leaf_130_clk;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire clknet_leaf_124_clk;
 wire _08624_;
 wire net9627;
 wire net9647;
 wire _08627_;
 wire _08628_;
 wire net9678;
 wire net9797;
 wire _08631_;
 wire net10436;
 wire net9798;
 wire _08634_;
 wire net10111;
 wire _08636_;
 wire net10160;
 wire _08638_;
 wire net10129;
 wire net9665;
 wire _08641_;
 wire _08642_;
 wire net9688;
 wire net9667;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire net9666;
 wire _08649_;
 wire net9691;
 wire net9662;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire net9638;
 wire net9658;
 wire net9661;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire net9856;
 wire net10097;
 wire _08664_;
 wire net9639;
 wire net9640;
 wire net10811;
 wire _08668_;
 wire _08669_;
 wire net9847;
 wire net9852;
 wire net9659;
 wire _08673_;
 wire net10022;
 wire net9660;
 wire net9631;
 wire _08677_;
 wire _08678_;
 wire net9851;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire clknet_leaf_123_clk;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire net9629;
 wire net9935;
 wire _08693_;
 wire net9628;
 wire _08695_;
 wire clknet_leaf_122_clk;
 wire _08697_;
 wire _08698_;
 wire net10159;
 wire clknet_leaf_94_clk;
 wire _08701_;
 wire _08702_;
 wire clknet_leaf_87_clk;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire net9630;
 wire clknet_leaf_121_clk;
 wire _08709_;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_116_clk;
 wire _08712_;
 wire net10826;
 wire _08714_;
 wire clknet_leaf_90_clk;
 wire _08716_;
 wire net10245;
 wire net10809;
 wire _08719_;
 wire _08720_;
 wire net10805;
 wire _08722_;
 wire _08723_;
 wire net10808;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_18_clk;
 wire _08727_;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_25_clk;
 wire _08730_;
 wire clknet_leaf_20_clk;
 wire _08732_;
 wire _08733_;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_26_clk;
 wire _08737_;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_14_clk;
 wire _08740_;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_13_clk;
 wire _08743_;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_107_clk;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire clknet_leaf_102_clk;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire clknet_leaf_106_clk;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire clknet_leaf_104_clk;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire clknet_leaf_105_clk;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire clknet_leaf_111_clk;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire clknet_leaf_110_clk;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire clknet_leaf_108_clk;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire clknet_leaf_119_clk;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire clknet_leaf_118_clk;
 wire _08842_;
 wire clknet_leaf_117_clk;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire net10911;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire net10914;
 wire _08861_;
 wire net9673;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire net10908;
 wire clknet_leaf_22_clk;
 wire _08869_;
 wire net10913;
 wire _08871_;
 wire _08872_;
 wire net9635;
 wire net10754;
 wire net10756;
 wire net9664;
 wire net10749;
 wire net9633;
 wire _08879_;
 wire net10411;
 wire _08881_;
 wire net10916;
 wire net9759;
 wire net9757;
 wire _08885_;
 wire _08886_;
 wire net10856;
 wire net10861;
 wire net9760;
 wire _08890_;
 wire net9632;
 wire _08892_;
 wire _08893_;
 wire net10740;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire net9758;
 wire net10829;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire net10828;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire net10844;
 wire _08944_;
 wire _08945_;
 wire net10931;
 wire net10761;
 wire net10869;
 wire net10751;
 wire net10854;
 wire net10855;
 wire clknet_leaf_58_clk;
 wire net10932;
 wire net9668;
 wire _08955_;
 wire net9637;
 wire net9634;
 wire net10930;
 wire net10912;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire net10927;
 wire net10819;
 wire _08966_;
 wire net10764;
 wire _08968_;
 wire _08969_;
 wire net10815;
 wire _08971_;
 wire clknet_leaf_21_clk;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire net10813;
 wire net10817;
 wire _08983_;
 wire net10812;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire net10915;
 wire _08992_;
 wire net10919;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire net10840;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_56_clk;
 wire _09002_;
 wire net10843;
 wire _09004_;
 wire net10810;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire clknet_leaf_50_clk;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire clknet_leaf_55_clk;
 wire net10807;
 wire _09026_;
 wire net10806;
 wire clknet_leaf_101_clk;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire net10929;
 wire clknet_leaf_85_clk;
 wire _09034_;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_69_clk;
 wire net10835;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire net10830;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire net10832;
 wire _09048_;
 wire net10831;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire net10839;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire net10838;
 wire _09059_;
 wire net10842;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire net10837;
 wire _09067_;
 wire net10918;
 wire clknet_leaf_49_clk;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire clknet_leaf_32_clk;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire net10841;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire net10834;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_75_clk;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire net10836;
 wire clknet_leaf_51_clk;
 wire net10833;
 wire _09098_;
 wire _09099_;
 wire clknet_leaf_68_clk;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire net10909;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire net10910;
 wire _09117_;
 wire clknet_leaf_30_clk;
 wire _09119_;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire _09124_;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_28_clk;
 wire net10824;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire net10825;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire clknet_leaf_84_clk;
 wire net10933;
 wire net10818;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire net11032;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire net11020;
 wire _09157_;
 wire _09158_;
 wire net11024;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire net10821;
 wire _09164_;
 wire net10820;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_81_clk;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire net11053;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire clknet_leaf_60_clk;
 wire _09188_;
 wire _09189_;
 wire clknet_leaf_77_clk;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire net10934;
 wire net11030;
 wire _09196_;
 wire net11017;
 wire net11028;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire net11052;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire net10996;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire net11040;
 wire clknet_leaf_47_clk;
 wire net11051;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire net10983;
 wire _09232_;
 wire net10982;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire net10920;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire net10922;
 wire net10975;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire net10993;
 wire _09247_;
 wire net10997;
 wire net10947;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire net11029;
 wire _09256_;
 wire net10994;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire net10949;
 wire _09265_;
 wire net10988;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire net10995;
 wire net10973;
 wire net10948;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire net10816;
 wire net11033;
 wire net10823;
 wire _09300_;
 wire clknet_leaf_2_clk;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire net11019;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire net11018;
 wire _09312_;
 wire net11026;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire net11034;
 wire clknet_leaf_8_clk;
 wire net11031;
 wire clknet_leaf_83_clk;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire net11027;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire net10814;
 wire net11021;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire net11036;
 wire _09340_;
 wire clknet_leaf_82_clk;
 wire _09342_;
 wire net10822;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire net11025;
 wire net11058;
 wire _09349_;
 wire _09350_;
 wire clknet_leaf_7_clk;
 wire net11022;
 wire net11023;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire net11059;
 wire _09362_;
 wire _09363_;
 wire net10924;
 wire net10917;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire net10926;
 wire net11061;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire net11035;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire net10921;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire net10925;
 wire net11060;
 wire _09391_;
 wire clknet_leaf_4_clk;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire clknet_leaf_6_clk;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_136_clk;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire clknet_leaf_62_clk;
 wire _09422_;
 wire net10952;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire net11037;
 wire net10972;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire net10951;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire net10901;
 wire net11043;
 wire _09453_;
 wire net10900;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire net11000;
 wire _09459_;
 wire net11039;
 wire net10971;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire clknet_leaf_134_clk;
 wire net11042;
 wire _09470_;
 wire _09471_;
 wire net10999;
 wire net10998;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire net10895;
 wire net11057;
 wire net10950;
 wire net10899;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire clknet_leaf_42_clk;
 wire net11048;
 wire _09490_;
 wire net11050;
 wire _09492_;
 wire _09493_;
 wire net11055;
 wire clknet_leaf_131_clk;
 wire _09496_;
 wire net11056;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire net11041;
 wire _09502_;
 wire clknet_leaf_48_clk;
 wire _09504_;
 wire net11046;
 wire net11047;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire clknet_leaf_78_clk;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire net11049;
 wire clknet_leaf_72_clk;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire clknet_leaf_43_clk;
 wire net11038;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire net10928;
 wire net10923;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire net11044;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire clknet_leaf_61_clk;
 wire _09552_;
 wire net11045;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire clknet_leaf_65_clk;
 wire _09558_;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_70_clk;
 wire _09561_;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_63_clk;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire clknet_leaf_44_clk;
 wire _09568_;
 wire net10893;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire net11003;
 wire _09576_;
 wire clknet_leaf_73_clk;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire net11014;
 wire net10978;
 wire net11016;
 wire _09586_;
 wire _09587_;
 wire net11013;
 wire net11012;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire net11015;
 wire _09595_;
 wire net10970;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire net10969;
 wire net10958;
 wire net10935;
 wire _09610_;
 wire _09611_;
 wire net10953;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire clknet_leaf_76_clk;
 wire net10968;
 wire _09619_;
 wire net10976;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire net10874;
 wire net10873;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire net10872;
 wire _09635_;
 wire net10906;
 wire net10984;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire net10992;
 wire net10941;
 wire net10889;
 wire net10875;
 wire net10954;
 wire net10987;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire net10991;
 wire _09657_;
 wire net10986;
 wire _09659_;
 wire net10989;
 wire net10853;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire net10979;
 wire net10877;
 wire net10852;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire net10977;
 wire _09684_;
 wire _09685_;
 wire net10848;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire clknet_leaf_57_clk;
 wire net10990;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire net10981;
 wire net10980;
 wire net10867;
 wire _09709_;
 wire _09710_;
 wire net10850;
 wire _09712_;
 wire net10849;
 wire net10985;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire net10793;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire net10791;
 wire net10876;
 wire net10965;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire net10964;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire net10851;
 wire net10956;
 wire net10788;
 wire _09748_;
 wire _09749_;
 wire net10786;
 wire net10790;
 wire _09752_;
 wire net10789;
 wire net10787;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire clknet_leaf_59_clk;
 wire net10776;
 wire net10777;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire net10773;
 wire net10797;
 wire _09778_;
 wire net11009;
 wire net10897;
 wire net10884;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire net10902;
 wire net10866;
 wire _09794_;
 wire _09795_;
 wire net10758;
 wire net10784;
 wire _09798_;
 wire net10883;
 wire net10885;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire net10870;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire net10892;
 wire net10898;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire net10796;
 wire net10803;
 wire _09828_;
 wire net10750;
 wire net10709;
 wire net10698;
 wire net10695;
 wire net10696;
 wire net10846;
 wire _09835_;
 wire _09836_;
 wire net10693;
 wire net10692;
 wire net10691;
 wire net10903;
 wire net10690;
 wire _09842_;
 wire _09843_;
 wire net10904;
 wire _09845_;
 wire net10734;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire net10689;
 wire _09852_;
 wire net10688;
 wire net10741;
 wire net10753;
 wire _09856_;
 wire _09857_;
 wire net10726;
 wire net10755;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire net10694;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire net10699;
 wire net10802;
 wire _09871_;
 wire _09872_;
 wire net10683;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire net10859;
 wire net10682;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire net10681;
 wire net10687;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire net10779;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire net10686;
 wire net10679;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire net10678;
 wire net10778;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire net10677;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire net10781;
 wire net10676;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire net10680;
 wire net10675;
 wire _09922_;
 wire _09923_;
 wire net10742;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire net10685;
 wire net10780;
 wire net10774;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire net10684;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire net11011;
 wire net10894;
 wire _09941_;
 wire net11005;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire net10671;
 wire net10759;
 wire _09950_;
 wire net11002;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire net10670;
 wire net10858;
 wire _09957_;
 wire net10674;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire net10743;
 wire clknet_leaf_140_clk;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire net10673;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire net11008;
 wire net10746;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire net11007;
 wire net11006;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire net10697;
 wire net10886;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire net11004;
 wire net10757;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire net10733;
 wire net10715;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire net10800;
 wire net10668;
 wire net10672;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire net10716;
 wire net10745;
 wire _10026_;
 wire net10718;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire net10700;
 wire net10701;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire net10669;
 wire net10722;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire net10725;
 wire net10721;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire net10667;
 wire net10724;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_143_clk;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire net10702;
 wire net10706;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire net10703;
 wire net10663;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire net10705;
 wire net10704;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire net10707;
 wire net10655;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire net10662;
 wire net10666;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire net10654;
 wire net10653;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire net10650;
 wire net10644;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire net10639;
 wire _10126_;
 wire net10637;
 wire net10627;
 wire net10710;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire net10661;
 wire _10139_;
 wire _10140_;
 wire net10626;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire net10649;
 wire _10151_;
 wire _10152_;
 wire net10625;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire net10660;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire net10657;
 wire _10171_;
 wire net10624;
 wire net10647;
 wire net10623;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire net10622;
 wire _10184_;
 wire _10185_;
 wire net10633;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire net10628;
 wire _10196_;
 wire _10197_;
 wire net10618;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire net10629;
 wire _10213_;
 wire net10615;
 wire net10614;
 wire net10616;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire net10612;
 wire _10226_;
 wire _10227_;
 wire net10611;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire net10610;
 wire _10238_;
 wire _10239_;
 wire net10648;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire net10609;
 wire net10608;
 wire clknet_leaf_145_clk;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire net10652;
 wire _10266_;
 wire _10267_;
 wire net10607;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire net10621;
 wire _10278_;
 wire _10279_;
 wire clknet_leaf_150_clk;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire clknet_leaf_147_clk;
 wire net10606;
 wire net10619;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire clknet_leaf_149_clk;
 wire _10306_;
 wire _10307_;
 wire clknet_leaf_148_clk;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire net10656;
 wire _10318_;
 wire _10319_;
 wire net10643;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire net10651;
 wire net10640;
 wire net10642;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire net10603;
 wire _10348_;
 wire _10349_;
 wire net10636;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire net10632;
 wire _10360_;
 wire _10361_;
 wire net10658;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire net10631;
 wire net10605;
 wire net10596;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire net10595;
 wire _10388_;
 wire _10389_;
 wire net10613;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire net10593;
 wire _10400_;
 wire _10401_;
 wire net10594;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_151_clk;
 wire net10592;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire net10591;
 wire _10428_;
 wire _10429_;
 wire net10641;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire net10589;
 wire _10440_;
 wire _10441_;
 wire net10588;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire clknet_leaf_153_clk;
 wire net10601;
 wire net10586;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire clknet_leaf_154_clk;
 wire _10468_;
 wire _10469_;
 wire net10602;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire net10585;
 wire _10480_;
 wire _10481_;
 wire clknet_leaf_161_clk;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire clknet_leaf_160_clk;
 wire _10496_;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_155_clk;
 wire _10500_;
 wire net10590;
 wire _10502_;
 wire net10583;
 wire _10504_;
 wire clknet_leaf_158_clk;
 wire _10506_;
 wire net10587;
 wire _10508_;
 wire net10604;
 wire _10510_;
 wire net10630;
 wire _10512_;
 wire net10580;
 wire _10514_;
 wire net10579;
 wire net10645;
 wire _10517_;
 wire net10617;
 wire _10519_;
 wire net10620;
 wire net10584;
 wire _10522_;
 wire net10638;
 wire _10524_;
 wire net10635;
 wire _10526_;
 wire net10581;
 wire _10528_;
 wire net10600;
 wire _10530_;
 wire clknet_leaf_163_clk;
 wire _10532_;
 wire clknet_leaf_162_clk;
 wire _10534_;
 wire net10573;
 wire _10536_;
 wire net10574;
 wire net10582;
 wire _10539_;
 wire net10598;
 wire _10541_;
 wire net10570;
 wire net10567;
 wire _10544_;
 wire net10568;
 wire _10546_;
 wire net10569;
 wire _10548_;
 wire net10563;
 wire _10550_;
 wire net10566;
 wire _10552_;
 wire net10564;
 wire _10554_;
 wire net10560;
 wire _10556_;
 wire net10561;
 wire _10558_;
 wire clknet_leaf_164_clk;
 wire _10560_;
 wire net10559;
 wire _10562_;
 wire net10558;
 wire _10564_;
 wire clknet_leaf_170_clk;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire clknet_leaf_166_clk;
 wire net10554;
 wire net10556;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire clknet_leaf_172_clk;
 wire _10581_;
 wire _10582_;
 wire net10553;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire net10557;
 wire _10593_;
 wire _10594_;
 wire net10552;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire net10548;
 wire net10555;
 wire net10549;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire net10551;
 wire _10621_;
 wire _10622_;
 wire net10546;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire clknet_leaf_173_clk;
 wire _10633_;
 wire _10634_;
 wire net10547;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire net10550;
 wire clknet_leaf_174_clk;
 wire net10543;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire net10544;
 wire _10661_;
 wire _10662_;
 wire clknet_leaf_176_clk;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire net10539;
 wire _10673_;
 wire _10674_;
 wire clknet_leaf_177_clk;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire net10535;
 wire net10538;
 wire net10536;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire net10534;
 wire _10701_;
 wire _10702_;
 wire clknet_leaf_179_clk;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire net10533;
 wire _10713_;
 wire _10714_;
 wire net10531;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire clknet_leaf_182_clk;
 wire net10532;
 wire net10530;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire net10545;
 wire _10743_;
 wire _10744_;
 wire net10529;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire net10528;
 wire _10755_;
 wire _10756_;
 wire net10542;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire net10526;
 wire net10524;
 wire net10525;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire net10522;
 wire _10783_;
 wire _10784_;
 wire net10519;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire clknet_leaf_184_clk;
 wire _10795_;
 wire _10796_;
 wire net10518;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire net10523;
 wire net10516;
 wire net10517;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire net10515;
 wire _10823_;
 wire _10824_;
 wire clknet_leaf_186_clk;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire net10514;
 wire _10835_;
 wire _10836_;
 wire clknet_leaf_188_clk;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire net10513;
 wire clknet_leaf_194_clk;
 wire net10512;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire clknet_leaf_195_clk;
 wire _10863_;
 wire _10864_;
 wire net10511;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire clknet_leaf_197_clk;
 wire _10875_;
 wire _10876_;
 wire clknet_leaf_196_clk;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire net10510;
 wire clknet_leaf_198_clk;
 wire net10509;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire clknet_leaf_200_clk;
 wire _10904_;
 wire _10905_;
 wire net10508;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire net10507;
 wire _10916_;
 wire _10917_;
 wire net10506;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire net10505;
 wire _10932_;
 wire net10504;
 wire net10503;
 wire net10502;
 wire _10936_;
 wire net10501;
 wire _10938_;
 wire net10500;
 wire _10940_;
 wire net10499;
 wire _10942_;
 wire net10498;
 wire _10944_;
 wire net10497;
 wire _10946_;
 wire net10496;
 wire _10948_;
 wire clknet_leaf_201_clk;
 wire _10950_;
 wire net10495;
 wire clknet_leaf_203_clk;
 wire _10953_;
 wire net10494;
 wire _10955_;
 wire net10493;
 wire clknet_leaf_204_clk;
 wire _10958_;
 wire net10521;
 wire _10960_;
 wire clknet_leaf_205_clk;
 wire _10962_;
 wire net10491;
 wire _10964_;
 wire net10492;
 wire _10966_;
 wire net10490;
 wire _10968_;
 wire net10541;
 wire _10970_;
 wire net10520;
 wire _10972_;
 wire net10537;
 wire net10485;
 wire _10975_;
 wire clknet_leaf_207_clk;
 wire _10977_;
 wire net10484;
 wire net10483;
 wire _10980_;
 wire net10482;
 wire _10982_;
 wire clknet_leaf_208_clk;
 wire _10984_;
 wire net10487;
 wire _10986_;
 wire net10486;
 wire _10988_;
 wire clknet_leaf_212_clk;
 wire _10990_;
 wire net10479;
 wire _10992_;
 wire net10478;
 wire _10994_;
 wire clknet_leaf_214_clk;
 wire _10996_;
 wire net10477;
 wire _10998_;
 wire net10489;
 wire _11000_;
 wire net10481;
 wire _11002_;
 wire _11003_;
 wire net10480;
 wire net10476;
 wire net10540;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire net10471;
 wire _11016_;
 wire _11017_;
 wire clknet_leaf_221_clk;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire clknet_leaf_220_clk;
 wire _11028_;
 wire _11029_;
 wire clknet_leaf_218_clk;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire clknet_leaf_216_clk;
 wire net10470;
 wire net10562;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire net10576;
 wire _11056_;
 wire _11057_;
 wire net10720;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire clknet_leaf_226_clk;
 wire _11068_;
 wire _11069_;
 wire net10475;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire net10473;
 wire net10527;
 wire net10571;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire net10488;
 wire _11096_;
 wire _11097_;
 wire clknet_leaf_231_clk;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire clknet_leaf_229_clk;
 wire _11108_;
 wire _11109_;
 wire net10468;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire net10634;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_227_clk;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire net10462;
 wire _11136_;
 wire _11137_;
 wire clknet_leaf_233_clk;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire clknet_leaf_232_clk;
 wire _11148_;
 wire _11149_;
 wire net10469;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire net10474;
 wire net10461;
 wire net10467;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire net10565;
 wire _11177_;
 wire _11178_;
 wire net10597;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire net10466;
 wire _11189_;
 wire _11190_;
 wire net10464;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire clknet_leaf_234_clk;
 wire net10460;
 wire net10472;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire net10575;
 wire _11217_;
 wire _11218_;
 wire net10646;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire net10463;
 wire _11229_;
 wire _11230_;
 wire net10465;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_240_clk;
 wire net10457;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire net10665;
 wire _11257_;
 wire _11258_;
 wire net10458;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire net10455;
 wire _11269_;
 wire _11270_;
 wire clknet_leaf_238_clk;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_244_clk;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire net10578;
 wire _11297_;
 wire _11298_;
 wire clknet_leaf_243_clk;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire clknet_leaf_242_clk;
 wire _11309_;
 wire _11310_;
 wire net10577;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire net10572;
 wire net10447;
 wire net10452;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire net10459;
 wire _11337_;
 wire _11338_;
 wire net10453;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire net10456;
 wire _11349_;
 wire _11350_;
 wire net10719;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire net10664;
 wire net10445;
 wire net10744;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire net10450;
 wire _11377_;
 wire _11378_;
 wire net10763;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire net10446;
 wire _11389_;
 wire _11390_;
 wire net10717;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire net10712;
 wire _11407_;
 wire _11408_;
 wire net10441;
 wire _11410_;
 wire _11411_;
 wire net10711;
 wire _11413_;
 wire net10748;
 wire net10752;
 wire _11416_;
 wire net10440;
 wire _11418_;
 wire net10723;
 wire net10713;
 wire net10439;
 wire _11422_;
 wire net10739;
 wire net10444;
 wire net10442;
 wire net10433;
 wire _11427_;
 wire _11428_;
 wire net10727;
 wire _11430_;
 wire net10432;
 wire _11432_;
 wire _11433_;
 wire net10425;
 wire net10729;
 wire _11436_;
 wire net10431;
 wire _11438_;
 wire _11439_;
 wire net10420;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire net10419;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire net10422;
 wire net10409;
 wire net10404;
 wire _11462_;
 wire net10417;
 wire clknet_leaf_248_clk;
 wire _11465_;
 wire _11466_;
 wire net10714;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire net10416;
 wire _11477_;
 wire _11478_;
 wire net10396;
 wire _11480_;
 wire _11481_;
 wire clknet_leaf_247_clk;
 wire _11483_;
 wire _11484_;
 wire clknet_leaf_246_clk;
 wire _11486_;
 wire clknet_leaf_245_clk;
 wire _11488_;
 wire net10448;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire net10430;
 wire _11500_;
 wire _11501_;
 wire net10728;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire net10454;
 wire _11510_;
 wire _11511_;
 wire net10449;
 wire _11513_;
 wire _11514_;
 wire net10423;
 wire _11516_;
 wire _11517_;
 wire net10397;
 wire _11519_;
 wire _11520_;
 wire net10418;
 wire _11522_;
 wire _11523_;
 wire net10403;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire clknet_leaf_266_clk;
 wire _11529_;
 wire _11530_;
 wire clknet_leaf_254_clk;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire net10424;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire net10410;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire net10405;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire net10414;
 wire clknet_leaf_250_clk;
 wire net10402;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire clknet_leaf_265_clk;
 wire _11602_;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_256_clk;
 wire _11605_;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_257_clk;
 wire net10407;
 wire _11611_;
 wire _11612_;
 wire net10401;
 wire net10863;
 wire net10395;
 wire _11616_;
 wire net10747;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire net10400;
 wire _11625_;
 wire net10799;
 wire net10864;
 wire net10408;
 wire net10394;
 wire _11630_;
 wire net10438;
 wire net10443;
 wire _11633_;
 wire _11634_;
 wire net10385;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire net10427;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire net10801;
 wire _11680_;
 wire net10413;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire net10426;
 wire net10412;
 wire _11689_;
 wire _11690_;
 wire net10599;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire net10737;
 wire _11735_;
 wire net10708;
 wire _11737_;
 wire net10659;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire net10384;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire net10382;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire net10389;
 wire _11794_;
 wire _11795_;
 wire net10738;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire net10406;
 wire _11808_;
 wire net10731;
 wire net10434;
 wire net10399;
 wire net10730;
 wire _11813_;
 wire _11814_;
 wire net10367;
 wire net10366;
 wire _11817_;
 wire net10383;
 wire _11819_;
 wire _11820_;
 wire net10804;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire net10437;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire net10373;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire net10435;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire clknet_leaf_268_clk;
 wire _11838_;
 wire clknet_leaf_267_clk;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire net10371;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire net10362;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire net10451;
 wire net10381;
 wire _11854_;
 wire net10392;
 wire _11856_;
 wire _11857_;
 wire net10369;
 wire _11859_;
 wire net10363;
 wire net10365;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire net10370;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire net10388;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire net10368;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire net10386;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire net10358;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire net10387;
 wire _11887_;
 wire net10364;
 wire _11889_;
 wire net10380;
 wire _11891_;
 wire _11892_;
 wire net10357;
 wire _11894_;
 wire _11895_;
 wire net10372;
 wire _11897_;
 wire _11898_;
 wire net10334;
 wire _11900_;
 wire net10345;
 wire _11902_;
 wire net10348;
 wire _11904_;
 wire _11905_;
 wire net10343;
 wire _11907_;
 wire net10350;
 wire net10356;
 wire net10354;
 wire net10374;
 wire net10359;
 wire _11913_;
 wire net10355;
 wire _11915_;
 wire _11916_;
 wire net10335;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire net10361;
 wire _11928_;
 wire net10338;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire net10375;
 wire _11937_;
 wire _11938_;
 wire net10337;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire net10336;
 wire clknet_leaf_269_clk;
 wire net10325;
 wire net10317;
 wire _11948_;
 wire net10324;
 wire net10360;
 wire _11951_;
 wire _11952_;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_270_clk;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire net10318;
 wire net10323;
 wire net10311;
 wire net10320;
 wire net10310;
 wire net10314;
 wire net10322;
 wire net10313;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire net10312;
 wire net10306;
 wire net10321;
 wire net10305;
 wire net10308;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_272_clk;
 wire _11984_;
 wire net10316;
 wire net10300;
 wire _11987_;
 wire _11988_;
 wire net10319;
 wire net10298;
 wire net10344;
 wire _11992_;
 wire _11993_;
 wire net10303;
 wire _11995_;
 wire _11996_;
 wire net10309;
 wire net10302;
 wire clknet_leaf_276_clk;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire net10301;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire net10295;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire net10297;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire net10292;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire net10293;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire net10299;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire clk;
 wire gpio_in1;
 wire gpio_in2;
 wire gpio_io1_oe;
 wire gpio_io2_oe;
 wire gpio_out1;
 wire gpio_out2;
 wire pwm_out;
 wire resetn;
 wire ser_rx;
 wire ser_tx;
 wire spi_flash_clk;
 wire spi_flash_cs_n;
 wire spi_flash_io0_di;
 wire spi_flash_io0_do;
 wire spi_flash_io0_oe;
 wire spi_flash_io1_di;
 wire spi_flash_io1_do;
 wire spi_flash_io1_oe;
 wire spi_flash_io2_di;
 wire spi_flash_io2_do;
 wire spi_flash_io2_oe;
 wire spi_flash_io3_di;
 wire spi_flash_io3_do;
 wire spi_flash_io3_oe;
 wire spi_sensor_clk;
 wire spi_sensor_cs_n;
 wire spi_sensor_miso;
 wire spi_sensor_mosi;
 wire \u_ac_controller_soc_inst.cbus_addr[10] ;
 wire \u_ac_controller_soc_inst.cbus_addr[11] ;
 wire \u_ac_controller_soc_inst.cbus_addr[12] ;
 wire \u_ac_controller_soc_inst.cbus_addr[13] ;
 wire \u_ac_controller_soc_inst.cbus_addr[14] ;
 wire \u_ac_controller_soc_inst.cbus_addr[15] ;
 wire \u_ac_controller_soc_inst.cbus_addr[16] ;
 wire \u_ac_controller_soc_inst.cbus_addr[17] ;
 wire \u_ac_controller_soc_inst.cbus_addr[18] ;
 wire \u_ac_controller_soc_inst.cbus_addr[19] ;
 wire \u_ac_controller_soc_inst.cbus_addr[20] ;
 wire \u_ac_controller_soc_inst.cbus_addr[21] ;
 wire \u_ac_controller_soc_inst.cbus_addr[22] ;
 wire \u_ac_controller_soc_inst.cbus_addr[23] ;
 wire \u_ac_controller_soc_inst.cbus_addr[24] ;
 wire \u_ac_controller_soc_inst.cbus_addr[25] ;
 wire \u_ac_controller_soc_inst.cbus_addr[26] ;
 wire \u_ac_controller_soc_inst.cbus_addr[27] ;
 wire \u_ac_controller_soc_inst.cbus_addr[28] ;
 wire \u_ac_controller_soc_inst.cbus_addr[29] ;
 wire \u_ac_controller_soc_inst.cbus_addr[2] ;
 wire \u_ac_controller_soc_inst.cbus_addr[30] ;
 wire \u_ac_controller_soc_inst.cbus_addr[31] ;
 wire \u_ac_controller_soc_inst.cbus_addr[3] ;
 wire \u_ac_controller_soc_inst.cbus_addr[4] ;
 wire \u_ac_controller_soc_inst.cbus_addr[5] ;
 wire \u_ac_controller_soc_inst.cbus_addr[6] ;
 wire \u_ac_controller_soc_inst.cbus_addr[7] ;
 wire \u_ac_controller_soc_inst.cbus_addr[8] ;
 wire \u_ac_controller_soc_inst.cbus_addr[9] ;
 wire \u_ac_controller_soc_inst.cbus_valid ;
 wire \u_ac_controller_soc_inst.cbus_wdata[0] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[10] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[11] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[12] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[13] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[14] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[15] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[16] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[17] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[18] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[19] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[1] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[20] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[21] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[22] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[23] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[24] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[25] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[26] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[27] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[28] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[29] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[2] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[30] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[31] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[3] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[4] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[5] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[6] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[7] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[8] ;
 wire \u_ac_controller_soc_inst.cbus_wdata[9] ;
 wire \u_ac_controller_soc_inst.cbus_wstrb[0] ;
 wire \u_ac_controller_soc_inst.cbus_wstrb[1] ;
 wire \u_ac_controller_soc_inst.cbus_wstrb[2] ;
 wire \u_ac_controller_soc_inst.cbus_wstrb[3] ;
 wire \u_ac_controller_soc_inst.io_rdata[0] ;
 wire \u_ac_controller_soc_inst.io_rdata[10] ;
 wire \u_ac_controller_soc_inst.io_rdata[11] ;
 wire \u_ac_controller_soc_inst.io_rdata[12] ;
 wire \u_ac_controller_soc_inst.io_rdata[13] ;
 wire \u_ac_controller_soc_inst.io_rdata[14] ;
 wire \u_ac_controller_soc_inst.io_rdata[15] ;
 wire \u_ac_controller_soc_inst.io_rdata[16] ;
 wire \u_ac_controller_soc_inst.io_rdata[17] ;
 wire \u_ac_controller_soc_inst.io_rdata[18] ;
 wire \u_ac_controller_soc_inst.io_rdata[19] ;
 wire \u_ac_controller_soc_inst.io_rdata[1] ;
 wire \u_ac_controller_soc_inst.io_rdata[20] ;
 wire \u_ac_controller_soc_inst.io_rdata[21] ;
 wire \u_ac_controller_soc_inst.io_rdata[22] ;
 wire \u_ac_controller_soc_inst.io_rdata[23] ;
 wire \u_ac_controller_soc_inst.io_rdata[24] ;
 wire \u_ac_controller_soc_inst.io_rdata[25] ;
 wire \u_ac_controller_soc_inst.io_rdata[26] ;
 wire \u_ac_controller_soc_inst.io_rdata[27] ;
 wire \u_ac_controller_soc_inst.io_rdata[28] ;
 wire \u_ac_controller_soc_inst.io_rdata[29] ;
 wire \u_ac_controller_soc_inst.io_rdata[2] ;
 wire \u_ac_controller_soc_inst.io_rdata[30] ;
 wire \u_ac_controller_soc_inst.io_rdata[31] ;
 wire \u_ac_controller_soc_inst.io_rdata[3] ;
 wire \u_ac_controller_soc_inst.io_rdata[4] ;
 wire \u_ac_controller_soc_inst.io_rdata[5] ;
 wire \u_ac_controller_soc_inst.io_rdata[6] ;
 wire \u_ac_controller_soc_inst.io_rdata[7] ;
 wire \u_ac_controller_soc_inst.io_rdata[8] ;
 wire \u_ac_controller_soc_inst.io_rdata[9] ;
 wire \u_ac_controller_soc_inst.io_ready ;
 wire \u_ac_controller_soc_inst.spi_flash_cfg_rdata[16] ;
 wire \u_ac_controller_soc_inst.spi_flash_cfg_rdata[17] ;
 wire \u_ac_controller_soc_inst.spi_flash_cfg_rdata[18] ;
 wire \u_ac_controller_soc_inst.spi_flash_cfg_rdata[19] ;
 wire \u_ac_controller_soc_inst.spi_flash_cfg_rdata[20] ;
 wire \u_ac_controller_soc_inst.spi_flash_cfg_rdata[21] ;
 wire \u_ac_controller_soc_inst.spi_flash_cfg_rdata[22] ;
 wire \u_ac_controller_soc_inst.spi_flash_cfg_rdata[31] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[0] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[10] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[11] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[12] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[13] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[14] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[15] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[16] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[17] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[18] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[19] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[1] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[20] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[21] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[22] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[23] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[24] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[25] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[26] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[27] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[28] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[29] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[2] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[30] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[31] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[3] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[4] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[5] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[6] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[7] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[8] ;
 wire \u_ac_controller_soc_inst.spi_flash_rdata[9] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[0] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[10] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[11] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[12] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[13] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[14] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[15] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[16] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[17] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[18] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[19] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[1] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[20] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[21] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[22] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[23] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[24] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[25] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[26] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[27] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[28] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[29] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[2] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[30] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[31] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[3] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[4] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[5] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[6] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[7] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[8] ;
 wire \u_ac_controller_soc_inst.spi_sensor_rdata[9] ;
 wire \u_ac_controller_soc_inst.spi_sensor_ready ;
 wire \u_ac_controller_soc_inst.sram_ready ;
 wire \u_ac_controller_soc_inst.trap ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[11] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[12] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[13] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[15] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[16] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[17] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[18] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[19] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[20] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[23] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[25] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[27] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[28] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[29] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[30] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[31] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[6] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[7] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[8] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[10] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[11] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[12] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[13] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[14] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[15] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[16] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[17] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[18] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[19] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[20] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[21] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[22] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[23] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[24] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[25] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[26] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[27] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[28] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[29] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[30] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[31] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[6] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[7] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[8] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[9] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in1_sync ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in1_sync1 ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in2_sync ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in2_sync1 ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[10] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[11] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[12] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[13] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[14] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[15] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[16] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[17] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[18] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[19] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[20] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[21] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[22] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[23] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[24] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[25] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[26] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[27] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[28] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[29] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[30] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[31] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[6] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[7] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[8] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[9] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_enable ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[10] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[11] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[12] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[13] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[14] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[15] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[16] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[17] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[18] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[19] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[20] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[21] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[22] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[23] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[24] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[25] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[26] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[27] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[28] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[29] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[30] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[31] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[6] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[7] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[8] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[9] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[10] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[11] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[12] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[13] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[14] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[15] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[16] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[17] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[18] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[19] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[20] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[21] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[22] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[23] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[24] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[25] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[26] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[27] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[28] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[29] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[30] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[31] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[32] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[33] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[34] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[35] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[36] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[37] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[38] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[39] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[6] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[7] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[8] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[9] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[10] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[11] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[12] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[15] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[16] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[17] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[18] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[19] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[20] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[21] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[23] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[24] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[25] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[26] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[27] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[28] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[29] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[30] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[31] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[6] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[7] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[8] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[6] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[7] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[8] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync1 ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.start_bit ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.stop_bit ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[6] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[7] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[8] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_ready ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[10] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[11] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[12] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[13] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[14] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[15] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[16] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[17] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[18] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[19] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[20] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[21] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[22] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[23] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[24] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[25] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[26] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[27] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[28] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[29] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[30] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[31] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[6] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[7] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[8] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[9] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_done ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[0] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[10] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[11] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[12] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[13] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[14] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[15] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[16] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[17] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[18] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[19] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[1] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[20] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[21] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[22] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[23] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[24] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[25] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[26] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[27] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[28] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[29] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[2] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[30] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[31] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[3] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[4] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[5] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[6] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[7] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[8] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[9] ;
 wire \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfering ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.alu_out_q[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[32] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[33] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[34] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[35] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[36] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[37] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[38] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[39] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[40] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[41] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[42] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[43] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[44] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[45] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[46] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[47] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[48] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[49] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[50] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[51] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[52] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[53] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[54] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[55] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[56] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[57] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[58] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[59] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[60] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[61] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[62] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[63] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_cycle[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[32] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[33] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[34] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[35] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[36] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[37] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[38] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[39] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[40] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[41] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[42] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[43] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[44] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[45] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[46] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[47] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[48] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[49] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[50] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[51] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[52] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[53] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[54] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[55] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[56] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[57] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[58] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[59] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[60] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[61] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[62] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[63] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.count_instr[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpu_state[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpu_state[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpu_state[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpu_state[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpu_state[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpu_state[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpu_state[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_rd[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_rd[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_rd[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_rd[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoded_rd[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoder_pseudo_trigger ;
 wire \u_ac_controller_soc_inst.u_picorv32.decoder_trigger ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_add ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_addi ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_and ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_andi ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_auipc ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_beq ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_bge ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_bgeu ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_blt ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_bltu ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_bne ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_fence ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_jal ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_jalr ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_lb ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_lbu ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_lh ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_lhu ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_lui ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_lw ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_or ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_ori ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_rdcycle ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_rdcycleh ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_rdinstr ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_sb ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_sh ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_sll ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_slli ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_slt ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_slti ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_sltiu ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_sltu ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_sra ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_srai ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_srl ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_srli ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_sub ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_sw ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_xor ;
 wire \u_ac_controller_soc_inst.u_picorv32.instr_xori ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_alu_reg_imm ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_alu_reg_reg ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_beq_bne_blt_bge_bltu_bgeu ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_compare ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_jalr_addi_slti_sltiu_xori_ori_andi ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_lb_lh_lw_lbu_lhu ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_lui_auipc_jal ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_sb_sh_sw ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_sll_srl_sra ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_slli_srli_srai ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_slti_blt_slt ;
 wire \u_ac_controller_soc_inst.u_picorv32.is_sltiu_bltu_sltu ;
 wire \u_ac_controller_soc_inst.u_picorv32.latched_branch ;
 wire \u_ac_controller_soc_inst.u_picorv32.latched_is_lb ;
 wire \u_ac_controller_soc_inst.u_picorv32.latched_is_lh ;
 wire \u_ac_controller_soc_inst.u_picorv32.latched_rd[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.latched_rd[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.latched_rd[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.latched_rd[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.latched_rd[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.latched_stalu ;
 wire \u_ac_controller_soc_inst.u_picorv32.latched_store ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_do_prefetch ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_do_rdata ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_do_rinst ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_do_wdata ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[11] ;
 wire clknet_leaf_446_clk;
 wire clknet_leaf_452_clk;
 wire clknet_leaf_443_clk;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_state[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_state[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_wordsize[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_wordsize[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.mem_wordsize[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_out[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[10] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[11] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[12] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[13] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[14] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[15] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[16] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[17] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[18] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[19] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[20] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[21] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[22] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[23] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[24] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[25] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[26] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[27] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[28] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[29] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[30] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[31] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[4] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[5] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[6] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[7] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[8] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_pc[9] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_sh[0] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_sh[1] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_sh[2] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_sh[3] ;
 wire \u_ac_controller_soc_inst.u_picorv32.reg_sh[4] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[10] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[11] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[12] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[13] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[14] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[15] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[16] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[17] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[18] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[19] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[20] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[21] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[22] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[23] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[3] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[4] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[5] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[6] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[7] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[8] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[9] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.config_clk ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.config_csb ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[3] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[3] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[3] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[4] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[5] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[6] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[7] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_ddr ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_qspi ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_rd ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.din_valid ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[3] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[4] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[5] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[6] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[7] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[10] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[11] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[12] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[13] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[14] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[16] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[17] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[18] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[22] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[3] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[4] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[5] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[6] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[7] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[8] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[9] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_inc ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_valid ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.rd_wait ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.softreset ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[10] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[11] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[12] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[3] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[4] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[5] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[6] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[7] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[8] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.state[9] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[3] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[3] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.fetch ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_csb ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io0_do ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io1_do ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io2_do ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io3_do ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.last_fetch ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[3] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[4] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[5] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[6] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[7] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.resetn ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr_q ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_qspi ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_rd ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[0] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[1] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[2] ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io0_90 ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io1_90 ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io2_90 ;
 wire \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io3_90 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire clknet_leaf_833_clk;
 wire clknet_leaf_834_clk;
 wire clknet_leaf_835_clk;
 wire clknet_leaf_836_clk;
 wire clknet_leaf_837_clk;
 wire clknet_leaf_838_clk;
 wire clknet_leaf_840_clk;
 wire clknet_leaf_841_clk;
 wire clknet_leaf_842_clk;
 wire clknet_leaf_845_clk;
 wire clknet_leaf_847_clk;
 wire clknet_leaf_848_clk;
 wire clknet_leaf_849_clk;
 wire clknet_leaf_850_clk;
 wire clknet_leaf_851_clk;
 wire clknet_leaf_852_clk;
 wire clknet_leaf_853_clk;
 wire clknet_leaf_854_clk;
 wire clknet_leaf_857_clk;
 wire clknet_leaf_858_clk;
 wire clknet_leaf_859_clk;
 wire clknet_leaf_860_clk;
 wire clknet_leaf_861_clk;
 wire clknet_leaf_863_clk;
 wire clknet_leaf_865_clk;
 wire clknet_leaf_867_clk;
 wire clknet_leaf_868_clk;
 wire clknet_leaf_869_clk;
 wire clknet_leaf_870_clk;
 wire clknet_leaf_873_clk;
 wire clknet_leaf_874_clk;
 wire clknet_leaf_875_clk;
 wire clknet_leaf_877_clk;
 wire clknet_leaf_878_clk;
 wire clknet_leaf_879_clk;
 wire clknet_leaf_882_clk;
 wire clknet_leaf_883_clk;
 wire clknet_leaf_884_clk;
 wire clknet_leaf_886_clk;
 wire clknet_leaf_887_clk;
 wire clknet_leaf_888_clk;
 wire clknet_leaf_890_clk;
 wire clknet_leaf_891_clk;
 wire clknet_leaf_892_clk;
 wire clknet_leaf_893_clk;
 wire clknet_leaf_894_clk;
 wire clknet_leaf_896_clk;
 wire clknet_leaf_898_clk;
 wire clknet_leaf_899_clk;
 wire clknet_leaf_900_clk;
 wire clknet_leaf_902_clk;
 wire clknet_leaf_903_clk;
 wire clknet_leaf_904_clk;
 wire clknet_leaf_905_clk;
 wire clknet_leaf_907_clk;
 wire clknet_leaf_909_clk;
 wire clknet_leaf_910_clk;
 wire clknet_leaf_912_clk;
 wire clknet_leaf_914_clk;
 wire clknet_leaf_916_clk;
 wire clknet_leaf_917_clk;
 wire clknet_leaf_920_clk;
 wire clknet_leaf_921_clk;
 wire clknet_leaf_923_clk;
 wire clknet_leaf_924_clk;
 wire clknet_leaf_926_clk;
 wire clknet_leaf_927_clk;
 wire clknet_leaf_929_clk;
 wire clknet_leaf_930_clk;
 wire clknet_leaf_931_clk;
 wire clknet_leaf_932_clk;
 wire clknet_leaf_933_clk;
 wire clknet_leaf_934_clk;
 wire clknet_leaf_935_clk;
 wire clknet_leaf_936_clk;
 wire clknet_leaf_937_clk;
 wire clknet_leaf_938_clk;
 wire clknet_leaf_941_clk;
 wire clknet_leaf_942_clk;
 wire clknet_leaf_943_clk;
 wire clknet_leaf_946_clk;
 wire clknet_leaf_948_clk;
 wire clknet_leaf_949_clk;
 wire clknet_leaf_951_clk;
 wire clknet_leaf_952_clk;
 wire clknet_leaf_953_clk;
 wire clknet_leaf_954_clk;
 wire clknet_leaf_955_clk;
 wire clknet_leaf_956_clk;
 wire clknet_leaf_957_clk;
 wire clknet_leaf_960_clk;
 wire clknet_leaf_961_clk;
 wire clknet_leaf_962_clk;
 wire clknet_leaf_963_clk;
 wire clknet_leaf_965_clk;
 wire clknet_leaf_966_clk;
 wire clknet_leaf_968_clk;
 wire clknet_leaf_969_clk;
 wire clknet_leaf_972_clk;
 wire clknet_leaf_974_clk;
 wire clknet_leaf_978_clk;
 wire clknet_leaf_982_clk;
 wire clknet_leaf_988_clk;
 wire clknet_leaf_990_clk;
 wire clknet_leaf_991_clk;
 wire clknet_leaf_994_clk;
 wire clknet_leaf_995_clk;
 wire clknet_leaf_997_clk;
 wire clknet_leaf_998_clk;
 wire clknet_leaf_999_clk;
 wire clknet_leaf_1000_clk;
 wire clknet_leaf_1003_clk;
 wire clknet_leaf_1004_clk;
 wire clknet_leaf_1005_clk;
 wire clknet_leaf_1006_clk;
 wire clknet_leaf_1007_clk;
 wire clknet_leaf_1009_clk;
 wire clknet_leaf_1010_clk;
 wire clknet_leaf_1011_clk;
 wire clknet_leaf_1012_clk;
 wire clknet_leaf_1015_clk;
 wire clknet_leaf_1017_clk;
 wire clknet_leaf_1018_clk;
 wire clknet_leaf_1019_clk;
 wire clknet_leaf_1020_clk;
 wire clknet_leaf_1021_clk;
 wire clknet_leaf_1022_clk;
 wire clknet_leaf_1023_clk;
 wire clknet_leaf_1026_clk;
 wire clknet_leaf_1027_clk;
 wire clknet_leaf_1028_clk;
 wire clknet_leaf_1031_clk;
 wire clknet_leaf_1032_clk;
 wire clknet_leaf_1033_clk;
 wire clknet_leaf_1034_clk;
 wire clknet_leaf_1035_clk;
 wire clknet_leaf_1037_clk;
 wire clknet_leaf_1038_clk;
 wire clknet_leaf_1040_clk;
 wire clknet_leaf_1041_clk;
 wire clknet_leaf_1043_clk;
 wire clknet_leaf_1044_clk;
 wire clknet_leaf_1045_clk;
 wire clknet_leaf_1046_clk;
 wire clknet_leaf_1047_clk;
 wire clknet_leaf_1048_clk;
 wire clknet_leaf_1049_clk;
 wire clknet_leaf_1051_clk;
 wire clknet_leaf_1052_clk;
 wire clknet_leaf_1053_clk;
 wire clknet_leaf_1054_clk;
 wire clknet_leaf_1055_clk;
 wire clknet_leaf_1056_clk;
 wire clknet_leaf_1057_clk;
 wire clknet_leaf_1058_clk;
 wire clknet_leaf_1060_clk;
 wire clknet_leaf_1061_clk;
 wire clknet_leaf_1062_clk;
 wire clknet_leaf_1063_clk;
 wire clknet_leaf_1065_clk;
 wire clknet_leaf_1066_clk;
 wire clknet_leaf_1067_clk;
 wire clknet_leaf_1069_clk;
 wire clknet_leaf_1070_clk;
 wire clknet_leaf_1071_clk;
 wire clknet_leaf_1072_clk;
 wire clknet_leaf_1073_clk;
 wire clknet_leaf_1074_clk;
 wire clknet_leaf_1075_clk;
 wire clknet_leaf_1076_clk;
 wire clknet_leaf_1077_clk;
 wire clknet_leaf_1078_clk;
 wire clknet_leaf_1079_clk;
 wire clknet_leaf_1080_clk;
 wire clknet_leaf_1081_clk;
 wire clknet_leaf_1083_clk;
 wire clknet_leaf_1084_clk;
 wire clknet_leaf_1085_clk;
 wire clknet_leaf_1086_clk;
 wire clknet_leaf_1087_clk;
 wire clknet_leaf_1088_clk;
 wire clknet_leaf_1089_clk;
 wire clknet_leaf_1090_clk;
 wire clknet_leaf_1091_clk;
 wire clknet_leaf_1092_clk;
 wire clknet_leaf_1093_clk;
 wire clknet_leaf_1096_clk;
 wire clknet_leaf_1097_clk;
 wire clknet_leaf_1098_clk;
 wire clknet_leaf_1099_clk;
 wire clknet_leaf_1101_clk;
 wire clknet_leaf_1104_clk;
 wire clknet_leaf_1105_clk;
 wire clknet_leaf_1106_clk;
 wire clknet_leaf_1109_clk;
 wire clknet_leaf_1110_clk;
 wire clknet_leaf_1112_clk;
 wire clknet_leaf_1113_clk;
 wire clknet_leaf_1114_clk;
 wire clknet_leaf_1116_clk;
 wire clknet_leaf_1120_clk;
 wire clknet_leaf_1122_clk;
 wire clknet_leaf_1124_clk;
 wire clknet_leaf_1125_clk;
 wire clknet_leaf_1126_clk;
 wire clknet_leaf_1127_clk;
 wire clknet_leaf_1128_clk;
 wire clknet_leaf_1129_clk;
 wire clknet_leaf_1131_clk;
 wire clknet_leaf_1133_clk;
 wire clknet_leaf_1134_clk;
 wire clknet_leaf_1135_clk;
 wire clknet_leaf_1136_clk;
 wire clknet_leaf_1138_clk;
 wire clknet_leaf_1139_clk;
 wire clknet_leaf_1140_clk;
 wire clknet_leaf_1142_clk;
 wire clknet_leaf_1144_clk;
 wire clknet_leaf_1145_clk;
 wire clknet_leaf_1146_clk;
 wire clknet_leaf_1147_clk;
 wire clknet_leaf_1148_clk;
 wire clknet_leaf_1149_clk;
 wire clknet_leaf_1150_clk;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_0_1_clk;
 wire clknet_1_1_0_clk;
 wire clknet_1_1_1_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_0_1_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_1_1_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_2_1_clk;
 wire clknet_2_3_0_clk;
 wire clknet_2_3_1_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0_0_clk;
 wire clknet_5_1_0_clk;
 wire clknet_5_2_0_clk;
 wire clknet_5_3_0_clk;
 wire clknet_5_4_0_clk;
 wire clknet_5_5_0_clk;
 wire clknet_5_6_0_clk;
 wire clknet_5_7_0_clk;
 wire clknet_5_8_0_clk;
 wire clknet_5_9_0_clk;
 wire clknet_5_10_0_clk;
 wire clknet_5_11_0_clk;
 wire clknet_5_12_0_clk;
 wire clknet_5_13_0_clk;
 wire clknet_5_14_0_clk;
 wire clknet_5_15_0_clk;
 wire clknet_5_16_0_clk;
 wire clknet_5_17_0_clk;
 wire clknet_5_18_0_clk;
 wire clknet_5_19_0_clk;
 wire clknet_5_20_0_clk;
 wire clknet_5_21_0_clk;
 wire clknet_5_22_0_clk;
 wire clknet_5_23_0_clk;
 wire clknet_5_24_0_clk;
 wire clknet_5_25_0_clk;
 wire clknet_5_26_0_clk;
 wire clknet_5_27_0_clk;
 wire clknet_5_28_0_clk;
 wire clknet_5_29_0_clk;
 wire clknet_5_30_0_clk;
 wire clknet_5_31_0_clk;
 wire clknet_6_0_0_clk;
 wire clknet_6_1_0_clk;
 wire clknet_6_2_0_clk;
 wire clknet_6_3_0_clk;
 wire clknet_6_4_0_clk;
 wire clknet_6_5_0_clk;
 wire clknet_6_6_0_clk;
 wire clknet_6_7_0_clk;
 wire clknet_6_8_0_clk;
 wire clknet_6_9_0_clk;
 wire clknet_6_10_0_clk;
 wire clknet_6_11_0_clk;
 wire clknet_6_12_0_clk;
 wire clknet_6_13_0_clk;
 wire clknet_6_14_0_clk;
 wire clknet_6_15_0_clk;
 wire clknet_6_16_0_clk;
 wire clknet_6_17_0_clk;
 wire clknet_6_18_0_clk;
 wire clknet_6_19_0_clk;
 wire clknet_6_20_0_clk;
 wire clknet_6_21_0_clk;
 wire clknet_6_22_0_clk;
 wire clknet_6_23_0_clk;
 wire clknet_6_24_0_clk;
 wire clknet_6_25_0_clk;
 wire clknet_6_26_0_clk;
 wire clknet_6_27_0_clk;
 wire clknet_6_28_0_clk;
 wire clknet_6_29_0_clk;
 wire clknet_6_30_0_clk;
 wire clknet_6_31_0_clk;
 wire clknet_6_32_0_clk;
 wire clknet_6_33_0_clk;
 wire clknet_6_34_0_clk;
 wire clknet_6_35_0_clk;
 wire clknet_6_36_0_clk;
 wire clknet_6_37_0_clk;
 wire clknet_6_38_0_clk;
 wire clknet_6_39_0_clk;
 wire clknet_6_40_0_clk;
 wire clknet_6_41_0_clk;
 wire clknet_6_42_0_clk;
 wire clknet_6_43_0_clk;
 wire clknet_6_44_0_clk;
 wire clknet_6_45_0_clk;
 wire clknet_6_46_0_clk;
 wire clknet_6_47_0_clk;
 wire clknet_6_48_0_clk;
 wire clknet_6_49_0_clk;
 wire clknet_6_50_0_clk;
 wire clknet_6_51_0_clk;
 wire clknet_6_52_0_clk;
 wire clknet_6_53_0_clk;
 wire clknet_6_54_0_clk;
 wire clknet_6_55_0_clk;
 wire clknet_6_56_0_clk;
 wire clknet_6_57_0_clk;
 wire clknet_6_58_0_clk;
 wire clknet_6_59_0_clk;
 wire clknet_6_60_0_clk;
 wire clknet_6_61_0_clk;
 wire clknet_6_62_0_clk;
 wire clknet_6_63_0_clk;
 wire clknet_7_0_0_clk;
 wire clknet_7_1_0_clk;
 wire clknet_7_2_0_clk;
 wire clknet_7_3_0_clk;
 wire clknet_7_4_0_clk;
 wire clknet_7_5_0_clk;
 wire clknet_7_6_0_clk;
 wire clknet_7_7_0_clk;
 wire clknet_7_8_0_clk;
 wire clknet_7_9_0_clk;
 wire clknet_7_10_0_clk;
 wire clknet_7_11_0_clk;
 wire clknet_7_12_0_clk;
 wire clknet_7_13_0_clk;
 wire clknet_7_14_0_clk;
 wire clknet_7_15_0_clk;
 wire clknet_7_16_0_clk;
 wire clknet_7_17_0_clk;
 wire clknet_7_18_0_clk;
 wire clknet_7_19_0_clk;
 wire clknet_7_20_0_clk;
 wire clknet_7_21_0_clk;
 wire clknet_7_22_0_clk;
 wire clknet_7_23_0_clk;
 wire clknet_7_24_0_clk;
 wire clknet_7_25_0_clk;
 wire clknet_7_26_0_clk;
 wire clknet_7_27_0_clk;
 wire clknet_7_28_0_clk;
 wire clknet_7_29_0_clk;
 wire clknet_7_30_0_clk;
 wire clknet_7_31_0_clk;
 wire clknet_7_32_0_clk;
 wire clknet_7_33_0_clk;
 wire clknet_7_34_0_clk;
 wire clknet_7_35_0_clk;
 wire clknet_7_36_0_clk;
 wire clknet_7_37_0_clk;
 wire clknet_7_38_0_clk;
 wire clknet_7_39_0_clk;
 wire clknet_7_40_0_clk;
 wire clknet_7_41_0_clk;
 wire clknet_7_42_0_clk;
 wire clknet_7_43_0_clk;
 wire clknet_7_44_0_clk;
 wire clknet_7_45_0_clk;
 wire clknet_7_46_0_clk;
 wire clknet_7_47_0_clk;
 wire clknet_7_48_0_clk;
 wire clknet_7_49_0_clk;
 wire clknet_7_50_0_clk;
 wire clknet_7_51_0_clk;
 wire clknet_7_52_0_clk;
 wire clknet_7_53_0_clk;
 wire clknet_7_54_0_clk;
 wire clknet_7_55_0_clk;
 wire clknet_7_56_0_clk;
 wire clknet_7_57_0_clk;
 wire clknet_7_58_0_clk;
 wire clknet_7_59_0_clk;
 wire clknet_7_60_0_clk;
 wire clknet_7_61_0_clk;
 wire clknet_7_62_0_clk;
 wire clknet_7_63_0_clk;
 wire clknet_7_64_0_clk;
 wire clknet_7_65_0_clk;
 wire clknet_7_66_0_clk;
 wire clknet_7_67_0_clk;
 wire clknet_7_68_0_clk;
 wire clknet_7_69_0_clk;
 wire clknet_7_70_0_clk;
 wire clknet_7_71_0_clk;
 wire clknet_7_72_0_clk;
 wire clknet_7_73_0_clk;
 wire clknet_7_74_0_clk;
 wire clknet_7_75_0_clk;
 wire clknet_7_76_0_clk;
 wire clknet_7_77_0_clk;
 wire clknet_7_78_0_clk;
 wire clknet_7_79_0_clk;
 wire clknet_7_80_0_clk;
 wire clknet_7_81_0_clk;
 wire clknet_7_82_0_clk;
 wire clknet_7_83_0_clk;
 wire clknet_7_84_0_clk;
 wire clknet_7_85_0_clk;
 wire clknet_7_86_0_clk;
 wire clknet_7_87_0_clk;
 wire clknet_7_88_0_clk;
 wire clknet_7_89_0_clk;
 wire clknet_7_90_0_clk;
 wire clknet_7_91_0_clk;
 wire clknet_7_92_0_clk;
 wire clknet_7_93_0_clk;
 wire clknet_7_94_0_clk;
 wire clknet_7_95_0_clk;
 wire clknet_7_96_0_clk;
 wire clknet_7_97_0_clk;
 wire clknet_7_98_0_clk;
 wire clknet_7_99_0_clk;
 wire clknet_7_100_0_clk;
 wire clknet_7_101_0_clk;
 wire clknet_7_102_0_clk;
 wire clknet_7_103_0_clk;
 wire clknet_7_104_0_clk;
 wire clknet_7_105_0_clk;
 wire clknet_7_106_0_clk;
 wire clknet_7_107_0_clk;
 wire clknet_7_108_0_clk;
 wire clknet_7_109_0_clk;
 wire clknet_7_110_0_clk;
 wire clknet_7_111_0_clk;
 wire clknet_7_112_0_clk;
 wire clknet_7_113_0_clk;
 wire clknet_7_114_0_clk;
 wire clknet_7_115_0_clk;
 wire clknet_7_116_0_clk;
 wire clknet_7_117_0_clk;
 wire clknet_7_118_0_clk;
 wire clknet_7_119_0_clk;
 wire clknet_7_120_0_clk;
 wire clknet_7_121_0_clk;
 wire clknet_7_122_0_clk;
 wire clknet_7_123_0_clk;
 wire clknet_7_124_0_clk;
 wire clknet_7_125_0_clk;
 wire clknet_7_126_0_clk;
 wire clknet_7_127_0_clk;
 wire clknet_8_0_0_clk;
 wire clknet_8_1_0_clk;
 wire clknet_8_2_0_clk;
 wire clknet_8_3_0_clk;
 wire clknet_8_4_0_clk;
 wire clknet_8_5_0_clk;
 wire clknet_8_6_0_clk;
 wire clknet_8_7_0_clk;
 wire clknet_8_8_0_clk;
 wire clknet_8_9_0_clk;
 wire clknet_8_10_0_clk;
 wire clknet_8_11_0_clk;
 wire clknet_8_12_0_clk;
 wire clknet_8_13_0_clk;
 wire clknet_8_14_0_clk;
 wire clknet_8_15_0_clk;
 wire clknet_8_16_0_clk;
 wire clknet_8_17_0_clk;
 wire clknet_8_18_0_clk;
 wire clknet_8_19_0_clk;
 wire clknet_8_20_0_clk;
 wire clknet_8_21_0_clk;
 wire clknet_8_22_0_clk;
 wire clknet_8_23_0_clk;
 wire clknet_8_24_0_clk;
 wire clknet_8_25_0_clk;
 wire clknet_8_26_0_clk;
 wire clknet_8_27_0_clk;
 wire clknet_8_28_0_clk;
 wire clknet_8_29_0_clk;
 wire clknet_8_30_0_clk;
 wire clknet_8_31_0_clk;
 wire clknet_8_32_0_clk;
 wire clknet_8_33_0_clk;
 wire clknet_8_34_0_clk;
 wire clknet_8_35_0_clk;
 wire clknet_8_36_0_clk;
 wire clknet_8_37_0_clk;
 wire clknet_8_38_0_clk;
 wire clknet_8_39_0_clk;
 wire clknet_8_40_0_clk;
 wire clknet_8_41_0_clk;
 wire clknet_8_42_0_clk;
 wire clknet_8_43_0_clk;
 wire clknet_8_44_0_clk;
 wire clknet_8_45_0_clk;
 wire clknet_8_46_0_clk;
 wire clknet_8_47_0_clk;
 wire clknet_8_48_0_clk;
 wire clknet_8_49_0_clk;
 wire clknet_8_50_0_clk;
 wire clknet_8_51_0_clk;
 wire clknet_8_52_0_clk;
 wire clknet_8_53_0_clk;
 wire clknet_8_54_0_clk;
 wire clknet_8_55_0_clk;
 wire clknet_8_56_0_clk;
 wire clknet_8_57_0_clk;
 wire clknet_8_58_0_clk;
 wire clknet_8_59_0_clk;
 wire clknet_8_60_0_clk;
 wire clknet_8_61_0_clk;
 wire clknet_8_62_0_clk;
 wire clknet_8_63_0_clk;
 wire clknet_8_64_0_clk;
 wire clknet_8_65_0_clk;
 wire clknet_8_66_0_clk;
 wire clknet_8_67_0_clk;
 wire clknet_8_68_0_clk;
 wire clknet_8_69_0_clk;
 wire clknet_8_70_0_clk;
 wire clknet_8_71_0_clk;
 wire clknet_8_72_0_clk;
 wire clknet_8_73_0_clk;
 wire clknet_8_74_0_clk;
 wire clknet_8_75_0_clk;
 wire clknet_8_76_0_clk;
 wire clknet_8_77_0_clk;
 wire clknet_8_78_0_clk;
 wire clknet_8_79_0_clk;
 wire clknet_8_80_0_clk;
 wire clknet_8_81_0_clk;
 wire clknet_8_82_0_clk;
 wire clknet_8_83_0_clk;
 wire clknet_8_84_0_clk;
 wire clknet_8_85_0_clk;
 wire clknet_8_86_0_clk;
 wire clknet_8_87_0_clk;
 wire clknet_8_88_0_clk;
 wire clknet_8_89_0_clk;
 wire clknet_8_90_0_clk;
 wire clknet_8_91_0_clk;
 wire clknet_8_92_0_clk;
 wire clknet_8_93_0_clk;
 wire clknet_8_94_0_clk;
 wire clknet_8_95_0_clk;
 wire clknet_8_96_0_clk;
 wire clknet_8_97_0_clk;
 wire clknet_8_98_0_clk;
 wire clknet_8_99_0_clk;
 wire clknet_8_100_0_clk;
 wire clknet_8_101_0_clk;
 wire clknet_8_102_0_clk;
 wire clknet_8_103_0_clk;
 wire clknet_8_104_0_clk;
 wire clknet_8_105_0_clk;
 wire clknet_8_106_0_clk;
 wire clknet_8_107_0_clk;
 wire clknet_8_108_0_clk;
 wire clknet_8_109_0_clk;
 wire clknet_8_110_0_clk;
 wire clknet_8_111_0_clk;
 wire clknet_8_112_0_clk;
 wire clknet_8_113_0_clk;
 wire clknet_8_114_0_clk;
 wire clknet_8_115_0_clk;
 wire clknet_8_116_0_clk;
 wire clknet_8_117_0_clk;
 wire clknet_8_118_0_clk;
 wire clknet_8_119_0_clk;
 wire clknet_8_120_0_clk;
 wire clknet_8_121_0_clk;
 wire clknet_8_122_0_clk;
 wire clknet_8_123_0_clk;
 wire clknet_8_124_0_clk;
 wire clknet_8_125_0_clk;
 wire clknet_8_126_0_clk;
 wire clknet_8_127_0_clk;
 wire clknet_8_128_0_clk;
 wire clknet_8_129_0_clk;
 wire clknet_8_130_0_clk;
 wire clknet_8_131_0_clk;
 wire clknet_8_132_0_clk;
 wire clknet_8_133_0_clk;
 wire clknet_8_134_0_clk;
 wire clknet_8_135_0_clk;
 wire clknet_8_136_0_clk;
 wire clknet_8_137_0_clk;
 wire clknet_8_138_0_clk;
 wire clknet_8_139_0_clk;
 wire clknet_8_140_0_clk;
 wire clknet_8_141_0_clk;
 wire clknet_8_142_0_clk;
 wire clknet_8_143_0_clk;
 wire clknet_8_144_0_clk;
 wire clknet_8_145_0_clk;
 wire clknet_8_146_0_clk;
 wire clknet_8_147_0_clk;
 wire clknet_8_148_0_clk;
 wire clknet_8_149_0_clk;
 wire clknet_8_150_0_clk;
 wire clknet_8_151_0_clk;
 wire clknet_8_152_0_clk;
 wire clknet_8_153_0_clk;
 wire clknet_8_154_0_clk;
 wire clknet_8_155_0_clk;
 wire clknet_8_156_0_clk;
 wire clknet_8_157_0_clk;
 wire clknet_8_158_0_clk;
 wire clknet_8_159_0_clk;
 wire clknet_8_160_0_clk;
 wire clknet_8_161_0_clk;
 wire clknet_8_162_0_clk;
 wire clknet_8_163_0_clk;
 wire clknet_8_164_0_clk;
 wire clknet_8_165_0_clk;
 wire clknet_8_166_0_clk;
 wire clknet_8_167_0_clk;
 wire clknet_8_168_0_clk;
 wire clknet_8_169_0_clk;
 wire clknet_8_170_0_clk;
 wire clknet_8_171_0_clk;
 wire clknet_8_172_0_clk;
 wire clknet_8_173_0_clk;
 wire clknet_8_174_0_clk;
 wire clknet_8_175_0_clk;
 wire clknet_8_176_0_clk;
 wire clknet_8_177_0_clk;
 wire clknet_8_178_0_clk;
 wire clknet_8_179_0_clk;
 wire clknet_8_180_0_clk;
 wire clknet_8_181_0_clk;
 wire clknet_8_182_0_clk;
 wire clknet_8_183_0_clk;
 wire clknet_8_184_0_clk;
 wire clknet_8_185_0_clk;
 wire clknet_8_186_0_clk;
 wire clknet_8_187_0_clk;
 wire clknet_8_188_0_clk;
 wire clknet_8_189_0_clk;
 wire clknet_8_190_0_clk;
 wire clknet_8_191_0_clk;
 wire clknet_8_192_0_clk;
 wire clknet_8_193_0_clk;
 wire clknet_8_194_0_clk;
 wire clknet_8_195_0_clk;
 wire clknet_8_196_0_clk;
 wire clknet_8_197_0_clk;
 wire clknet_8_198_0_clk;
 wire clknet_8_199_0_clk;
 wire clknet_8_200_0_clk;
 wire clknet_8_201_0_clk;
 wire clknet_8_202_0_clk;
 wire clknet_8_203_0_clk;
 wire clknet_8_204_0_clk;
 wire clknet_8_205_0_clk;
 wire clknet_8_206_0_clk;
 wire clknet_8_207_0_clk;
 wire clknet_8_208_0_clk;
 wire clknet_8_209_0_clk;
 wire clknet_8_210_0_clk;
 wire clknet_8_211_0_clk;
 wire clknet_8_212_0_clk;
 wire clknet_8_213_0_clk;
 wire clknet_8_214_0_clk;
 wire clknet_8_215_0_clk;
 wire clknet_8_216_0_clk;
 wire clknet_8_217_0_clk;
 wire clknet_8_218_0_clk;
 wire clknet_8_219_0_clk;
 wire clknet_8_220_0_clk;
 wire clknet_8_221_0_clk;
 wire clknet_8_222_0_clk;
 wire clknet_8_223_0_clk;
 wire clknet_8_224_0_clk;
 wire clknet_8_225_0_clk;
 wire clknet_8_226_0_clk;
 wire clknet_8_227_0_clk;
 wire clknet_8_228_0_clk;
 wire clknet_8_229_0_clk;
 wire clknet_8_230_0_clk;
 wire clknet_8_231_0_clk;
 wire clknet_8_232_0_clk;
 wire clknet_8_233_0_clk;
 wire clknet_8_234_0_clk;
 wire clknet_8_235_0_clk;
 wire clknet_8_236_0_clk;
 wire clknet_8_237_0_clk;
 wire clknet_8_238_0_clk;
 wire clknet_8_239_0_clk;
 wire clknet_8_240_0_clk;
 wire clknet_8_241_0_clk;
 wire clknet_8_242_0_clk;
 wire clknet_8_243_0_clk;
 wire clknet_8_244_0_clk;
 wire clknet_8_245_0_clk;
 wire clknet_8_246_0_clk;
 wire clknet_8_247_0_clk;
 wire clknet_8_248_0_clk;
 wire clknet_8_249_0_clk;
 wire clknet_8_250_0_clk;
 wire clknet_8_251_0_clk;
 wire clknet_8_252_0_clk;
 wire clknet_8_253_0_clk;
 wire clknet_8_254_0_clk;
 wire clknet_8_255_0_clk;

 sg13g2_buf_16 clkbuf_leaf_832_clk (.X(clknet_leaf_832_clk),
    .A(clknet_8_175_0_clk));
 sg13g2_inv_4 _14114_ (.A(_00085_),
    .Y(_07697_));
 sg13g2_buf_16 clkbuf_leaf_831_clk (.X(clknet_leaf_831_clk),
    .A(clknet_8_175_0_clk));
 sg13g2_nand2b_1 _14116_ (.Y(_07699_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_state[0] ),
    .A_N(_00087_));
 sg13g2_buf_16 clkbuf_leaf_829_clk (.X(clknet_leaf_829_clk),
    .A(clknet_8_174_0_clk));
 sg13g2_inv_8 _14118_ (.Y(_07701_),
    .A(net10606));
 sg13g2_buf_16 clkbuf_leaf_828_clk (.X(clknet_leaf_828_clk),
    .A(clknet_8_174_0_clk));
 sg13g2_buf_16 clkbuf_leaf_824_clk (.X(clknet_leaf_824_clk),
    .A(clknet_8_171_0_clk));
 sg13g2_buf_16 clkbuf_leaf_823_clk (.X(clknet_leaf_823_clk),
    .A(clknet_8_170_0_clk));
 sg13g2_or3_1 _14122_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_do_rinst ),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_do_rdata ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_do_wdata ),
    .X(_07705_));
 sg13g2_buf_16 clkbuf_leaf_821_clk (.X(clknet_leaf_821_clk),
    .A(clknet_8_170_0_clk));
 sg13g2_inv_4 _14124_ (.A(net10617),
    .Y(_07707_));
 sg13g2_buf_16 clkbuf_leaf_820_clk (.X(clknet_leaf_820_clk),
    .A(clknet_8_170_0_clk));
 sg13g2_buf_16 clkbuf_leaf_817_clk (.X(clknet_leaf_817_clk),
    .A(clknet_8_184_0_clk));
 sg13g2_nor4_2 _14127_ (.A(\u_ac_controller_soc_inst.cbus_addr[27] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[26] ),
    .C(\u_ac_controller_soc_inst.cbus_addr[25] ),
    .Y(_07710_),
    .D(\u_ac_controller_soc_inst.cbus_addr[24] ));
 sg13g2_buf_16 clkbuf_leaf_816_clk (.X(clknet_leaf_816_clk),
    .A(clknet_8_184_0_clk));
 sg13g2_buf_16 clkbuf_leaf_815_clk (.X(clknet_leaf_815_clk),
    .A(clknet_8_178_0_clk));
 sg13g2_buf_16 clkbuf_leaf_814_clk (.X(clknet_leaf_814_clk),
    .A(clknet_8_184_0_clk));
 sg13g2_nor2_2 _14131_ (.A(\u_ac_controller_soc_inst.cbus_addr[28] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[29] ),
    .Y(_07714_));
 sg13g2_buf_16 clkbuf_leaf_813_clk (.X(clknet_leaf_813_clk),
    .A(clknet_8_184_0_clk));
 sg13g2_buf_16 clkbuf_leaf_811_clk (.X(clknet_leaf_811_clk),
    .A(clknet_8_186_0_clk));
 sg13g2_buf_16 clkbuf_leaf_810_clk (.X(clknet_leaf_810_clk),
    .A(clknet_8_186_0_clk));
 sg13g2_nor2_2 _14135_ (.A(\u_ac_controller_soc_inst.cbus_addr[30] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[31] ),
    .Y(_07718_));
 sg13g2_buf_16 clkbuf_leaf_808_clk (.X(clknet_leaf_808_clk),
    .A(clknet_8_186_0_clk));
 sg13g2_nand3_1 _14137_ (.B(_07714_),
    .C(_07718_),
    .A(_07710_),
    .Y(_07720_));
 sg13g2_buf_16 clkbuf_leaf_807_clk (.X(clknet_leaf_807_clk),
    .A(clknet_8_185_0_clk));
 sg13g2_buf_16 clkbuf_leaf_806_clk (.X(clknet_leaf_806_clk),
    .A(clknet_8_187_0_clk));
 sg13g2_buf_16 clkbuf_leaf_803_clk (.X(clknet_leaf_803_clk),
    .A(clknet_8_190_0_clk));
 sg13g2_o21ai_1 _14141_ (.B1(net10477),
    .Y(_07724_),
    .A1(_07707_),
    .A2(net10299));
 sg13g2_buf_16 clkbuf_leaf_801_clk (.X(clknet_leaf_801_clk),
    .A(clknet_8_187_0_clk));
 sg13g2_buf_16 clkbuf_leaf_800_clk (.X(clknet_leaf_800_clk),
    .A(clknet_8_185_0_clk));
 sg13g2_nand4_1 _14144_ (.B(_07710_),
    .C(_07714_),
    .A(\u_ac_controller_soc_inst.cbus_addr[16] ),
    .Y(_07727_),
    .D(_07718_));
 sg13g2_buf_16 clkbuf_leaf_799_clk (.X(clknet_leaf_799_clk),
    .A(clknet_8_188_0_clk));
 sg13g2_nand4_1 _14146_ (.B(_07710_),
    .C(_07714_),
    .A(\u_ac_controller_soc_inst.cbus_addr[14] ),
    .Y(_07729_),
    .D(_07718_));
 sg13g2_buf_16 clkbuf_leaf_798_clk (.X(clknet_leaf_798_clk),
    .A(clknet_8_177_0_clk));
 sg13g2_buf_16 clkbuf_leaf_797_clk (.X(clknet_leaf_797_clk),
    .A(clknet_8_177_0_clk));
 sg13g2_a22oi_1 _14149_ (.Y(_07732_),
    .B1(_07729_),
    .B2(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[14] ),
    .A2(_07727_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[16] ));
 sg13g2_and2_1 _14150_ (.A(_07724_),
    .B(_07732_),
    .X(_07733_));
 sg13g2_buf_16 clkbuf_leaf_795_clk (.X(clknet_leaf_795_clk),
    .A(clknet_8_179_0_clk));
 sg13g2_inv_1 _14152_ (.Y(_07735_),
    .A(\u_ac_controller_soc_inst.cbus_addr[22] ));
 sg13g2_buf_16 clkbuf_leaf_794_clk (.X(clknet_leaf_794_clk),
    .A(clknet_8_185_0_clk));
 sg13g2_o21ai_1 _14154_ (.B1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[22] ),
    .Y(_07737_),
    .A1(_07735_),
    .A2(_07720_));
 sg13g2_buf_16 clkbuf_leaf_793_clk (.X(clknet_leaf_793_clk),
    .A(clknet_8_178_0_clk));
 sg13g2_inv_2 _14156_ (.Y(_07739_),
    .A(\u_ac_controller_soc_inst.cbus_addr[12] ));
 sg13g2_buf_16 clkbuf_leaf_792_clk (.X(clknet_leaf_792_clk),
    .A(clknet_8_178_0_clk));
 sg13g2_o21ai_1 _14158_ (.B1(net10483),
    .Y(_07741_),
    .A1(_07739_),
    .A2(_07720_));
 sg13g2_inv_2 _14159_ (.Y(_07742_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_valid ));
 sg13g2_buf_16 clkbuf_leaf_791_clk (.X(clknet_leaf_791_clk),
    .A(clknet_8_174_0_clk));
 sg13g2_nand4_1 _14161_ (.B(_07710_),
    .C(_07714_),
    .A(\u_ac_controller_soc_inst.cbus_valid ),
    .Y(_07744_),
    .D(_07718_));
 sg13g2_buf_16 clkbuf_leaf_790_clk (.X(clknet_leaf_790_clk),
    .A(clknet_8_178_0_clk));
 sg13g2_nand2b_2 _14163_ (.Y(_07746_),
    .B(\u_ac_controller_soc_inst.cbus_addr[12] ),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[12] ));
 sg13g2_nand2b_1 _14164_ (.Y(_07747_),
    .B(\u_ac_controller_soc_inst.cbus_addr[14] ),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[14] ));
 sg13g2_nand2b_1 _14165_ (.Y(_07748_),
    .B(\u_ac_controller_soc_inst.cbus_addr[4] ),
    .A_N(net10477));
 sg13g2_nand3_1 _14166_ (.B(_07747_),
    .C(_07748_),
    .A(_07746_),
    .Y(_07749_));
 sg13g2_nand2b_1 _14167_ (.Y(_07750_),
    .B(\u_ac_controller_soc_inst.cbus_addr[22] ),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[22] ));
 sg13g2_nand2b_1 _14168_ (.Y(_07751_),
    .B(\u_ac_controller_soc_inst.cbus_addr[16] ),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[16] ));
 sg13g2_buf_16 clkbuf_leaf_789_clk (.X(clknet_leaf_789_clk),
    .A(clknet_8_179_0_clk));
 sg13g2_buf_16 clkbuf_leaf_788_clk (.X(clknet_leaf_788_clk),
    .A(clknet_8_179_0_clk));
 sg13g2_xnor2_1 _14171_ (.Y(_07754_),
    .A(\u_ac_controller_soc_inst.cbus_addr[6] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[6] ));
 sg13g2_buf_16 clkbuf_leaf_787_clk (.X(clknet_leaf_787_clk),
    .A(clknet_8_179_0_clk));
 sg13g2_buf_16 clkbuf_leaf_786_clk (.X(clknet_leaf_786_clk),
    .A(clknet_8_176_0_clk));
 sg13g2_nand2b_1 _14174_ (.Y(_07757_),
    .B(\u_ac_controller_soc_inst.cbus_addr[18] ),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[18] ));
 sg13g2_nand4_1 _14175_ (.B(_07751_),
    .C(_07754_),
    .A(_07750_),
    .Y(_07758_),
    .D(_07757_));
 sg13g2_nor4_1 _14176_ (.A(_07742_),
    .B(_07744_),
    .C(_07749_),
    .D(_07758_),
    .Y(_07759_));
 sg13g2_inv_4 _14177_ (.A(\u_ac_controller_soc_inst.cbus_addr[18] ),
    .Y(_07760_));
 sg13g2_o21ai_1 _14178_ (.B1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[18] ),
    .Y(_07761_),
    .A1(_07760_),
    .A2(net10299));
 sg13g2_and4_1 _14179_ (.A(_07737_),
    .B(_07741_),
    .C(_07759_),
    .D(_07761_),
    .X(_07762_));
 sg13g2_buf_16 clkbuf_leaf_781_clk (.X(clknet_leaf_781_clk),
    .A(clknet_8_176_0_clk));
 sg13g2_buf_16 clkbuf_leaf_780_clk (.X(clknet_leaf_780_clk),
    .A(clknet_8_173_0_clk));
 sg13g2_buf_16 clkbuf_leaf_778_clk (.X(clknet_leaf_778_clk),
    .A(clknet_8_180_0_clk));
 sg13g2_buf_16 clkbuf_leaf_777_clk (.X(clknet_leaf_777_clk),
    .A(clknet_8_181_0_clk));
 sg13g2_xnor2_1 _14184_ (.Y(_07767_),
    .A(net10622),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23] ));
 sg13g2_and3_1 _14185_ (.X(_07768_),
    .A(\u_ac_controller_soc_inst.cbus_addr[8] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[8] ),
    .C(_07767_));
 sg13g2_inv_1 _14186_ (.Y(_07769_),
    .A(net10622));
 sg13g2_inv_1 _14187_ (.Y(_07770_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23] ));
 sg13g2_nor4_1 _14188_ (.A(\u_ac_controller_soc_inst.cbus_addr[8] ),
    .B(_07769_),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[8] ),
    .D(_07770_),
    .Y(_07771_));
 sg13g2_or4_1 _14189_ (.A(\u_ac_controller_soc_inst.cbus_addr[27] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[26] ),
    .C(\u_ac_controller_soc_inst.cbus_addr[25] ),
    .D(\u_ac_controller_soc_inst.cbus_addr[24] ),
    .X(_07772_));
 sg13g2_or2_1 _14190_ (.X(_07773_),
    .B(\u_ac_controller_soc_inst.cbus_addr[31] ),
    .A(\u_ac_controller_soc_inst.cbus_addr[30] ));
 sg13g2_nor4_2 _14191_ (.A(\u_ac_controller_soc_inst.cbus_addr[28] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[29] ),
    .C(_07772_),
    .Y(_07774_),
    .D(_07773_));
 sg13g2_buf_16 clkbuf_leaf_776_clk (.X(clknet_leaf_776_clk),
    .A(clknet_8_180_0_clk));
 sg13g2_o21ai_1 _14193_ (.B1(net10295),
    .Y(_07776_),
    .A1(_07768_),
    .A2(_07771_));
 sg13g2_nor2_1 _14194_ (.A(\u_ac_controller_soc_inst.cbus_addr[8] ),
    .B(net10622),
    .Y(_07777_));
 sg13g2_buf_16 clkbuf_leaf_775_clk (.X(clknet_leaf_775_clk),
    .A(clknet_8_180_0_clk));
 sg13g2_nor2_1 _14196_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[8] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23] ),
    .Y(_07779_));
 sg13g2_o21ai_1 _14197_ (.B1(_07779_),
    .Y(_07780_),
    .A1(net10300),
    .A2(_07777_));
 sg13g2_buf_16 clkbuf_leaf_774_clk (.X(clknet_leaf_774_clk),
    .A(clknet_8_177_0_clk));
 sg13g2_buf_16 clkbuf_leaf_773_clk (.X(clknet_leaf_773_clk),
    .A(clknet_8_180_0_clk));
 sg13g2_buf_16 clkbuf_leaf_772_clk (.X(clknet_leaf_772_clk),
    .A(clknet_8_183_0_clk));
 sg13g2_buf_16 clkbuf_leaf_771_clk (.X(clknet_leaf_771_clk),
    .A(clknet_8_181_0_clk));
 sg13g2_xnor2_1 _14202_ (.Y(_07785_),
    .A(\u_ac_controller_soc_inst.cbus_addr[10] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[10] ));
 sg13g2_and3_1 _14203_ (.X(_07786_),
    .A(\u_ac_controller_soc_inst.cbus_addr[17] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[17] ),
    .C(_07785_));
 sg13g2_inv_1 _14204_ (.Y(_07787_),
    .A(\u_ac_controller_soc_inst.cbus_addr[10] ));
 sg13g2_inv_4 _14205_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[10] ),
    .Y(_07788_));
 sg13g2_nor4_1 _14206_ (.A(\u_ac_controller_soc_inst.cbus_addr[17] ),
    .B(_07787_),
    .C(_07788_),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[17] ),
    .Y(_07789_));
 sg13g2_o21ai_1 _14207_ (.B1(net10295),
    .Y(_07790_),
    .A1(_07786_),
    .A2(_07789_));
 sg13g2_nor2_1 _14208_ (.A(\u_ac_controller_soc_inst.cbus_addr[17] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[10] ),
    .Y(_07791_));
 sg13g2_nor2_1 _14209_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[10] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[17] ),
    .Y(_07792_));
 sg13g2_o21ai_1 _14210_ (.B1(_07792_),
    .Y(_07793_),
    .A1(net10300),
    .A2(_07791_));
 sg13g2_a22oi_1 _14211_ (.Y(_07794_),
    .B1(_07790_),
    .B2(_07793_),
    .A2(_07780_),
    .A1(_07776_));
 sg13g2_buf_16 clkbuf_leaf_770_clk (.X(clknet_leaf_770_clk),
    .A(clknet_8_183_0_clk));
 sg13g2_buf_16 clkbuf_leaf_769_clk (.X(clknet_leaf_769_clk),
    .A(clknet_8_233_0_clk));
 sg13g2_buf_16 clkbuf_leaf_768_clk (.X(clknet_leaf_768_clk),
    .A(clknet_8_233_0_clk));
 sg13g2_buf_16 clkbuf_leaf_767_clk (.X(clknet_leaf_767_clk),
    .A(clknet_8_183_0_clk));
 sg13g2_buf_16 clkbuf_leaf_765_clk (.X(clknet_leaf_765_clk),
    .A(clknet_8_183_0_clk));
 sg13g2_xnor2_1 _14217_ (.Y(_07800_),
    .A(net10625),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[13] ));
 sg13g2_and3_1 _14218_ (.X(_07801_),
    .A(net10619),
    .B(net10478),
    .C(_07800_));
 sg13g2_nand3b_1 _14219_ (.B(net10625),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[13] ),
    .Y(_07802_),
    .A_N(net10619));
 sg13g2_nor2_1 _14220_ (.A(net10478),
    .B(_07802_),
    .Y(_07803_));
 sg13g2_o21ai_1 _14221_ (.B1(net10295),
    .Y(_07804_),
    .A1(_07801_),
    .A2(_07803_));
 sg13g2_nor2_1 _14222_ (.A(\u_ac_controller_soc_inst.cbus_addr[3] ),
    .B(net10625),
    .Y(_07805_));
 sg13g2_nor2_1 _14223_ (.A(net10478),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[13] ),
    .Y(_07806_));
 sg13g2_o21ai_1 _14224_ (.B1(_07806_),
    .Y(_07807_),
    .A1(net10299),
    .A2(_07805_));
 sg13g2_buf_16 clkbuf_leaf_759_clk (.X(clknet_leaf_759_clk),
    .A(clknet_8_182_0_clk));
 sg13g2_buf_16 clkbuf_leaf_758_clk (.X(clknet_leaf_758_clk),
    .A(clknet_8_188_0_clk));
 sg13g2_nand4_1 _14227_ (.B(_07710_),
    .C(_07714_),
    .A(\u_ac_controller_soc_inst.cbus_addr[7] ),
    .Y(_07810_),
    .D(_07718_));
 sg13g2_xnor2_1 _14228_ (.Y(_07811_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[7] ),
    .B(_07810_));
 sg13g2_a21oi_1 _14229_ (.A1(_07804_),
    .A2(_07807_),
    .Y(_07812_),
    .B1(_07811_));
 sg13g2_nand4_1 _14230_ (.B(_07762_),
    .C(_07794_),
    .A(_07733_),
    .Y(_07813_),
    .D(_07812_));
 sg13g2_buf_16 clkbuf_leaf_757_clk (.X(clknet_leaf_757_clk),
    .A(clknet_8_188_0_clk));
 sg13g2_buf_16 clkbuf_leaf_755_clk (.X(clknet_leaf_755_clk),
    .A(clknet_8_190_0_clk));
 sg13g2_buf_16 clkbuf_leaf_754_clk (.X(clknet_leaf_754_clk),
    .A(clknet_8_190_0_clk));
 sg13g2_buf_16 clkbuf_leaf_753_clk (.X(clknet_leaf_753_clk),
    .A(clknet_8_190_0_clk));
 sg13g2_buf_16 clkbuf_leaf_752_clk (.X(clknet_leaf_752_clk),
    .A(clknet_8_190_0_clk));
 sg13g2_xnor2_1 _14236_ (.Y(_07819_),
    .A(\u_ac_controller_soc_inst.cbus_addr[19] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19] ));
 sg13g2_and3_1 _14237_ (.X(_07820_),
    .A(\u_ac_controller_soc_inst.cbus_addr[2] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2] ),
    .C(_07819_));
 sg13g2_nand3b_1 _14238_ (.B(\u_ac_controller_soc_inst.cbus_addr[19] ),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19] ),
    .Y(_07821_),
    .A_N(\u_ac_controller_soc_inst.cbus_addr[2] ));
 sg13g2_nor2_1 _14239_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2] ),
    .B(_07821_),
    .Y(_07822_));
 sg13g2_o21ai_1 _14240_ (.B1(_07774_),
    .Y(_07823_),
    .A1(_07820_),
    .A2(_07822_));
 sg13g2_nor2_1 _14241_ (.A(\u_ac_controller_soc_inst.cbus_addr[2] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[19] ),
    .Y(_07824_));
 sg13g2_nor2_1 _14242_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19] ),
    .Y(_07825_));
 sg13g2_o21ai_1 _14243_ (.B1(_07825_),
    .Y(_07826_),
    .A1(net10299),
    .A2(_07824_));
 sg13g2_nand2_1 _14244_ (.Y(_07827_),
    .A(_07823_),
    .B(_07826_));
 sg13g2_buf_16 clkbuf_leaf_750_clk (.X(clknet_leaf_750_clk),
    .A(clknet_8_191_0_clk));
 sg13g2_buf_16 clkbuf_leaf_749_clk (.X(clknet_leaf_749_clk),
    .A(clknet_8_191_0_clk));
 sg13g2_xnor2_1 _14247_ (.Y(_07830_),
    .A(net10626),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[11] ));
 sg13g2_buf_16 clkbuf_leaf_748_clk (.X(clknet_leaf_748_clk),
    .A(clknet_8_191_0_clk));
 sg13g2_buf_16 clkbuf_leaf_747_clk (.X(clknet_leaf_747_clk),
    .A(clknet_8_234_0_clk));
 sg13g2_and2_1 _14250_ (.A(\u_ac_controller_soc_inst.cbus_addr[15] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15] ),
    .X(_07833_));
 sg13g2_nor2b_1 _14251_ (.A(\u_ac_controller_soc_inst.cbus_addr[15] ),
    .B_N(net10626),
    .Y(_07834_));
 sg13g2_nor2b_1 _14252_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15] ),
    .B_N(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[11] ),
    .Y(_07835_));
 sg13g2_a22oi_1 _14253_ (.Y(_07836_),
    .B1(_07834_),
    .B2(_07835_),
    .A2(_07833_),
    .A1(_07830_));
 sg13g2_nor2_1 _14254_ (.A(\u_ac_controller_soc_inst.cbus_addr[15] ),
    .B(net10626),
    .Y(_07837_));
 sg13g2_buf_16 clkbuf_leaf_744_clk (.X(clknet_leaf_744_clk),
    .A(clknet_8_189_0_clk));
 sg13g2_nor2_1 _14256_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[11] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15] ),
    .Y(_07839_));
 sg13g2_o21ai_1 _14257_ (.B1(_07839_),
    .Y(_07840_),
    .A1(net10299),
    .A2(_07837_));
 sg13g2_o21ai_1 _14258_ (.B1(_07840_),
    .Y(_07841_),
    .A1(net10299),
    .A2(_07836_));
 sg13g2_buf_16 clkbuf_leaf_743_clk (.X(clknet_leaf_743_clk),
    .A(clknet_8_189_0_clk));
 sg13g2_buf_16 clkbuf_leaf_742_clk (.X(clknet_leaf_742_clk),
    .A(clknet_8_232_0_clk));
 sg13g2_buf_16 clkbuf_leaf_740_clk (.X(clknet_leaf_740_clk),
    .A(clknet_8_238_0_clk));
 sg13g2_buf_16 clkbuf_leaf_739_clk (.X(clknet_leaf_739_clk),
    .A(clknet_8_232_0_clk));
 sg13g2_xnor2_1 _14263_ (.Y(_07846_),
    .A(net10624),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20] ));
 sg13g2_and3_1 _14264_ (.X(_07847_),
    .A(net10616),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[5] ),
    .C(_07846_));
 sg13g2_buf_16 clkbuf_leaf_738_clk (.X(clknet_leaf_738_clk),
    .A(clknet_8_238_0_clk));
 sg13g2_nand3b_1 _14266_ (.B(net10624),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20] ),
    .Y(_07849_),
    .A_N(net10616));
 sg13g2_nor2_1 _14267_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[5] ),
    .B(_07849_),
    .Y(_07850_));
 sg13g2_o21ai_1 _14268_ (.B1(_07774_),
    .Y(_07851_),
    .A1(_07847_),
    .A2(_07850_));
 sg13g2_nor2_1 _14269_ (.A(\u_ac_controller_soc_inst.cbus_addr[5] ),
    .B(net10624),
    .Y(_07852_));
 sg13g2_nor2_1 _14270_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[5] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20] ),
    .Y(_07853_));
 sg13g2_o21ai_1 _14271_ (.B1(_07853_),
    .Y(_07854_),
    .A1(_07720_),
    .A2(_07852_));
 sg13g2_nand2_1 _14272_ (.Y(_07855_),
    .A(_07851_),
    .B(_07854_));
 sg13g2_buf_16 clkbuf_leaf_736_clk (.X(clknet_leaf_736_clk),
    .A(clknet_8_234_0_clk));
 sg13g2_buf_16 clkbuf_leaf_734_clk (.X(clknet_leaf_734_clk),
    .A(clknet_8_234_0_clk));
 sg13g2_buf_16 clkbuf_leaf_733_clk (.X(clknet_leaf_733_clk),
    .A(clknet_8_235_0_clk));
 sg13g2_buf_16 clkbuf_leaf_731_clk (.X(clknet_leaf_731_clk),
    .A(clknet_8_235_0_clk));
 sg13g2_xnor2_1 _14277_ (.Y(_07860_),
    .A(net10623),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21] ));
 sg13g2_nand3_1 _14278_ (.B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[9] ),
    .C(_07860_),
    .A(\u_ac_controller_soc_inst.cbus_addr[9] ),
    .Y(_07861_));
 sg13g2_nor2_1 _14279_ (.A(\u_ac_controller_soc_inst.cbus_addr[9] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[9] ),
    .Y(_07862_));
 sg13g2_nand3_1 _14280_ (.B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21] ),
    .C(_07862_),
    .A(net10623),
    .Y(_07863_));
 sg13g2_and2_1 _14281_ (.A(_07861_),
    .B(_07863_),
    .X(_07864_));
 sg13g2_nor2_1 _14282_ (.A(\u_ac_controller_soc_inst.cbus_addr[9] ),
    .B(net10623),
    .Y(_07865_));
 sg13g2_nor2_1 _14283_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[9] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21] ),
    .Y(_07866_));
 sg13g2_o21ai_1 _14284_ (.B1(_07866_),
    .Y(_07867_),
    .A1(net10299),
    .A2(_07865_));
 sg13g2_o21ai_1 _14285_ (.B1(_07867_),
    .Y(_07868_),
    .A1(net10299),
    .A2(_07864_));
 sg13g2_nand4_1 _14286_ (.B(_07841_),
    .C(_07855_),
    .A(_07827_),
    .Y(_07869_),
    .D(_07868_));
 sg13g2_nor2_1 _14287_ (.A(\u_ac_controller_soc_inst.cbus_addr[23] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[22] ),
    .Y(_07870_));
 sg13g2_nor4_1 _14288_ (.A(\u_ac_controller_soc_inst.cbus_addr[21] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[20] ),
    .C(\u_ac_controller_soc_inst.cbus_addr[19] ),
    .D(\u_ac_controller_soc_inst.cbus_addr[18] ),
    .Y(_07871_));
 sg13g2_nand4_1 _14289_ (.B(_07718_),
    .C(_07870_),
    .A(_07710_),
    .Y(_07872_),
    .D(_07871_));
 sg13g2_buf_16 clkbuf_leaf_730_clk (.X(clknet_leaf_730_clk),
    .A(clknet_8_239_0_clk));
 sg13g2_or2_1 _14291_ (.X(_07874_),
    .B(\u_ac_controller_soc_inst.cbus_addr[16] ),
    .A(\u_ac_controller_soc_inst.cbus_addr[17] ));
 sg13g2_buf_16 clkbuf_leaf_728_clk (.X(clknet_leaf_728_clk),
    .A(clknet_8_239_0_clk));
 sg13g2_or4_1 _14293_ (.A(\u_ac_controller_soc_inst.cbus_addr[9] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[15] ),
    .C(\u_ac_controller_soc_inst.cbus_addr[12] ),
    .D(\u_ac_controller_soc_inst.cbus_addr[11] ),
    .X(_07876_));
 sg13g2_buf_16 clkbuf_leaf_727_clk (.X(clknet_leaf_727_clk),
    .A(clknet_8_239_0_clk));
 sg13g2_or3_1 _14295_ (.A(\u_ac_controller_soc_inst.cbus_addr[14] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[13] ),
    .C(\u_ac_controller_soc_inst.cbus_addr[10] ),
    .X(_07878_));
 sg13g2_buf_16 clkbuf_leaf_726_clk (.X(clknet_leaf_726_clk),
    .A(clknet_8_239_0_clk));
 sg13g2_or3_1 _14297_ (.A(_07874_),
    .B(_07876_),
    .C(_07878_),
    .X(_07880_));
 sg13g2_nor2_2 _14298_ (.A(\u_ac_controller_soc_inst.cbus_addr[7] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[6] ),
    .Y(_07881_));
 sg13g2_nor4_2 _14299_ (.A(\u_ac_controller_soc_inst.cbus_addr[3] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[2] ),
    .C(\u_ac_controller_soc_inst.cbus_addr[5] ),
    .Y(_07882_),
    .D(\u_ac_controller_soc_inst.cbus_addr[4] ));
 sg13g2_inv_1 _14300_ (.Y(_07883_),
    .A(\u_ac_controller_soc_inst.cbus_addr[8] ));
 sg13g2_a21oi_2 _14301_ (.B1(_07883_),
    .Y(_07884_),
    .A2(_07882_),
    .A1(_07881_));
 sg13g2_nand2b_1 _14302_ (.Y(_07885_),
    .B(\u_ac_controller_soc_inst.cbus_addr[29] ),
    .A_N(\u_ac_controller_soc_inst.cbus_addr[28] ));
 sg13g2_nor4_2 _14303_ (.A(_07872_),
    .B(_07880_),
    .C(_07884_),
    .Y(_07886_),
    .D(_07885_));
 sg13g2_and2_1 _14304_ (.A(\u_ac_controller_soc_inst.cbus_valid ),
    .B(_07886_),
    .X(_07887_));
 sg13g2_buf_16 clkbuf_leaf_725_clk (.X(clknet_leaf_725_clk),
    .A(clknet_8_236_0_clk));
 sg13g2_inv_1 _14306_ (.Y(_07889_),
    .A(\u_ac_controller_soc_inst.io_ready ));
 sg13g2_or2_1 _14307_ (.X(_07890_),
    .B(\u_ac_controller_soc_inst.cbus_addr[22] ),
    .A(net10622));
 sg13g2_buf_16 clkbuf_leaf_724_clk (.X(clknet_leaf_724_clk),
    .A(clknet_8_236_0_clk));
 sg13g2_or4_1 _14309_ (.A(net10623),
    .B(net10624),
    .C(\u_ac_controller_soc_inst.cbus_addr[19] ),
    .D(\u_ac_controller_soc_inst.cbus_addr[18] ),
    .X(_07892_));
 sg13g2_buf_16 clkbuf_leaf_723_clk (.X(clknet_leaf_723_clk),
    .A(clknet_8_236_0_clk));
 sg13g2_nor4_1 _14311_ (.A(_07772_),
    .B(_07773_),
    .C(_07890_),
    .D(_07892_),
    .Y(_07894_));
 sg13g2_nor4_2 _14312_ (.A(\u_ac_controller_soc_inst.cbus_addr[8] ),
    .B(_07874_),
    .C(_07876_),
    .Y(_07895_),
    .D(_07878_));
 sg13g2_buf_16 clkbuf_leaf_722_clk (.X(clknet_leaf_722_clk),
    .A(clknet_8_238_0_clk));
 sg13g2_nand4_1 _14314_ (.B(\u_ac_controller_soc_inst.cbus_addr[29] ),
    .C(_07894_),
    .A(\u_ac_controller_soc_inst.cbus_addr[28] ),
    .Y(_07897_),
    .D(_07895_));
 sg13g2_buf_16 clkbuf_leaf_721_clk (.X(clknet_leaf_721_clk),
    .A(clknet_8_238_0_clk));
 sg13g2_and2_1 _14316_ (.A(_07710_),
    .B(_07714_),
    .X(_07899_));
 sg13g2_buf_16 clkbuf_leaf_718_clk (.X(clknet_leaf_718_clk),
    .A(clknet_8_232_0_clk));
 sg13g2_nor2b_2 _14318_ (.A(\u_ac_controller_soc_inst.cbus_addr[31] ),
    .B_N(\u_ac_controller_soc_inst.cbus_addr[30] ),
    .Y(_07901_));
 sg13g2_and3_2 _14319_ (.X(_07902_),
    .A(_07870_),
    .B(_07871_),
    .C(_07901_));
 sg13g2_nand4_1 _14320_ (.B(_07899_),
    .C(_07895_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_ready ),
    .Y(_07903_),
    .D(_07902_));
 sg13g2_o21ai_1 _14321_ (.B1(_07903_),
    .Y(_07904_),
    .A1(_07889_),
    .A2(_07897_));
 sg13g2_inv_2 _14322_ (.Y(_07905_),
    .A(\u_ac_controller_soc_inst.cbus_valid ));
 sg13g2_nor3_1 _14323_ (.A(\u_ac_controller_soc_inst.cbus_addr[29] ),
    .B(_07905_),
    .C(_07874_),
    .Y(_07906_));
 sg13g2_and3_2 _14324_ (.X(_07907_),
    .A(\u_ac_controller_soc_inst.cbus_addr[28] ),
    .B(_07894_),
    .C(_07906_));
 sg13g2_buf_16 clkbuf_leaf_717_clk (.X(clknet_leaf_717_clk),
    .A(clknet_8_233_0_clk));
 sg13g2_and2_1 _14326_ (.A(\u_ac_controller_soc_inst.sram_ready ),
    .B(_07907_),
    .X(_07909_));
 sg13g2_a221oi_1 _14327_ (.B2(_07701_),
    .C1(_07909_),
    .B1(_07904_),
    .A1(\u_ac_controller_soc_inst.spi_sensor_ready ),
    .Y(_07910_),
    .A2(_07887_));
 sg13g2_o21ai_1 _14328_ (.B1(_07910_),
    .Y(_07911_),
    .A1(_07813_),
    .A2(_07869_));
 sg13g2_nand3_1 _14329_ (.B(_07705_),
    .C(_07911_),
    .A(_07701_),
    .Y(_07912_));
 sg13g2_buf_16 clkbuf_leaf_714_clk (.X(clknet_leaf_714_clk),
    .A(clknet_8_227_0_clk));
 sg13g2_inv_1 _14331_ (.Y(_07914_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_state[1] ));
 sg13g2_a21oi_2 _14332_ (.B1(_07914_),
    .Y(_07915_),
    .A2(_07912_),
    .A1(_07699_));
 sg13g2_inv_2 _14333_ (.Y(_07916_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_state[0] ));
 sg13g2_inv_1 _14334_ (.Y(_07917_),
    .A(_07705_));
 sg13g2_and3_1 _14335_ (.X(_07918_),
    .A(_07732_),
    .B(_07737_),
    .C(_07759_));
 sg13g2_and3_1 _14336_ (.X(_07919_),
    .A(_07724_),
    .B(_07741_),
    .C(_07761_));
 sg13g2_a21oi_1 _14337_ (.A1(_07823_),
    .A2(_07826_),
    .Y(_07920_),
    .B1(_07811_));
 sg13g2_a22oi_1 _14338_ (.Y(_07921_),
    .B1(_07851_),
    .B2(_07854_),
    .A2(_07807_),
    .A1(_07804_));
 sg13g2_and4_2 _14339_ (.A(_07918_),
    .B(_07919_),
    .C(_07920_),
    .D(_07921_),
    .X(_07922_));
 sg13g2_and3_2 _14340_ (.X(_07923_),
    .A(_07794_),
    .B(_07841_),
    .C(_07868_));
 sg13g2_and4_2 _14341_ (.A(\u_ac_controller_soc_inst.cbus_addr[28] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[29] ),
    .C(_07894_),
    .D(_07895_),
    .X(_07924_));
 sg13g2_buf_16 clkbuf_leaf_712_clk (.X(clknet_leaf_712_clk),
    .A(clknet_8_227_0_clk));
 sg13g2_nor2_2 _14343_ (.A(_07890_),
    .B(_07892_),
    .Y(_07926_));
 sg13g2_and4_2 _14344_ (.A(_07899_),
    .B(_07926_),
    .C(_07895_),
    .D(_07901_),
    .X(_07927_));
 sg13g2_buf_16 clkbuf_leaf_711_clk (.X(clknet_leaf_711_clk),
    .A(clknet_8_230_0_clk));
 sg13g2_a22oi_1 _14346_ (.Y(_07929_),
    .B1(_07927_),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_ready ),
    .A2(_07924_),
    .A1(\u_ac_controller_soc_inst.io_ready ));
 sg13g2_or4_1 _14347_ (.A(_07874_),
    .B(_07876_),
    .C(_07878_),
    .D(_07885_),
    .X(_07930_));
 sg13g2_nor4_2 _14348_ (.A(_07905_),
    .B(_07872_),
    .C(_07884_),
    .Y(_07931_),
    .D(_07930_));
 sg13g2_buf_16 clkbuf_leaf_708_clk (.X(clknet_leaf_708_clk),
    .A(clknet_8_230_0_clk));
 sg13g2_a22oi_1 _14350_ (.Y(_07933_),
    .B1(_07931_),
    .B2(\u_ac_controller_soc_inst.spi_sensor_ready ),
    .A2(_07907_),
    .A1(\u_ac_controller_soc_inst.sram_ready ));
 sg13g2_o21ai_1 _14351_ (.B1(_07933_),
    .Y(_07934_),
    .A1(net10606),
    .A2(_07929_));
 sg13g2_a21oi_2 _14352_ (.B1(_07934_),
    .Y(_07935_),
    .A2(_07923_),
    .A1(_07922_));
 sg13g2_or2_1 _14353_ (.X(_07936_),
    .B(_07935_),
    .A(_00086_));
 sg13g2_buf_16 clkbuf_leaf_707_clk (.X(clknet_leaf_707_clk),
    .A(clknet_8_230_0_clk));
 sg13g2_nor3_2 _14355_ (.A(_07916_),
    .B(_07917_),
    .C(_07936_),
    .Y(_07938_));
 sg13g2_buf_16 clkbuf_leaf_706_clk (.X(clknet_leaf_706_clk),
    .A(clknet_8_254_0_clk));
 sg13g2_o21ai_1 _14357_ (.B1(net11050),
    .Y(_07940_),
    .A1(_07915_),
    .A2(_07938_));
 sg13g2_buf_16 clkbuf_leaf_705_clk (.X(clknet_leaf_705_clk),
    .A(clknet_8_228_0_clk));
 sg13g2_and2_1 _14359_ (.A(_07697_),
    .B(_07940_),
    .X(_07942_));
 sg13g2_buf_16 clkbuf_leaf_704_clk (.X(clknet_leaf_704_clk),
    .A(clknet_8_231_0_clk));
 sg13g2_buf_16 clkbuf_leaf_703_clk (.X(clknet_leaf_703_clk),
    .A(clknet_8_254_0_clk));
 sg13g2_buf_16 clkbuf_leaf_701_clk (.X(clknet_leaf_701_clk),
    .A(clknet_8_254_0_clk));
 sg13g2_nand2b_2 _14363_ (.Y(_07946_),
    .B(net11050),
    .A_N(_07942_));
 sg13g2_or2_1 _14364_ (.X(_07947_),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_lhu ),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_lh ));
 sg13g2_buf_16 clkbuf_leaf_700_clk (.X(clknet_leaf_700_clk),
    .A(clknet_8_254_0_clk));
 sg13g2_inv_8 _14366_ (.Y(_07949_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[6] ));
 sg13g2_buf_16 clkbuf_leaf_699_clk (.X(clknet_leaf_699_clk),
    .A(clknet_8_251_0_clk));
 sg13g2_nor2_1 _14368_ (.A(net10610),
    .B(_07949_),
    .Y(_07951_));
 sg13g2_buf_16 clkbuf_leaf_698_clk (.X(clknet_leaf_698_clk),
    .A(clknet_8_224_0_clk));
 sg13g2_inv_2 _14370_ (.Y(_07953_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[5] ));
 sg13g2_nor2_2 _14371_ (.A(net10609),
    .B(_07953_),
    .Y(_07954_));
 sg13g2_a22oi_1 _14372_ (.Y(_07955_),
    .B1(_07954_),
    .B2(\u_ac_controller_soc_inst.u_picorv32.instr_sh ),
    .A2(_07951_),
    .A1(_07947_));
 sg13g2_nor2_2 _14373_ (.A(_07915_),
    .B(_07938_),
    .Y(_07956_));
 sg13g2_buf_16 clkbuf_leaf_697_clk (.X(clknet_leaf_697_clk),
    .A(clknet_8_225_0_clk));
 sg13g2_nor3_2 _14375_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_sh ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_sb ),
    .C(\u_ac_controller_soc_inst.u_picorv32.instr_sw ),
    .Y(_07958_));
 sg13g2_nor2_1 _14376_ (.A(net10609),
    .B(_00089_),
    .Y(_07959_));
 sg13g2_a22oi_1 _14377_ (.Y(_07960_),
    .B1(_07958_),
    .B2(_07959_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpu_state[5] ),
    .A1(net10609));
 sg13g2_or2_1 _14378_ (.X(_07961_),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_lbu ),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_lb ));
 sg13g2_nor3_2 _14379_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_lw ),
    .B(_07947_),
    .C(_07961_),
    .Y(_07962_));
 sg13g2_buf_16 clkbuf_leaf_696_clk (.X(clknet_leaf_696_clk),
    .A(clknet_8_226_0_clk));
 sg13g2_nor2_1 _14381_ (.A(net10610),
    .B(_00088_),
    .Y(_07964_));
 sg13g2_a22oi_1 _14382_ (.Y(_07965_),
    .B1(_07962_),
    .B2(_07964_),
    .A2(net10695),
    .A1(net10610));
 sg13g2_a22oi_1 _14383_ (.Y(_07966_),
    .B1(_07960_),
    .B2(_07965_),
    .A2(_07956_),
    .A1(_07697_));
 sg13g2_nand2_2 _14384_ (.Y(_07967_),
    .A(_07697_),
    .B(_07956_));
 sg13g2_nand2_1 _14385_ (.Y(_07968_),
    .A(_00088_),
    .B(_00089_));
 sg13g2_inv_1 _14386_ (.Y(_07969_),
    .A(_07968_));
 sg13g2_nor2_1 _14387_ (.A(_07967_),
    .B(_07969_),
    .Y(_07970_));
 sg13g2_buf_16 clkbuf_leaf_695_clk (.X(clknet_leaf_695_clk),
    .A(clknet_8_226_0_clk));
 sg13g2_nand2_2 _14389_ (.Y(_07972_),
    .A(_07949_),
    .B(_07953_));
 sg13g2_o21ai_1 _14390_ (.B1(net11050),
    .Y(_07973_),
    .A1(net10722),
    .A2(_07972_));
 sg13g2_nor3_2 _14391_ (.A(_07966_),
    .B(_07970_),
    .C(_07973_),
    .Y(_07974_));
 sg13g2_buf_16 clkbuf_leaf_694_clk (.X(clknet_leaf_694_clk),
    .A(clknet_8_233_0_clk));
 sg13g2_buf_16 clkbuf_leaf_693_clk (.X(clknet_leaf_693_clk),
    .A(clknet_8_226_0_clk));
 sg13g2_nand2b_1 _14394_ (.Y(_07977_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[2] ),
    .A_N(_07974_));
 sg13g2_o21ai_1 _14395_ (.B1(_07977_),
    .Y(_00019_),
    .A1(_07946_),
    .A2(_07955_));
 sg13g2_buf_16 clkbuf_leaf_692_clk (.X(clknet_leaf_692_clk),
    .A(clknet_8_226_0_clk));
 sg13g2_nor2_2 _14397_ (.A(_07905_),
    .B(_07720_),
    .Y(_07979_));
 sg13g2_buf_16 clkbuf_leaf_690_clk (.X(clknet_leaf_690_clk),
    .A(clknet_8_225_0_clk));
 sg13g2_buf_16 clkbuf_leaf_689_clk (.X(clknet_leaf_689_clk),
    .A(clknet_8_225_0_clk));
 sg13g2_o21ai_1 _14400_ (.B1(_07979_),
    .Y(_07982_),
    .A1(_07813_),
    .A2(_07869_));
 sg13g2_buf_16 clkbuf_leaf_688_clk (.X(clknet_leaf_688_clk),
    .A(clknet_8_225_0_clk));
 sg13g2_buf_16 clkbuf_leaf_687_clk (.X(clknet_leaf_687_clk),
    .A(clknet_8_224_0_clk));
 sg13g2_buf_16 clkbuf_leaf_685_clk (.X(clknet_leaf_685_clk),
    .A(clknet_8_181_0_clk));
 sg13g2_inv_1 _14404_ (.Y(_07986_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[17] ));
 sg13g2_nand2_1 _14405_ (.Y(_07987_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[16] ));
 sg13g2_and4_2 _14406_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[10] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[11] ),
    .C(net10483),
    .D(net10482),
    .X(_07988_));
 sg13g2_nand2_2 _14407_ (.Y(_07989_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[14] ),
    .B(_07988_));
 sg13g2_nand3_1 _14408_ (.B(net10478),
    .C(net10477),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2] ),
    .Y(_07990_));
 sg13g2_buf_16 clkbuf_leaf_684_clk (.X(clknet_leaf_684_clk),
    .A(clknet_8_224_0_clk));
 sg13g2_nand3_1 _14410_ (.B(net10475),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[7] ),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[5] ),
    .Y(_07992_));
 sg13g2_buf_16 clkbuf_leaf_682_clk (.X(clknet_leaf_682_clk),
    .A(clknet_8_172_0_clk));
 sg13g2_nor2_2 _14412_ (.A(_07990_),
    .B(_07992_),
    .Y(_07994_));
 sg13g2_buf_16 clkbuf_leaf_681_clk (.X(clknet_leaf_681_clk),
    .A(clknet_8_251_0_clk));
 sg13g2_nand3_1 _14414_ (.B(net10473),
    .C(_07994_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[8] ),
    .Y(_07996_));
 sg13g2_buf_16 clkbuf_leaf_680_clk (.X(clknet_leaf_680_clk),
    .A(clknet_8_251_0_clk));
 sg13g2_nor4_2 _14416_ (.A(_07986_),
    .B(_07987_),
    .C(_07989_),
    .Y(_07998_),
    .D(_07996_));
 sg13g2_buf_16 clkbuf_leaf_679_clk (.X(clknet_leaf_679_clk),
    .A(clknet_8_250_0_clk));
 sg13g2_and4_2 _14418_ (.A(net10481),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19] ),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20] ),
    .D(_07998_),
    .X(_08000_));
 sg13g2_buf_16 clkbuf_leaf_678_clk (.X(clknet_leaf_678_clk),
    .A(clknet_8_251_0_clk));
 sg13g2_and2_1 _14420_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21] ),
    .B(_08000_),
    .X(_08002_));
 sg13g2_buf_16 clkbuf_leaf_677_clk (.X(clknet_leaf_677_clk),
    .A(clknet_8_224_0_clk));
 sg13g2_or3_1 _14422_ (.A(net10480),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23] ),
    .C(_08002_),
    .X(_08004_));
 sg13g2_and4_1 _14423_ (.A(net10481),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19] ),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20] ),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21] ),
    .X(_08005_));
 sg13g2_nor3_1 _14424_ (.A(_07987_),
    .B(_07989_),
    .C(_07996_),
    .Y(_08006_));
 sg13g2_and2_1 _14425_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[17] ),
    .B(_08006_),
    .X(_08007_));
 sg13g2_buf_16 clkbuf_leaf_676_clk (.X(clknet_leaf_676_clk),
    .A(clknet_8_250_0_clk));
 sg13g2_nand4_1 _14427_ (.B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23] ),
    .C(_08005_),
    .A(net10480),
    .Y(_08009_),
    .D(_08007_));
 sg13g2_a22oi_1 _14428_ (.Y(_08010_),
    .B1(_08004_),
    .B2(_08009_),
    .A2(_07890_),
    .A1(net10296));
 sg13g2_nand2b_1 _14429_ (.Y(_08011_),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23] ),
    .A_N(net10480));
 sg13g2_nand4_1 _14430_ (.B(_07770_),
    .C(_07998_),
    .A(net10480),
    .Y(_08012_),
    .D(_08005_));
 sg13g2_o21ai_1 _14431_ (.B1(_08012_),
    .Y(_08013_),
    .A1(_08002_),
    .A2(_08011_));
 sg13g2_nand3_1 _14432_ (.B(_07735_),
    .C(_08013_),
    .A(net10622),
    .Y(_08014_));
 sg13g2_xnor2_1 _14433_ (.Y(_08015_),
    .A(net10480),
    .B(_08002_));
 sg13g2_nand3b_1 _14434_ (.B(_07767_),
    .C(\u_ac_controller_soc_inst.cbus_addr[22] ),
    .Y(_08016_),
    .A_N(_08015_));
 sg13g2_a21oi_1 _14435_ (.A1(_08014_),
    .A2(_08016_),
    .Y(_08017_),
    .B1(net10301));
 sg13g2_nor2_2 _14436_ (.A(_07989_),
    .B(_07996_),
    .Y(_08018_));
 sg13g2_nand2_2 _14437_ (.Y(_08019_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15] ),
    .B(_08018_));
 sg13g2_xnor2_1 _14438_ (.Y(_08020_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[16] ),
    .B(_08019_));
 sg13g2_xnor2_1 _14439_ (.Y(_08021_),
    .A(net10481),
    .B(_07998_));
 sg13g2_nor4_1 _14440_ (.A(\u_ac_controller_soc_inst.cbus_addr[16] ),
    .B(_07760_),
    .C(_08020_),
    .D(_08021_),
    .Y(_08022_));
 sg13g2_xnor2_1 _14441_ (.Y(_08023_),
    .A(_07760_),
    .B(_08021_));
 sg13g2_and3_1 _14442_ (.X(_08024_),
    .A(\u_ac_controller_soc_inst.cbus_addr[16] ),
    .B(_08020_),
    .C(_08023_));
 sg13g2_o21ai_1 _14443_ (.B1(_07774_),
    .Y(_08025_),
    .A1(_08022_),
    .A2(_08024_));
 sg13g2_o21ai_1 _14444_ (.B1(_07774_),
    .Y(_08026_),
    .A1(\u_ac_controller_soc_inst.cbus_addr[16] ),
    .A2(\u_ac_controller_soc_inst.cbus_addr[18] ));
 sg13g2_nand3b_1 _14445_ (.B(_08021_),
    .C(_08026_),
    .Y(_08027_),
    .A_N(_08020_));
 sg13g2_nor2_1 _14446_ (.A(net10625),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15] ),
    .Y(_08028_));
 sg13g2_inv_1 _14447_ (.Y(_08029_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15] ));
 sg13g2_nand2_2 _14448_ (.Y(_08030_),
    .A(net10474),
    .B(net10473));
 sg13g2_nor4_2 _14449_ (.A(_07788_),
    .B(_07990_),
    .C(_07992_),
    .Y(_08031_),
    .D(_08030_));
 sg13g2_buf_16 clkbuf_leaf_672_clk (.X(clknet_leaf_672_clk),
    .A(clknet_8_250_0_clk));
 sg13g2_nand3_1 _14451_ (.B(net10483),
    .C(_08031_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[11] ),
    .Y(_08033_));
 sg13g2_buf_16 clkbuf_leaf_671_clk (.X(clknet_leaf_671_clk),
    .A(clknet_8_249_0_clk));
 sg13g2_xor2_1 _14453_ (.B(_08033_),
    .A(net10482),
    .X(_08035_));
 sg13g2_nand2b_1 _14454_ (.Y(_08036_),
    .B(net10482),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[14] ));
 sg13g2_mux2_1 _14455_ (.A0(_08036_),
    .A1(net10482),
    .S(_08033_),
    .X(_08037_));
 sg13g2_nand2_2 _14456_ (.Y(_08038_),
    .A(net10625),
    .B(_07774_));
 sg13g2_mux2_1 _14457_ (.A0(_08035_),
    .A1(_08037_),
    .S(_08038_),
    .X(_08039_));
 sg13g2_nor2_1 _14458_ (.A(_08029_),
    .B(_08039_),
    .Y(_08040_));
 sg13g2_a21oi_1 _14459_ (.A1(_08018_),
    .A2(_08028_),
    .Y(_08041_),
    .B1(_08040_));
 sg13g2_inv_1 _14460_ (.Y(_08042_),
    .A(_08019_));
 sg13g2_nor2_1 _14461_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15] ),
    .B(_08039_),
    .Y(_08043_));
 sg13g2_a21oi_1 _14462_ (.A1(_08042_),
    .A2(_08038_),
    .Y(_08044_),
    .B1(_08043_));
 sg13g2_nand2_1 _14463_ (.Y(_08045_),
    .A(\u_ac_controller_soc_inst.cbus_addr[15] ),
    .B(_07774_));
 sg13g2_mux2_1 _14464_ (.A0(_08041_),
    .A1(_08044_),
    .S(_08045_),
    .X(_08046_));
 sg13g2_a21oi_2 _14465_ (.B1(_08046_),
    .Y(_08047_),
    .A2(_08027_),
    .A1(_08025_));
 sg13g2_o21ai_1 _14466_ (.B1(_08047_),
    .Y(_08048_),
    .A1(_08010_),
    .A2(_08017_));
 sg13g2_xor2_1 _14467_ (.B(net10291),
    .A(net10484),
    .X(_08049_));
 sg13g2_nand2_1 _14468_ (.Y(_08050_),
    .A(_07739_),
    .B(net10483));
 sg13g2_and3_1 _14469_ (.X(_08051_),
    .A(_07746_),
    .B(_08049_),
    .C(_08050_));
 sg13g2_inv_1 _14470_ (.Y(_08052_),
    .A(net10483));
 sg13g2_and2_1 _14471_ (.A(_08052_),
    .B(net10291),
    .X(_08053_));
 sg13g2_nor3_1 _14472_ (.A(net10484),
    .B(_08052_),
    .C(net10291),
    .Y(_08054_));
 sg13g2_a21oi_1 _14473_ (.A1(net10484),
    .A2(_08053_),
    .Y(_08055_),
    .B1(_08054_));
 sg13g2_nor3_1 _14474_ (.A(_07739_),
    .B(net10626),
    .C(_08055_),
    .Y(_08056_));
 sg13g2_a21oi_1 _14475_ (.A1(net10626),
    .A2(_08051_),
    .Y(_08057_),
    .B1(_08056_));
 sg13g2_nor2_1 _14476_ (.A(\u_ac_controller_soc_inst.cbus_addr[12] ),
    .B(net10626),
    .Y(_08058_));
 sg13g2_nor3_1 _14477_ (.A(net10484),
    .B(net10483),
    .C(net10291),
    .Y(_08059_));
 sg13g2_nand3_1 _14478_ (.B(net10483),
    .C(net10291),
    .A(net10484),
    .Y(_08060_));
 sg13g2_nand2b_1 _14479_ (.Y(_08061_),
    .B(_08060_),
    .A_N(_08059_));
 sg13g2_o21ai_1 _14480_ (.B1(_08061_),
    .Y(_08062_),
    .A1(net10300),
    .A2(_08058_));
 sg13g2_o21ai_1 _14481_ (.B1(_08062_),
    .Y(_08063_),
    .A1(net10300),
    .A2(_08057_));
 sg13g2_and3_2 _14482_ (.X(_08064_),
    .A(net10479),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[3] ),
    .C(net10477));
 sg13g2_buf_16 clkbuf_leaf_669_clk (.X(clknet_leaf_669_clk),
    .A(clknet_8_255_0_clk));
 sg13g2_and3_2 _14484_ (.X(_08066_),
    .A(net10476),
    .B(net10475),
    .C(_08064_));
 sg13g2_buf_16 clkbuf_leaf_668_clk (.X(clknet_leaf_668_clk),
    .A(clknet_8_252_0_clk));
 sg13g2_nor3_1 _14486_ (.A(net10476),
    .B(net10475),
    .C(_08064_),
    .Y(_08068_));
 sg13g2_buf_16 clkbuf_leaf_667_clk (.X(clknet_leaf_667_clk),
    .A(clknet_8_252_0_clk));
 sg13g2_o21ai_1 _14488_ (.B1(net10297),
    .Y(_08070_),
    .A1(net10616),
    .A2(net10614));
 sg13g2_o21ai_1 _14489_ (.B1(_08070_),
    .Y(_08071_),
    .A1(_08066_),
    .A2(_08068_));
 sg13g2_xnor2_1 _14490_ (.Y(_08072_),
    .A(net10476),
    .B(_07990_));
 sg13g2_nor3_1 _14491_ (.A(net10616),
    .B(net10476),
    .C(_08064_),
    .Y(_08073_));
 sg13g2_a21o_1 _14492_ (.A2(_08072_),
    .A1(net10616),
    .B1(_08073_),
    .X(_08074_));
 sg13g2_nand2_1 _14493_ (.Y(_08075_),
    .A(net10476),
    .B(_08064_));
 sg13g2_nor3_1 _14494_ (.A(net10616),
    .B(net10475),
    .C(_08075_),
    .Y(_08076_));
 sg13g2_a21o_1 _14495_ (.A2(_08074_),
    .A1(net10475),
    .B1(_08076_),
    .X(_08077_));
 sg13g2_inv_2 _14496_ (.Y(_08078_),
    .A(net10615));
 sg13g2_nor3_1 _14497_ (.A(_08078_),
    .B(net10614),
    .C(net10475),
    .Y(_08079_));
 sg13g2_a22oi_1 _14498_ (.Y(_08080_),
    .B1(_08079_),
    .B2(_08072_),
    .A2(_08077_),
    .A1(net10614));
 sg13g2_nand2b_1 _14499_ (.Y(_08081_),
    .B(net10296),
    .A_N(_08080_));
 sg13g2_inv_2 _14500_ (.Y(_08082_),
    .A(net10620));
 sg13g2_buf_16 clkbuf_leaf_666_clk (.X(clknet_leaf_666_clk),
    .A(clknet_8_252_0_clk));
 sg13g2_buf_16 clkbuf_leaf_660_clk (.X(clknet_leaf_660_clk),
    .A(clknet_8_244_0_clk));
 sg13g2_xnor2_1 _14503_ (.Y(_08085_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[7] ),
    .B(_08066_));
 sg13g2_xnor2_1 _14504_ (.Y(_08086_),
    .A(net10613),
    .B(_08085_));
 sg13g2_nor3_1 _14505_ (.A(_08082_),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2] ),
    .C(_08086_),
    .Y(_08087_));
 sg13g2_nand2_1 _14506_ (.Y(_08088_),
    .A(net10613),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2] ));
 sg13g2_nor3_1 _14507_ (.A(net10621),
    .B(_08085_),
    .C(_08088_),
    .Y(_08089_));
 sg13g2_o21ai_1 _14508_ (.B1(net10296),
    .Y(_08090_),
    .A1(_08087_),
    .A2(_08089_));
 sg13g2_o21ai_1 _14509_ (.B1(net10296),
    .Y(_08091_),
    .A1(net10621),
    .A2(net10613));
 sg13g2_nand3_1 _14510_ (.B(_08085_),
    .C(_08091_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2] ),
    .Y(_08092_));
 sg13g2_a22oi_1 _14511_ (.Y(_08093_),
    .B1(_08090_),
    .B2(_08092_),
    .A2(_08081_),
    .A1(_08071_));
 sg13g2_nor2_1 _14512_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[17] ),
    .B(_08006_),
    .Y(_08094_));
 sg13g2_or2_1 _14513_ (.X(_08095_),
    .B(_08094_),
    .A(_07998_));
 sg13g2_inv_1 _14514_ (.Y(_08096_),
    .A(net10481));
 sg13g2_a21oi_1 _14515_ (.A1(_08096_),
    .A2(_07998_),
    .Y(_08097_),
    .B1(_08094_));
 sg13g2_nand2_2 _14516_ (.Y(_08098_),
    .A(\u_ac_controller_soc_inst.cbus_addr[17] ),
    .B(net10295));
 sg13g2_mux2_1 _14517_ (.A0(_08095_),
    .A1(_08097_),
    .S(_08098_),
    .X(_08099_));
 sg13g2_nand2_2 _14518_ (.Y(_08100_),
    .A(\u_ac_controller_soc_inst.cbus_addr[19] ),
    .B(_07774_));
 sg13g2_xnor2_1 _14519_ (.Y(_08101_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19] ),
    .B(_08100_));
 sg13g2_nand4_1 _14520_ (.B(_08007_),
    .C(_08098_),
    .A(net10481),
    .Y(_08102_),
    .D(_08101_));
 sg13g2_o21ai_1 _14521_ (.B1(_08102_),
    .Y(_08103_),
    .A1(_08099_),
    .A2(_08101_));
 sg13g2_xnor2_1 _14522_ (.Y(_08104_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[14] ),
    .B(_07729_));
 sg13g2_nor3_2 _14523_ (.A(_07990_),
    .B(_07992_),
    .C(_08030_),
    .Y(_08105_));
 sg13g2_nand2_1 _14524_ (.Y(_08106_),
    .A(_07988_),
    .B(_08105_));
 sg13g2_xnor2_1 _14525_ (.Y(_08107_),
    .A(_08104_),
    .B(_08106_));
 sg13g2_nand2_2 _14526_ (.Y(_08108_),
    .A(\u_ac_controller_soc_inst.cbus_addr[10] ),
    .B(net10295));
 sg13g2_xnor2_1 _14527_ (.Y(_08109_),
    .A(_07788_),
    .B(_08108_));
 sg13g2_xnor2_1 _14528_ (.Y(_08110_),
    .A(_08105_),
    .B(_08109_));
 sg13g2_nand2_1 _14529_ (.Y(_08111_),
    .A(net10623),
    .B(net10296));
 sg13g2_xnor2_1 _14530_ (.Y(_08112_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21] ),
    .B(_08111_));
 sg13g2_xnor2_1 _14531_ (.Y(_08113_),
    .A(_08000_),
    .B(_08112_));
 sg13g2_nand2_1 _14532_ (.Y(_08114_),
    .A(net10624),
    .B(net10296));
 sg13g2_xnor2_1 _14533_ (.Y(_08115_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20] ),
    .B(_08114_));
 sg13g2_and3_2 _14534_ (.X(_08116_),
    .A(net10481),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19] ),
    .C(_08007_));
 sg13g2_buf_16 clkbuf_leaf_658_clk (.X(clknet_leaf_658_clk),
    .A(clknet_8_246_0_clk));
 sg13g2_xnor2_1 _14536_ (.Y(_08118_),
    .A(_08115_),
    .B(_08116_));
 sg13g2_buf_16 clkbuf_leaf_657_clk (.X(clknet_leaf_657_clk),
    .A(clknet_8_245_0_clk));
 sg13g2_xor2_1 _14538_ (.B(net10478),
    .A(net10479),
    .X(_08120_));
 sg13g2_nor3_1 _14539_ (.A(net10619),
    .B(net10479),
    .C(net10478),
    .Y(_08121_));
 sg13g2_a21o_1 _14540_ (.A2(_08120_),
    .A1(net10619),
    .B1(_08121_),
    .X(_08122_));
 sg13g2_nand2_1 _14541_ (.Y(_08123_),
    .A(net10479),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[3] ));
 sg13g2_nor3_1 _14542_ (.A(net10619),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[4] ),
    .C(_08123_),
    .Y(_08124_));
 sg13g2_a21o_1 _14543_ (.A2(_08122_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[4] ),
    .B1(_08124_),
    .X(_08125_));
 sg13g2_inv_8 _14544_ (.Y(_08126_),
    .A(\u_ac_controller_soc_inst.cbus_addr[3] ));
 sg13g2_nor3_1 _14545_ (.A(_08126_),
    .B(\u_ac_controller_soc_inst.cbus_addr[4] ),
    .C(net10477),
    .Y(_08127_));
 sg13g2_a22oi_1 _14546_ (.Y(_08128_),
    .B1(_08127_),
    .B2(_08120_),
    .A2(_08125_),
    .A1(\u_ac_controller_soc_inst.cbus_addr[4] ));
 sg13g2_nor3_1 _14547_ (.A(net10479),
    .B(net10478),
    .C(net10477),
    .Y(_08129_));
 sg13g2_o21ai_1 _14548_ (.B1(net10296),
    .Y(_08130_),
    .A1(net10619),
    .A2(\u_ac_controller_soc_inst.cbus_addr[4] ));
 sg13g2_o21ai_1 _14549_ (.B1(_08130_),
    .Y(_08131_),
    .A1(_08064_),
    .A2(_08129_));
 sg13g2_o21ai_1 _14550_ (.B1(_08131_),
    .Y(_08132_),
    .A1(net10301),
    .A2(_08128_));
 sg13g2_nand4_1 _14551_ (.B(_08113_),
    .C(_08118_),
    .A(_08009_),
    .Y(_08133_),
    .D(_08132_));
 sg13g2_buf_16 clkbuf_leaf_656_clk (.X(clknet_leaf_656_clk),
    .A(clknet_8_245_0_clk));
 sg13g2_o21ai_1 _14553_ (.B1(net10295),
    .Y(_08135_),
    .A1(net10612),
    .A2(net10611));
 sg13g2_or2_1 _14554_ (.X(_08136_),
    .B(net10473),
    .A(net10474));
 sg13g2_o21ai_1 _14555_ (.B1(_07996_),
    .Y(_08137_),
    .A1(_07994_),
    .A2(_08136_));
 sg13g2_xor2_1 _14556_ (.B(_07994_),
    .A(net10474),
    .X(_08138_));
 sg13g2_nor3_1 _14557_ (.A(net10612),
    .B(net10474),
    .C(_07994_),
    .Y(_08139_));
 sg13g2_a21oi_1 _14558_ (.A1(net10612),
    .A2(_08138_),
    .Y(_08140_),
    .B1(_08139_));
 sg13g2_nor2b_1 _14559_ (.A(_08140_),
    .B_N(net10473),
    .Y(_08141_));
 sg13g2_nand2_1 _14560_ (.Y(_08142_),
    .A(net10474),
    .B(_07994_));
 sg13g2_nor3_1 _14561_ (.A(net10612),
    .B(net10473),
    .C(_08142_),
    .Y(_08143_));
 sg13g2_o21ai_1 _14562_ (.B1(\u_ac_controller_soc_inst.cbus_addr[9] ),
    .Y(_08144_),
    .A1(_08141_),
    .A2(_08143_));
 sg13g2_nand3_1 _14563_ (.B(_07862_),
    .C(_08138_),
    .A(net10612),
    .Y(_08145_));
 sg13g2_nand2_1 _14564_ (.Y(_08146_),
    .A(_08144_),
    .B(_08145_));
 sg13g2_a22oi_1 _14565_ (.Y(_08147_),
    .B1(_08146_),
    .B2(net10295),
    .A2(_08137_),
    .A1(_08135_));
 sg13g2_nor4_1 _14566_ (.A(_08107_),
    .B(_08110_),
    .C(_08133_),
    .D(_08147_),
    .Y(_08148_));
 sg13g2_nand4_1 _14567_ (.B(_08093_),
    .C(_08103_),
    .A(_08063_),
    .Y(_08149_),
    .D(_08148_));
 sg13g2_o21ai_1 _14568_ (.B1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_valid ),
    .Y(_08150_),
    .A1(_08048_),
    .A2(_08149_));
 sg13g2_nor2_2 _14569_ (.A(_07982_),
    .B(_08150_),
    .Y(_08151_));
 sg13g2_buf_16 clkbuf_leaf_654_clk (.X(clknet_leaf_654_clk),
    .A(clknet_8_247_0_clk));
 sg13g2_buf_16 clkbuf_leaf_653_clk (.X(clknet_leaf_653_clk),
    .A(clknet_8_246_0_clk));
 sg13g2_buf_16 clkbuf_leaf_652_clk (.X(clknet_leaf_652_clk),
    .A(clknet_8_247_0_clk));
 sg13g2_buf_16 clkbuf_leaf_650_clk (.X(clknet_leaf_650_clk),
    .A(clknet_8_246_0_clk));
 sg13g2_buf_16 clkbuf_leaf_648_clk (.X(clknet_leaf_648_clk),
    .A(clknet_8_194_0_clk));
 sg13g2_buf_16 clkbuf_leaf_647_clk (.X(clknet_leaf_647_clk),
    .A(clknet_8_194_0_clk));
 sg13g2_nor3_1 _14576_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[0] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1] ),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[3] ),
    .Y(_08158_));
 sg13g2_nor2b_1 _14577_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2] ),
    .B_N(_08158_),
    .Y(_08159_));
 sg13g2_buf_16 clkbuf_leaf_646_clk (.X(clknet_leaf_646_clk),
    .A(clknet_8_252_0_clk));
 sg13g2_buf_16 clkbuf_leaf_645_clk (.X(clknet_leaf_645_clk),
    .A(clknet_8_247_0_clk));
 sg13g2_nor2_1 _14580_ (.A(net10467),
    .B(net10466),
    .Y(_08162_));
 sg13g2_nor2_1 _14581_ (.A(_08159_),
    .B(_08162_),
    .Y(_08163_));
 sg13g2_xor2_1 _14582_ (.B(_08163_),
    .A(_00093_),
    .X(_08164_));
 sg13g2_buf_16 clkbuf_leaf_644_clk (.X(clknet_leaf_644_clk),
    .A(clknet_8_246_0_clk));
 sg13g2_buf_16 clkbuf_leaf_641_clk (.X(clknet_leaf_641_clk),
    .A(clknet_8_253_0_clk));
 sg13g2_nand2_1 _14585_ (.Y(_08167_),
    .A(_00092_),
    .B(net10465));
 sg13g2_nor3_1 _14586_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[0] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1] ),
    .C(_08167_),
    .Y(_08168_));
 sg13g2_buf_16 clkbuf_leaf_640_clk (.X(clknet_leaf_640_clk),
    .A(clknet_8_255_0_clk));
 sg13g2_buf_16 clkbuf_leaf_636_clk (.X(clknet_leaf_636_clk),
    .A(clknet_8_253_0_clk));
 sg13g2_or4_1 _14589_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[0] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1] ),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2] ),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[3] ),
    .X(_08171_));
 sg13g2_buf_16 clkbuf_leaf_634_clk (.X(clknet_leaf_634_clk),
    .A(clknet_8_195_0_clk));
 sg13g2_xor2_1 _14591_ (.B(_08171_),
    .A(_00091_),
    .X(_08173_));
 sg13g2_nor2_1 _14592_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1] ),
    .B(net10467),
    .Y(_08174_));
 sg13g2_a21oi_1 _14593_ (.A1(net10467),
    .A2(_08173_),
    .Y(_08175_),
    .B1(_08174_));
 sg13g2_nand2_1 _14594_ (.Y(_08176_),
    .A(_00091_),
    .B(net10467));
 sg13g2_nor3_1 _14595_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2] ),
    .B(_08158_),
    .C(_08176_),
    .Y(_08177_));
 sg13g2_a21o_1 _14596_ (.A2(_08176_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2] ),
    .B1(_08177_),
    .X(_08178_));
 sg13g2_buf_16 clkbuf_leaf_633_clk (.X(clknet_leaf_633_clk),
    .A(clknet_8_200_0_clk));
 sg13g2_nand2b_2 _14598_ (.Y(_08180_),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi ),
    .A_N(net10465));
 sg13g2_buf_16 clkbuf_leaf_631_clk (.X(clknet_leaf_631_clk),
    .A(clknet_8_200_0_clk));
 sg13g2_nand2b_1 _14600_ (.Y(_08182_),
    .B(_00092_),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[0] ));
 sg13g2_nor4_1 _14601_ (.A(_08175_),
    .B(_08178_),
    .C(_08180_),
    .D(_08182_),
    .Y(_08183_));
 sg13g2_a21oi_1 _14602_ (.A1(_08164_),
    .A2(_08168_),
    .Y(_08184_),
    .B1(_08183_));
 sg13g2_nor2b_1 _14603_ (.A(_00093_),
    .B_N(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2] ),
    .Y(_08185_));
 sg13g2_nand3_1 _14604_ (.B(_00094_),
    .C(_08171_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk ),
    .Y(_08186_));
 sg13g2_buf_16 clkbuf_leaf_627_clk (.X(clknet_leaf_627_clk),
    .A(clknet_8_204_0_clk));
 sg13g2_nor2_2 _14606_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1] ),
    .B(_08186_),
    .Y(_08188_));
 sg13g2_mux2_1 _14607_ (.A0(_00093_),
    .A1(_08185_),
    .S(_08188_),
    .X(_08189_));
 sg13g2_nor3_2 _14608_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2] ),
    .C(_08186_),
    .Y(_08190_));
 sg13g2_nor2_1 _14609_ (.A(_00092_),
    .B(_00093_),
    .Y(_08191_));
 sg13g2_a22oi_1 _14610_ (.Y(_08192_),
    .B1(_08190_),
    .B2(_08191_),
    .A2(_08189_),
    .A1(_00092_));
 sg13g2_inv_1 _14611_ (.Y(_08193_),
    .A(_00094_));
 sg13g2_xnor2_1 _14612_ (.Y(_08194_),
    .A(_08193_),
    .B(_08171_));
 sg13g2_nor2_1 _14613_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[0] ),
    .B(net10467),
    .Y(_08195_));
 sg13g2_a21oi_1 _14614_ (.A1(net10467),
    .A2(_08194_),
    .Y(_08196_),
    .B1(_08195_));
 sg13g2_nor3_2 _14615_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi ),
    .B(net10462),
    .C(net10466),
    .Y(_08197_));
 sg13g2_buf_16 clkbuf_leaf_625_clk (.X(clknet_leaf_625_clk),
    .A(clknet_8_204_0_clk));
 sg13g2_nand2_1 _14617_ (.Y(_08199_),
    .A(_00091_),
    .B(_08197_));
 sg13g2_or3_1 _14618_ (.A(_08192_),
    .B(_08196_),
    .C(_08199_),
    .X(_08200_));
 sg13g2_buf_16 clkbuf_leaf_624_clk (.X(clknet_leaf_624_clk),
    .A(clknet_8_206_0_clk));
 sg13g2_buf_16 clkbuf_leaf_622_clk (.X(clknet_leaf_622_clk),
    .A(clknet_8_207_0_clk));
 sg13g2_buf_16 clkbuf_leaf_621_clk (.X(clknet_leaf_621_clk),
    .A(clknet_8_203_0_clk));
 sg13g2_or4_1 _14622_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[0] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[1] ),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[3] ),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[2] ),
    .X(_08204_));
 sg13g2_buf_16 clkbuf_leaf_620_clk (.X(clknet_leaf_620_clk),
    .A(clknet_8_202_0_clk));
 sg13g2_a21oi_2 _14624_ (.B1(_08204_),
    .Y(_08206_),
    .A2(_08200_),
    .A1(_08184_));
 sg13g2_and2_1 _14625_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_valid ),
    .B(_08206_),
    .X(_08207_));
 sg13g2_buf_16 clkbuf_leaf_618_clk (.X(clknet_leaf_618_clk),
    .A(clknet_8_201_0_clk));
 sg13g2_nand2_1 _14627_ (.Y(_08209_),
    .A(net10461),
    .B(net9747));
 sg13g2_buf_16 clkbuf_leaf_615_clk (.X(clknet_leaf_615_clk),
    .A(clknet_8_202_0_clk));
 sg13g2_buf_16 clkbuf_leaf_613_clk (.X(clknet_leaf_613_clk),
    .A(clknet_8_237_0_clk));
 sg13g2_nand2_1 _14630_ (.Y(_08212_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[0] ),
    .B(net9727));
 sg13g2_inv_4 _14631_ (.A(net11056),
    .Y(_08213_));
 sg13g2_buf_16 clkbuf_leaf_611_clk (.X(clknet_leaf_611_clk),
    .A(clknet_8_228_0_clk));
 sg13g2_nor2_2 _14633_ (.A(net10979),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.softreset ),
    .Y(_08215_));
 sg13g2_o21ai_1 _14634_ (.B1(_08215_),
    .Y(_00020_),
    .A1(_08151_),
    .A2(_08212_));
 sg13g2_buf_16 clkbuf_leaf_609_clk (.X(clknet_leaf_609_clk),
    .A(clknet_8_229_0_clk));
 sg13g2_nand2_1 _14636_ (.Y(_08217_),
    .A(net10470),
    .B(net9728));
 sg13g2_buf_16 clkbuf_leaf_608_clk (.X(clknet_leaf_608_clk),
    .A(clknet_8_255_0_clk));
 sg13g2_buf_16 clkbuf_leaf_607_clk (.X(clknet_leaf_607_clk),
    .A(clknet_8_253_0_clk));
 sg13g2_inv_4 _14639_ (.A(net10461),
    .Y(_08220_));
 sg13g2_inv_4 _14640_ (.A(net9747),
    .Y(_08221_));
 sg13g2_nor2_1 _14641_ (.A(_08220_),
    .B(_08221_),
    .Y(_08222_));
 sg13g2_buf_16 clkbuf_leaf_606_clk (.X(clknet_leaf_606_clk),
    .A(clknet_8_228_0_clk));
 sg13g2_buf_16 clkbuf_leaf_605_clk (.X(clknet_leaf_605_clk),
    .A(clknet_8_228_0_clk));
 sg13g2_buf_16 clkbuf_leaf_604_clk (.X(clknet_leaf_604_clk),
    .A(clknet_8_229_0_clk));
 sg13g2_or2_1 _14645_ (.X(_08226_),
    .B(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[21] ),
    .A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[22] ));
 sg13g2_nand3_1 _14646_ (.B(net9707),
    .C(_08226_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[12] ),
    .Y(_08227_));
 sg13g2_o21ai_1 _14647_ (.B1(_08215_),
    .Y(_08228_),
    .A1(_07982_),
    .A2(_08150_));
 sg13g2_buf_16 clkbuf_leaf_603_clk (.X(clknet_leaf_603_clk),
    .A(clknet_8_231_0_clk));
 sg13g2_buf_16 clkbuf_leaf_602_clk (.X(clknet_leaf_602_clk),
    .A(clknet_8_237_0_clk));
 sg13g2_a21oi_1 _14650_ (.A1(_08217_),
    .A2(_08227_),
    .Y(_00024_),
    .B1(_08228_));
 sg13g2_nand2b_2 _14651_ (.Y(_08231_),
    .B(net11040),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.softreset ));
 sg13g2_buf_16 clkbuf_leaf_601_clk (.X(clknet_leaf_601_clk),
    .A(clknet_8_231_0_clk));
 sg13g2_and2_1 _14653_ (.A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[20] ),
    .B(_08151_),
    .X(_08233_));
 sg13g2_buf_16 clkbuf_leaf_599_clk (.X(clknet_leaf_599_clk),
    .A(clknet_8_237_0_clk));
 sg13g2_buf_16 clkbuf_leaf_596_clk (.X(clknet_leaf_596_clk),
    .A(clknet_8_236_0_clk));
 sg13g2_buf_16 clkbuf_leaf_594_clk (.X(clknet_leaf_594_clk),
    .A(clknet_8_202_0_clk));
 sg13g2_nor2b_1 _14657_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.last_fetch ),
    .B_N(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr_q ),
    .Y(_08237_));
 sg13g2_nor2_1 _14658_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.fetch ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr_q ),
    .Y(_08238_));
 sg13g2_a22oi_1 _14659_ (.Y(_08239_),
    .B1(_08238_),
    .B2(_08206_),
    .A2(_08237_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.fetch ));
 sg13g2_nor2_2 _14660_ (.A(_00095_),
    .B(_08239_),
    .Y(_08240_));
 sg13g2_a221oi_1 _14661_ (.B2(\u_ac_controller_soc_inst.u_spi_flash_mem.state[10] ),
    .C1(_08151_),
    .B1(_08240_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[2] ),
    .Y(_08241_),
    .A2(net9727));
 sg13g2_nor3_1 _14662_ (.A(net10455),
    .B(_08233_),
    .C(_08241_),
    .Y(_00025_));
 sg13g2_buf_16 clkbuf_leaf_593_clk (.X(clknet_leaf_593_clk),
    .A(clknet_8_203_0_clk));
 sg13g2_nand2_2 _14664_ (.Y(_08243_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_wait ),
    .B(_07744_));
 sg13g2_nand2_1 _14665_ (.Y(_08244_),
    .A(net9707),
    .B(_08243_));
 sg13g2_buf_16 clkbuf_leaf_592_clk (.X(clknet_leaf_592_clk),
    .A(clknet_8_203_0_clk));
 sg13g2_a22oi_1 _14667_ (.Y(_08246_),
    .B1(_08244_),
    .B2(\u_ac_controller_soc_inst.u_spi_flash_mem.state[3] ),
    .A2(net9707),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[11] ));
 sg13g2_nor2_1 _14668_ (.A(_08228_),
    .B(_08246_),
    .Y(_00026_));
 sg13g2_buf_16 clkbuf_leaf_591_clk (.X(clknet_leaf_591_clk),
    .A(clknet_8_207_0_clk));
 sg13g2_a22oi_1 _14670_ (.Y(_08248_),
    .B1(_08240_),
    .B2(\u_ac_controller_soc_inst.u_spi_flash_mem.state[7] ),
    .A2(net9726),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[4] ));
 sg13g2_nor2_1 _14671_ (.A(net9653),
    .B(_08248_),
    .Y(_00027_));
 sg13g2_buf_16 clkbuf_leaf_590_clk (.X(clknet_leaf_590_clk),
    .A(clknet_8_206_0_clk));
 sg13g2_nand2_1 _14673_ (.Y(_08250_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[8] ),
    .B(net9705));
 sg13g2_buf_16 clkbuf_leaf_587_clk (.X(clknet_leaf_587_clk),
    .A(clknet_8_218_0_clk));
 sg13g2_nand2_1 _14675_ (.Y(_08252_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[5] ),
    .B(net9726));
 sg13g2_a21oi_1 _14676_ (.A1(_08250_),
    .A2(_08252_),
    .Y(_00028_),
    .B1(net9653));
 sg13g2_buf_16 clkbuf_leaf_586_clk (.X(clknet_leaf_586_clk),
    .A(clknet_8_207_0_clk));
 sg13g2_inv_1 _14678_ (.Y(_08254_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[9] ));
 sg13g2_or2_1 _14679_ (.X(_08255_),
    .B(_07982_),
    .A(_08254_));
 sg13g2_buf_16 clkbuf_leaf_585_clk (.X(clknet_leaf_585_clk),
    .A(clknet_8_218_0_clk));
 sg13g2_nor2_1 _14681_ (.A(net9727),
    .B(_08255_),
    .Y(_08257_));
 sg13g2_a21oi_1 _14682_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[6] ),
    .A2(net9727),
    .Y(_08258_),
    .B1(_08257_));
 sg13g2_nor2_1 _14683_ (.A(_08228_),
    .B(_08258_),
    .Y(_00029_));
 sg13g2_or2_1 _14684_ (.X(_08259_),
    .B(_08239_),
    .A(_00095_));
 sg13g2_buf_16 clkbuf_leaf_584_clk (.X(clknet_leaf_584_clk),
    .A(clknet_8_223_0_clk));
 sg13g2_a22oi_1 _14686_ (.Y(_08261_),
    .B1(_08259_),
    .B2(\u_ac_controller_soc_inst.u_spi_flash_mem.state[7] ),
    .A2(net9706),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[0] ));
 sg13g2_nor2_1 _14687_ (.A(net9653),
    .B(_08261_),
    .Y(_00030_));
 sg13g2_a21oi_1 _14688_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[3] ),
    .A2(_08243_),
    .Y(_08262_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[1] ));
 sg13g2_buf_16 clkbuf_leaf_583_clk (.X(clknet_leaf_583_clk),
    .A(clknet_8_223_0_clk));
 sg13g2_inv_4 _14690_ (.A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[21] ),
    .Y(_08264_));
 sg13g2_nand3b_1 _14691_ (.B(_08264_),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.state[12] ),
    .Y(_08265_),
    .A_N(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[22] ));
 sg13g2_a21oi_1 _14692_ (.A1(_08262_),
    .A2(_08265_),
    .Y(_08266_),
    .B1(net9727));
 sg13g2_a21oi_1 _14693_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[8] ),
    .A2(net9726),
    .Y(_08267_),
    .B1(_08266_));
 sg13g2_nor2_1 _14694_ (.A(net9653),
    .B(_08267_),
    .Y(_00031_));
 sg13g2_nand2_1 _14695_ (.Y(_08268_),
    .A(net10469),
    .B(net9707));
 sg13g2_mux2_1 _14696_ (.A0(_08268_),
    .A1(_00098_),
    .S(_08151_),
    .X(_08269_));
 sg13g2_a21oi_1 _14697_ (.A1(_08150_),
    .A2(net9727),
    .Y(_08270_),
    .B1(_07982_));
 sg13g2_nand2b_1 _14698_ (.Y(_08271_),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.state[9] ),
    .A_N(_08270_));
 sg13g2_a21oi_1 _14699_ (.A1(_08269_),
    .A2(_08271_),
    .Y(_00032_),
    .B1(net10455));
 sg13g2_a22oi_1 _14700_ (.Y(_08272_),
    .B1(_08259_),
    .B2(\u_ac_controller_soc_inst.u_spi_flash_mem.state[10] ),
    .A2(net9706),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[4] ));
 sg13g2_nor2_1 _14701_ (.A(net9653),
    .B(_08272_),
    .Y(_00021_));
 sg13g2_nand2_1 _14702_ (.Y(_08273_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[5] ),
    .B(net9706));
 sg13g2_nand2_1 _14703_ (.Y(_08274_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[11] ),
    .B(net9726));
 sg13g2_a21oi_1 _14704_ (.A1(_08273_),
    .A2(_08274_),
    .Y(_00022_),
    .B1(net9653));
 sg13g2_nand2_1 _14705_ (.Y(_08275_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[6] ),
    .B(net9707));
 sg13g2_nand2_1 _14706_ (.Y(_08276_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[12] ),
    .B(net9727));
 sg13g2_a21oi_1 _14707_ (.A1(_08275_),
    .A2(_08276_),
    .Y(_00023_),
    .B1(_08228_));
 sg13g2_buf_16 clkbuf_leaf_582_clk (.X(clknet_leaf_582_clk),
    .A(clknet_8_219_0_clk));
 sg13g2_buf_16 clkbuf_leaf_581_clk (.X(clknet_leaf_581_clk),
    .A(clknet_8_222_0_clk));
 sg13g2_buf_16 clkbuf_leaf_580_clk (.X(clknet_leaf_580_clk),
    .A(clknet_8_222_0_clk));
 sg13g2_buf_16 clkbuf_leaf_579_clk (.X(clknet_leaf_579_clk),
    .A(clknet_8_219_0_clk));
 sg13g2_o21ai_1 _14712_ (.B1(net10597),
    .Y(_08281_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[0] ));
 sg13g2_buf_16 clkbuf_leaf_578_clk (.X(clknet_leaf_578_clk),
    .A(clknet_8_217_0_clk));
 sg13g2_buf_16 clkbuf_leaf_574_clk (.X(clknet_leaf_574_clk),
    .A(clknet_8_218_0_clk));
 sg13g2_nand2_1 _14715_ (.Y(_08284_),
    .A(net10568),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[0] ));
 sg13g2_nor2_1 _14716_ (.A(net10610),
    .B(net10609),
    .Y(_08285_));
 sg13g2_a21oi_1 _14717_ (.A1(_08281_),
    .A2(_08284_),
    .Y(_08286_),
    .B1(_08285_));
 sg13g2_a21oi_2 _14718_ (.B1(_08286_),
    .Y(_08287_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_pc[1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_do_rinst ));
 sg13g2_buf_16 clkbuf_leaf_572_clk (.X(clknet_leaf_572_clk),
    .A(clknet_8_205_0_clk));
 sg13g2_nand2_1 _14720_ (.Y(_08289_),
    .A(net11050),
    .B(_08287_));
 sg13g2_buf_16 clkbuf_leaf_571_clk (.X(clknet_leaf_571_clk),
    .A(clknet_8_220_0_clk));
 sg13g2_buf_16 clkbuf_leaf_570_clk (.X(clknet_leaf_570_clk),
    .A(clknet_8_217_0_clk));
 sg13g2_nor2_2 _14723_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_or ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_ori ),
    .Y(_08292_));
 sg13g2_buf_16 clkbuf_leaf_569_clk (.X(clknet_leaf_569_clk),
    .A(clknet_8_222_0_clk));
 sg13g2_nor2_2 _14725_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_xor ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_xori ),
    .Y(_08294_));
 sg13g2_and2_1 _14726_ (.A(_08292_),
    .B(_08294_),
    .X(_08295_));
 sg13g2_nor4_2 _14727_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_addi ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_bltu ),
    .C(\u_ac_controller_soc_inst.u_picorv32.instr_blt ),
    .Y(_08296_),
    .D(\u_ac_controller_soc_inst.u_picorv32.instr_beq ));
 sg13g2_nor2_2 _14728_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_and ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_andi ),
    .Y(_08297_));
 sg13g2_buf_16 clkbuf_leaf_567_clk (.X(clknet_leaf_567_clk),
    .A(clknet_8_222_0_clk));
 sg13g2_buf_16 clkbuf_leaf_566_clk (.X(clknet_leaf_566_clk),
    .A(clknet_8_216_0_clk));
 sg13g2_buf_16 clkbuf_leaf_565_clk (.X(clknet_leaf_565_clk),
    .A(clknet_8_220_0_clk));
 sg13g2_nor4_1 _14732_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_fence ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_sub ),
    .C(\u_ac_controller_soc_inst.u_picorv32.instr_add ),
    .D(\u_ac_controller_soc_inst.u_picorv32.instr_jalr ),
    .Y(_08301_));
 sg13g2_nand4_1 _14733_ (.B(_08296_),
    .C(_08297_),
    .A(_08295_),
    .Y(_08302_),
    .D(_08301_));
 sg13g2_nor3_2 _14734_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_bgeu ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_bge ),
    .C(\u_ac_controller_soc_inst.u_picorv32.instr_bne ),
    .Y(_08303_));
 sg13g2_nor4_2 _14735_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_sltu ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_slt ),
    .C(\u_ac_controller_soc_inst.u_picorv32.instr_sltiu ),
    .Y(_08304_),
    .D(\u_ac_controller_soc_inst.u_picorv32.instr_slti ));
 sg13g2_buf_16 clkbuf_leaf_564_clk (.X(clknet_leaf_564_clk),
    .A(clknet_8_220_0_clk));
 sg13g2_or2_1 _14737_ (.X(_08306_),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_auipc ),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_lui ));
 sg13g2_buf_16 clkbuf_leaf_559_clk (.X(clknet_leaf_559_clk),
    .A(clknet_8_221_0_clk));
 sg13g2_nor2_1 _14739_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_jal ),
    .B(_08306_),
    .Y(_08308_));
 sg13g2_nand4_1 _14740_ (.B(_08303_),
    .C(_08304_),
    .A(_07958_),
    .Y(_08309_),
    .D(_08308_));
 sg13g2_or2_1 _14741_ (.X(_08310_),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_srli ),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_srl ));
 sg13g2_buf_16 clkbuf_leaf_558_clk (.X(clknet_leaf_558_clk),
    .A(clknet_8_223_0_clk));
 sg13g2_nor2_2 _14743_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_sra ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_srai ),
    .Y(_08312_));
 sg13g2_buf_16 clkbuf_leaf_557_clk (.X(clknet_leaf_557_clk),
    .A(clknet_8_223_0_clk));
 sg13g2_nand2b_2 _14745_ (.Y(_08314_),
    .B(_08312_),
    .A_N(_08310_));
 sg13g2_buf_16 clkbuf_leaf_556_clk (.X(clknet_leaf_556_clk),
    .A(clknet_8_221_0_clk));
 sg13g2_nor3_2 _14747_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_sll ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_slli ),
    .C(_08314_),
    .Y(_08316_));
 sg13g2_buf_16 clkbuf_leaf_555_clk (.X(clknet_leaf_555_clk),
    .A(clknet_8_215_0_clk));
 sg13g2_buf_16 clkbuf_leaf_554_clk (.X(clknet_leaf_554_clk),
    .A(clknet_8_215_0_clk));
 sg13g2_buf_16 clkbuf_leaf_553_clk (.X(clknet_leaf_553_clk),
    .A(clknet_8_215_0_clk));
 sg13g2_or3_1 _14751_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstr ),
    .C(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycleh ),
    .X(_08320_));
 sg13g2_buf_16 clkbuf_leaf_552_clk (.X(clknet_leaf_552_clk),
    .A(clknet_8_213_0_clk));
 sg13g2_nor2_2 _14753_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycle ),
    .B(net10435),
    .Y(_08322_));
 sg13g2_nand3_1 _14754_ (.B(_08316_),
    .C(_08322_),
    .A(_07962_),
    .Y(_08323_));
 sg13g2_nor3_2 _14755_ (.A(_08302_),
    .B(_08309_),
    .C(_08323_),
    .Y(_08324_));
 sg13g2_nor2_2 _14756_ (.A(_00101_),
    .B(_08324_),
    .Y(_08325_));
 sg13g2_or2_1 _14757_ (.X(_08326_),
    .B(_07938_),
    .A(_07915_));
 sg13g2_buf_16 clkbuf_leaf_550_clk (.X(clknet_leaf_550_clk),
    .A(clknet_8_213_0_clk));
 sg13g2_nand2_1 _14759_ (.Y(_08328_),
    .A(_00085_),
    .B(_08326_));
 sg13g2_buf_16 clkbuf_leaf_547_clk (.X(clknet_leaf_547_clk),
    .A(clknet_8_127_0_clk));
 sg13g2_a22oi_1 _14761_ (.Y(_08330_),
    .B1(_08328_),
    .B2(net10695),
    .A2(_08325_),
    .A1(net10714));
 sg13g2_nor2_1 _14762_ (.A(_08289_),
    .B(_08330_),
    .Y(_00016_));
 sg13g2_a22oi_1 _14763_ (.Y(_08331_),
    .B1(_07954_),
    .B2(\u_ac_controller_soc_inst.u_picorv32.instr_sw ),
    .A2(_07951_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_lw ));
 sg13g2_nand2_2 _14764_ (.Y(_08332_),
    .A(net11052),
    .B(net10722));
 sg13g2_buf_16 clkbuf_leaf_546_clk (.X(clknet_leaf_546_clk),
    .A(clknet_8_213_0_clk));
 sg13g2_o21ai_1 _14766_ (.B1(_08332_),
    .Y(_08334_),
    .A1(_07946_),
    .A2(_08331_));
 sg13g2_nand2b_1 _14767_ (.Y(_08335_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[0] ),
    .A_N(_07974_));
 sg13g2_nand2b_1 _14768_ (.Y(_00017_),
    .B(_08335_),
    .A_N(_08334_));
 sg13g2_a22oi_1 _14769_ (.Y(_08336_),
    .B1(_07961_),
    .B2(_07951_),
    .A2(_07954_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_sb ));
 sg13g2_buf_16 clkbuf_leaf_543_clk (.X(clknet_leaf_543_clk),
    .A(clknet_8_123_0_clk));
 sg13g2_buf_16 clkbuf_leaf_541_clk (.X(clknet_leaf_541_clk),
    .A(clknet_8_212_0_clk));
 sg13g2_nand2b_1 _14772_ (.Y(_08339_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[1] ),
    .A_N(_07974_));
 sg13g2_o21ai_1 _14773_ (.B1(_08339_),
    .Y(_00018_),
    .A1(_07946_),
    .A2(_08336_));
 sg13g2_buf_16 clkbuf_leaf_540_clk (.X(clknet_leaf_540_clk),
    .A(clknet_8_212_0_clk));
 sg13g2_inv_2 _14775_ (.Y(_08341_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_sb_sh_sw ));
 sg13g2_buf_16 clkbuf_leaf_539_clk (.X(clknet_leaf_539_clk),
    .A(clknet_8_212_0_clk));
 sg13g2_nor4_2 _14777_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycle ),
    .B(\u_ac_controller_soc_inst.u_picorv32.is_slli_srli_srai ),
    .C(net10435),
    .Y(_08343_),
    .D(_08324_));
 sg13g2_inv_2 _14778_ (.Y(_08344_),
    .A(_00101_));
 sg13g2_nand2_1 _14779_ (.Y(_08345_),
    .A(net11051),
    .B(\u_ac_controller_soc_inst.u_picorv32.cpu_state[2] ));
 sg13g2_buf_16 clkbuf_leaf_538_clk (.X(clknet_leaf_538_clk),
    .A(clknet_8_214_0_clk));
 sg13g2_buf_16 clkbuf_leaf_537_clk (.X(clknet_leaf_537_clk),
    .A(clknet_8_215_0_clk));
 sg13g2_or2_1 _14782_ (.X(_08348_),
    .B(\u_ac_controller_soc_inst.u_picorv32.is_jalr_addi_slti_sltiu_xori_ori_andi ),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_lui_auipc_jal ));
 sg13g2_buf_16 clkbuf_leaf_535_clk (.X(clknet_leaf_535_clk),
    .A(clknet_8_214_0_clk));
 sg13g2_nor3_1 _14784_ (.A(_08344_),
    .B(_08345_),
    .C(_08348_),
    .Y(_08350_));
 sg13g2_nand3_1 _14785_ (.B(_08343_),
    .C(_08350_),
    .A(_08287_),
    .Y(_08351_));
 sg13g2_buf_16 clkbuf_leaf_534_clk (.X(clknet_leaf_534_clk),
    .A(clknet_8_214_0_clk));
 sg13g2_nand4_1 _14787_ (.B(\u_ac_controller_soc_inst.u_picorv32.cpu_state[5] ),
    .C(_08287_),
    .A(net11050),
    .Y(_08353_),
    .D(_08328_));
 sg13g2_o21ai_1 _14788_ (.B1(_08353_),
    .Y(_00015_),
    .A1(_08341_),
    .A2(_08351_));
 sg13g2_buf_16 clkbuf_leaf_533_clk (.X(clknet_leaf_533_clk),
    .A(clknet_8_212_0_clk));
 sg13g2_buf_16 clkbuf_leaf_532_clk (.X(clknet_leaf_532_clk),
    .A(clknet_8_212_0_clk));
 sg13g2_buf_16 clkbuf_leaf_530_clk (.X(clknet_leaf_530_clk),
    .A(clknet_8_122_0_clk));
 sg13g2_buf_16 clkbuf_leaf_529_clk (.X(clknet_leaf_529_clk),
    .A(clknet_8_122_0_clk));
 sg13g2_buf_16 clkbuf_leaf_528_clk (.X(clknet_leaf_528_clk),
    .A(clknet_8_122_0_clk));
 sg13g2_buf_16 clkbuf_leaf_526_clk (.X(clknet_leaf_526_clk),
    .A(clknet_8_209_0_clk));
 sg13g2_buf_16 clkbuf_leaf_525_clk (.X(clknet_leaf_525_clk),
    .A(clknet_8_110_0_clk));
 sg13g2_buf_16 clkbuf_leaf_523_clk (.X(clknet_leaf_523_clk),
    .A(clknet_8_111_0_clk));
 sg13g2_buf_16 clkbuf_leaf_519_clk (.X(clknet_leaf_519_clk),
    .A(clknet_8_209_0_clk));
 sg13g2_or3_1 _14798_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_sh[2] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_sh[3] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.reg_sh[4] ),
    .X(_08363_));
 sg13g2_buf_16 clkbuf_leaf_518_clk (.X(clknet_leaf_518_clk),
    .A(clknet_8_208_0_clk));
 sg13g2_nor3_2 _14800_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_sh[1] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_sh[0] ),
    .C(_08363_),
    .Y(_08365_));
 sg13g2_buf_16 clkbuf_leaf_517_clk (.X(clknet_leaf_517_clk),
    .A(clknet_8_210_0_clk));
 sg13g2_inv_1 _14802_ (.Y(_08367_),
    .A(_08365_));
 sg13g2_a22oi_1 _14803_ (.Y(_08368_),
    .B1(net10708),
    .B2(_08367_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.is_slli_srli_srai ),
    .A1(net10714));
 sg13g2_buf_16 clkbuf_leaf_513_clk (.X(clknet_leaf_513_clk),
    .A(clknet_8_210_0_clk));
 sg13g2_nand4_1 _14805_ (.B(_08287_),
    .C(_08343_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_sll_srl_sra ),
    .Y(_08370_),
    .D(_08350_));
 sg13g2_o21ai_1 _14806_ (.B1(_08370_),
    .Y(_00014_),
    .A1(_08289_),
    .A2(_08368_));
 sg13g2_buf_16 clkbuf_leaf_512_clk (.X(clknet_leaf_512_clk),
    .A(clknet_8_211_0_clk));
 sg13g2_buf_16 clkbuf_leaf_511_clk (.X(clknet_leaf_511_clk),
    .A(clknet_8_211_0_clk));
 sg13g2_buf_16 clkbuf_leaf_509_clk (.X(clknet_leaf_509_clk),
    .A(clknet_8_217_0_clk));
 sg13g2_nand4_1 _14810_ (.B(net10714),
    .C(_08287_),
    .A(net11052),
    .Y(_08374_),
    .D(_08348_));
 sg13g2_or3_1 _14811_ (.A(\u_ac_controller_soc_inst.u_picorv32.is_sb_sh_sw ),
    .B(\u_ac_controller_soc_inst.u_picorv32.is_sll_srl_sra ),
    .C(_08351_),
    .X(_08375_));
 sg13g2_buf_16 clkbuf_leaf_508_clk (.X(clknet_leaf_508_clk),
    .A(clknet_8_214_0_clk));
 sg13g2_buf_16 clkbuf_leaf_507_clk (.X(clknet_leaf_507_clk),
    .A(clknet_8_217_0_clk));
 sg13g2_nand2_1 _14814_ (.Y(_08378_),
    .A(net11052),
    .B(\u_ac_controller_soc_inst.u_picorv32.cpu_state[3] ));
 sg13g2_nor2_1 _14815_ (.A(_00102_),
    .B(_08378_),
    .Y(_08379_));
 sg13g2_nand3_1 _14816_ (.B(_08287_),
    .C(_08379_),
    .A(_07956_),
    .Y(_08380_));
 sg13g2_nand3_1 _14817_ (.B(_08375_),
    .C(_08380_),
    .A(_08374_),
    .Y(_00013_));
 sg13g2_buf_16 clkbuf_leaf_506_clk (.X(clknet_leaf_506_clk),
    .A(clknet_8_216_0_clk));
 sg13g2_buf_16 clkbuf_leaf_505_clk (.X(clknet_leaf_505_clk),
    .A(clknet_8_216_0_clk));
 sg13g2_buf_16 clkbuf_leaf_502_clk (.X(clknet_leaf_502_clk),
    .A(clknet_8_197_0_clk));
 sg13g2_inv_1 _14821_ (.Y(_08384_),
    .A(_08287_));
 sg13g2_nor4_1 _14822_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_jal ),
    .B(_00107_),
    .C(_08384_),
    .D(_08332_),
    .Y(_00012_));
 sg13g2_inv_1 _14823_ (.Y(_00045_),
    .A(_08308_));
 sg13g2_or3_1 _14824_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_slt ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_slti ),
    .C(\u_ac_controller_soc_inst.u_picorv32.instr_blt ),
    .X(_00046_));
 sg13g2_or3_1 _14825_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_sltu ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_sltiu ),
    .C(\u_ac_controller_soc_inst.u_picorv32.instr_bltu ),
    .X(_00047_));
 sg13g2_buf_16 clkbuf_leaf_501_clk (.X(clknet_leaf_501_clk),
    .A(clknet_8_199_0_clk));
 sg13g2_buf_16 clkbuf_leaf_498_clk (.X(clknet_leaf_498_clk),
    .A(clknet_8_199_0_clk));
 sg13g2_nand4_1 _14828_ (.B(_00085_),
    .C(_08326_),
    .A(net11051),
    .Y(_08387_),
    .D(_07972_));
 sg13g2_buf_16 clkbuf_leaf_497_clk (.X(clknet_leaf_497_clk),
    .A(clknet_8_204_0_clk));
 sg13g2_buf_16 clkbuf_leaf_496_clk (.X(clknet_leaf_496_clk),
    .A(clknet_8_205_0_clk));
 sg13g2_inv_4 _14831_ (.A(net10714),
    .Y(_08390_));
 sg13g2_buf_16 clkbuf_leaf_495_clk (.X(clknet_leaf_495_clk),
    .A(clknet_8_205_0_clk));
 sg13g2_buf_16 clkbuf_leaf_493_clk (.X(clknet_leaf_493_clk),
    .A(clknet_8_205_0_clk));
 sg13g2_buf_16 clkbuf_leaf_492_clk (.X(clknet_leaf_492_clk),
    .A(clknet_8_204_0_clk));
 sg13g2_o21ai_1 _14835_ (.B1(net10660),
    .Y(_08394_),
    .A1(_00107_),
    .A2(_00108_));
 sg13g2_inv_8 _14836_ (.Y(_08395_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[3] ));
 sg13g2_buf_16 clkbuf_leaf_491_clk (.X(clknet_leaf_491_clk),
    .A(clknet_8_198_0_clk));
 sg13g2_o21ai_1 _14838_ (.B1(net11051),
    .Y(_08397_),
    .A1(_08395_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.is_beq_bne_blt_bge_bltu_bgeu ));
 sg13g2_buf_16 clkbuf_leaf_490_clk (.X(clknet_leaf_490_clk),
    .A(clknet_8_199_0_clk));
 sg13g2_a21oi_1 _14840_ (.A1(net10722),
    .A2(_08394_),
    .Y(_08399_),
    .B1(_08397_));
 sg13g2_o21ai_1 _14841_ (.B1(_08399_),
    .Y(_08400_),
    .A1(_08390_),
    .A2(_08322_));
 sg13g2_a221oi_1 _14842_ (.B2(_08326_),
    .C1(_08400_),
    .B1(_08379_),
    .A1(net10708),
    .Y(_08401_),
    .A2(_08365_));
 sg13g2_a22oi_1 _14843_ (.Y(_00011_),
    .B1(_08387_),
    .B2(_08401_),
    .A2(_08384_),
    .A1(net11051));
 sg13g2_buf_16 clkbuf_leaf_489_clk (.X(clknet_leaf_489_clk),
    .A(clknet_8_197_0_clk));
 sg13g2_buf_16 clkbuf_leaf_488_clk (.X(clknet_leaf_488_clk),
    .A(clknet_8_197_0_clk));
 sg13g2_buf_16 clkbuf_leaf_487_clk (.X(clknet_leaf_487_clk),
    .A(clknet_8_197_0_clk));
 sg13g2_nand2b_1 _14847_ (.Y(_08405_),
    .B(_08287_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.cpu_state[0] ));
 sg13g2_a21oi_1 _14848_ (.A1(net10714),
    .A2(_08324_),
    .Y(_08406_),
    .B1(_08405_));
 sg13g2_nor2_1 _14849_ (.A(net11014),
    .B(_08406_),
    .Y(_00010_));
 sg13g2_inv_1 _14850_ (.Y(_08407_),
    .A(\u_ac_controller_soc_inst.io_rdata[0] ));
 sg13g2_nand2_2 _14851_ (.Y(_08408_),
    .A(_07701_),
    .B(_07924_));
 sg13g2_buf_16 clkbuf_leaf_486_clk (.X(clknet_leaf_486_clk),
    .A(clknet_8_198_0_clk));
 sg13g2_nand4_1 _14853_ (.B(_07926_),
    .C(_07895_),
    .A(_07899_),
    .Y(_08410_),
    .D(_07901_));
 sg13g2_buf_16 clkbuf_leaf_485_clk (.X(clknet_leaf_485_clk),
    .A(clknet_8_196_0_clk));
 sg13g2_nor2_2 _14855_ (.A(net10606),
    .B(_08410_),
    .Y(_08412_));
 sg13g2_and2_1 _14856_ (.A(\u_ac_controller_soc_inst.spi_sensor_rdata[0] ),
    .B(_07887_),
    .X(_08413_));
 sg13g2_a221oi_1 _14857_ (.B2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[0] ),
    .C1(_08413_),
    .B1(_08412_),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[0] ),
    .Y(_08414_),
    .A2(_07979_));
 sg13g2_o21ai_1 _14858_ (.B1(_08414_),
    .Y(_08415_),
    .A1(_08407_),
    .A2(net10186));
 sg13g2_buf_16 clkbuf_leaf_482_clk (.X(clknet_leaf_482_clk),
    .A(clknet_8_196_0_clk));
 sg13g2_nor2_2 _14860_ (.A(_00086_),
    .B(_07935_),
    .Y(_08417_));
 sg13g2_buf_16 clkbuf_leaf_481_clk (.X(clknet_leaf_481_clk),
    .A(clknet_8_196_0_clk));
 sg13g2_buf_16 clkbuf_leaf_478_clk (.X(clknet_leaf_478_clk),
    .A(clknet_8_196_0_clk));
 sg13g2_mux2_1 _14863_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[0] ),
    .A1(_08415_),
    .S(net9804),
    .X(_00113_));
 sg13g2_and2_1 _14864_ (.A(_07701_),
    .B(_07924_),
    .X(_08420_));
 sg13g2_buf_16 clkbuf_leaf_477_clk (.X(clknet_leaf_477_clk),
    .A(clknet_8_208_0_clk));
 sg13g2_nand2_1 _14866_ (.Y(_08422_),
    .A(\u_ac_controller_soc_inst.io_rdata[1] ),
    .B(net10184));
 sg13g2_buf_16 clkbuf_leaf_475_clk (.X(clknet_leaf_475_clk),
    .A(clknet_8_208_0_clk));
 sg13g2_a22oi_1 _14868_ (.Y(_08424_),
    .B1(_07931_),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[1] ),
    .A2(net10230),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[1] ));
 sg13g2_and2_1 _14869_ (.A(_07701_),
    .B(_07927_),
    .X(_08425_));
 sg13g2_buf_16 clkbuf_leaf_474_clk (.X(clknet_leaf_474_clk),
    .A(clknet_8_110_0_clk));
 sg13g2_nand2_1 _14871_ (.Y(_08427_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[1] ),
    .B(_08425_));
 sg13g2_nand3_1 _14872_ (.B(_08424_),
    .C(_08427_),
    .A(_08422_),
    .Y(_08428_));
 sg13g2_mux2_1 _14873_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[1] ),
    .A1(_08428_),
    .S(net9804),
    .X(_00114_));
 sg13g2_buf_16 clkbuf_leaf_473_clk (.X(clknet_leaf_473_clk),
    .A(clknet_8_107_0_clk));
 sg13g2_buf_16 clkbuf_leaf_472_clk (.X(clknet_leaf_472_clk),
    .A(clknet_8_193_0_clk));
 sg13g2_inv_2 _14876_ (.Y(_08431_),
    .A(\u_ac_controller_soc_inst.spi_flash_rdata[2] ));
 sg13g2_a22oi_1 _14877_ (.Y(_08432_),
    .B1(_08412_),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[2] ),
    .A2(_07887_),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[2] ));
 sg13g2_o21ai_1 _14878_ (.B1(_08432_),
    .Y(_08433_),
    .A1(_08431_),
    .A2(_07744_));
 sg13g2_a21oi_2 _14879_ (.B1(_08433_),
    .Y(_08434_),
    .A2(net10184),
    .A1(\u_ac_controller_soc_inst.io_rdata[2] ));
 sg13g2_nand2_1 _14880_ (.Y(_08435_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[2] ),
    .B(net9811));
 sg13g2_o21ai_1 _14881_ (.B1(_08435_),
    .Y(_00115_),
    .A1(net9810),
    .A2(_08434_));
 sg13g2_inv_2 _14882_ (.Y(_08436_),
    .A(\u_ac_controller_soc_inst.spi_flash_rdata[3] ));
 sg13g2_a22oi_1 _14883_ (.Y(_08437_),
    .B1(_08412_),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[3] ),
    .A2(_07887_),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[3] ));
 sg13g2_o21ai_1 _14884_ (.B1(_08437_),
    .Y(_08438_),
    .A1(_08436_),
    .A2(_07744_));
 sg13g2_a21oi_2 _14885_ (.B1(_08438_),
    .Y(_08439_),
    .A2(net10184),
    .A1(\u_ac_controller_soc_inst.io_rdata[3] ));
 sg13g2_nand2_1 _14886_ (.Y(_08440_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[3] ),
    .B(net9810));
 sg13g2_o21ai_1 _14887_ (.B1(_08440_),
    .Y(_08441_),
    .A1(net9810),
    .A2(_08439_));
 sg13g2_buf_16 clkbuf_leaf_470_clk (.X(clknet_leaf_470_clk),
    .A(clknet_8_107_0_clk));
 sg13g2_buf_16 clkbuf_leaf_469_clk (.X(clknet_leaf_469_clk),
    .A(clknet_8_107_0_clk));
 sg13g2_buf_16 clkbuf_leaf_467_clk (.X(clknet_leaf_467_clk),
    .A(clknet_8_192_0_clk));
 sg13g2_mux2_1 _14891_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.config_clk ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk ),
    .S(net10486),
    .X(spi_flash_clk));
 sg13g2_nand2_1 _14892_ (.Y(_08444_),
    .A(\u_ac_controller_soc_inst.io_rdata[4] ),
    .B(net10184));
 sg13g2_buf_16 clkbuf_leaf_466_clk (.X(clknet_leaf_466_clk),
    .A(clknet_8_192_0_clk));
 sg13g2_a22oi_1 _14894_ (.Y(_08446_),
    .B1(_07931_),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[4] ),
    .A2(net10230),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[4] ));
 sg13g2_nand2_1 _14895_ (.Y(_08447_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[4] ),
    .B(_08425_));
 sg13g2_nand3_1 _14896_ (.B(_08446_),
    .C(_08447_),
    .A(_08444_),
    .Y(_08448_));
 sg13g2_mux2_1 _14897_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[4] ),
    .A1(_08448_),
    .S(net9804),
    .X(_08449_));
 sg13g2_buf_16 clkbuf_leaf_465_clk (.X(clknet_leaf_465_clk),
    .A(clknet_8_192_0_clk));
 sg13g2_mux2_1 _14899_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.config_csb ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_csb ),
    .S(net10486),
    .X(spi_flash_cs_n));
 sg13g2_nand2_1 _14900_ (.Y(_08450_),
    .A(\u_ac_controller_soc_inst.io_rdata[5] ),
    .B(net10184));
 sg13g2_buf_16 clkbuf_leaf_464_clk (.X(clknet_leaf_464_clk),
    .A(clknet_8_192_0_clk));
 sg13g2_a22oi_1 _14902_ (.Y(_08452_),
    .B1(net10242),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[5] ),
    .A2(net10231),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[5] ));
 sg13g2_nand2_1 _14903_ (.Y(_08453_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[5] ),
    .B(_08425_));
 sg13g2_nand3_1 _14904_ (.B(_08452_),
    .C(_08453_),
    .A(_08450_),
    .Y(_08454_));
 sg13g2_mux2_1 _14905_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[5] ),
    .A1(_08454_),
    .S(net9804),
    .X(_08455_));
 sg13g2_buf_16 clkbuf_leaf_463_clk (.X(clknet_leaf_463_clk),
    .A(clknet_8_195_0_clk));
 sg13g2_nand2_1 _14907_ (.Y(_08456_),
    .A(\u_ac_controller_soc_inst.io_rdata[6] ),
    .B(net10184));
 sg13g2_a22oi_1 _14908_ (.Y(_08457_),
    .B1(_07931_),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[6] ),
    .A2(net10230),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[6] ));
 sg13g2_nand2_1 _14909_ (.Y(_08458_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[6] ),
    .B(_08425_));
 sg13g2_nand3_1 _14910_ (.B(_08457_),
    .C(_08458_),
    .A(_08456_),
    .Y(_08459_));
 sg13g2_mux2_1 _14911_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[6] ),
    .A1(_08459_),
    .S(net9804),
    .X(_08460_));
 sg13g2_buf_16 clkbuf_leaf_461_clk (.X(clknet_leaf_461_clk),
    .A(clknet_8_194_0_clk));
 sg13g2_buf_16 clkbuf_leaf_457_clk (.X(clknet_leaf_457_clk),
    .A(clknet_8_245_0_clk));
 sg13g2_buf_16 clkbuf_leaf_456_clk (.X(clknet_leaf_456_clk),
    .A(clknet_8_244_0_clk));
 sg13g2_and2_1 _14915_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[13] ),
    .B(net10232),
    .X(_08463_));
 sg13g2_a221oi_1 _14916_ (.B2(\u_ac_controller_soc_inst.io_rdata[13] ),
    .C1(_08463_),
    .B1(net10183),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[13] ),
    .Y(_08464_),
    .A2(net10242));
 sg13g2_buf_16 clkbuf_leaf_455_clk (.X(clknet_leaf_455_clk),
    .A(clknet_8_244_0_clk));
 sg13g2_buf_16 clkbuf_leaf_453_clk (.X(clknet_leaf_453_clk),
    .A(clknet_8_31_0_clk));
 sg13g2_nand2_1 _14919_ (.Y(_08467_),
    .A(net10607),
    .B(net9811));
 sg13g2_o21ai_1 _14920_ (.B1(_08467_),
    .Y(_08468_),
    .A1(net9811),
    .A2(_08464_));
 sg13g2_buf_16 clkbuf_leaf_452_clk (.X(clknet_leaf_452_clk),
    .A(clknet_8_106_0_clk));
 sg13g2_and2_1 _14922_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[12] ),
    .B(net10232),
    .X(_08469_));
 sg13g2_a221oi_1 _14923_ (.B2(\u_ac_controller_soc_inst.io_rdata[12] ),
    .C1(_08469_),
    .B1(net10183),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[12] ),
    .Y(_08470_),
    .A2(net10242));
 sg13g2_buf_16 clkbuf_leaf_450_clk (.X(clknet_leaf_450_clk),
    .A(clknet_8_104_0_clk));
 sg13g2_buf_16 clkbuf_leaf_447_clk (.X(clknet_leaf_447_clk),
    .A(clknet_8_104_0_clk));
 sg13g2_nand2_1 _14926_ (.Y(_08473_),
    .A(net10608),
    .B(net9811));
 sg13g2_o21ai_1 _14927_ (.B1(_08473_),
    .Y(_08474_),
    .A1(net9811),
    .A2(_08470_));
 sg13g2_buf_16 clkbuf_leaf_446_clk (.X(clknet_leaf_446_clk),
    .A(clknet_8_98_0_clk));
 sg13g2_and2_1 _14929_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[14] ),
    .B(net10232),
    .X(_08475_));
 sg13g2_a221oi_1 _14930_ (.B2(\u_ac_controller_soc_inst.io_rdata[14] ),
    .C1(_08475_),
    .B1(net10185),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[14] ),
    .Y(_08476_),
    .A2(net10244));
 sg13g2_buf_16 clkbuf_leaf_445_clk (.X(clknet_leaf_445_clk),
    .A(clknet_8_98_0_clk));
 sg13g2_buf_16 clkbuf_leaf_444_clk (.X(clknet_leaf_444_clk),
    .A(clknet_8_98_0_clk));
 sg13g2_nand2_1 _14933_ (.Y(_08479_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[14] ),
    .B(net9811));
 sg13g2_o21ai_1 _14934_ (.B1(_08479_),
    .Y(_08480_),
    .A1(net9811),
    .A2(_08476_));
 sg13g2_buf_16 clkbuf_leaf_443_clk (.X(clknet_leaf_443_clk),
    .A(clknet_8_99_0_clk));
 sg13g2_inv_4 _14936_ (.A(\u_ac_controller_soc_inst.io_rdata[15] ),
    .Y(_08481_));
 sg13g2_a22oi_1 _14937_ (.Y(_08482_),
    .B1(net10245),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[15] ),
    .A2(net10233),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[15] ));
 sg13g2_o21ai_1 _14938_ (.B1(_08482_),
    .Y(_08483_),
    .A1(_08481_),
    .A2(_08408_));
 sg13g2_buf_16 clkbuf_leaf_442_clk (.X(clknet_leaf_442_clk),
    .A(clknet_8_99_0_clk));
 sg13g2_mux2_1 _14940_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[15] ),
    .A1(_08483_),
    .S(net9805),
    .X(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[15] ));
 sg13g2_buf_16 clkbuf_leaf_440_clk (.X(clknet_leaf_440_clk),
    .A(clknet_8_99_0_clk));
 sg13g2_nor2_1 _14942_ (.A(_07917_),
    .B(_07936_),
    .Y(_08486_));
 sg13g2_nand2_1 _14943_ (.Y(_08487_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_state[0] ),
    .B(_08486_));
 sg13g2_o21ai_1 _14944_ (.B1(\u_ac_controller_soc_inst.u_picorv32.mem_state[1] ),
    .Y(_08488_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_state[0] ),
    .A2(_08486_));
 sg13g2_nand2b_1 _14945_ (.Y(_08489_),
    .B(net11048),
    .A_N(_00087_));
 sg13g2_a21oi_2 _14946_ (.B1(_08489_),
    .Y(_08490_),
    .A2(_08488_),
    .A1(_08487_));
 sg13g2_buf_16 clkbuf_leaf_439_clk (.X(clknet_leaf_439_clk),
    .A(clknet_8_105_0_clk));
 sg13g2_buf_16 clkbuf_leaf_438_clk (.X(clknet_leaf_438_clk),
    .A(clknet_8_104_0_clk));
 sg13g2_mux2_1 _14949_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[15] ),
    .S(net9701),
    .X(_00038_));
 sg13g2_buf_16 clkbuf_leaf_437_clk (.X(clknet_leaf_437_clk),
    .A(clknet_8_106_0_clk));
 sg13g2_and2_1 _14951_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[16] ),
    .B(net10232),
    .X(_08494_));
 sg13g2_a221oi_1 _14952_ (.B2(\u_ac_controller_soc_inst.io_rdata[16] ),
    .C1(_08494_),
    .B1(net10185),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[16] ),
    .Y(_08495_),
    .A2(net10244));
 sg13g2_buf_16 clkbuf_leaf_436_clk (.X(clknet_leaf_436_clk),
    .A(clknet_8_104_0_clk));
 sg13g2_buf_16 clkbuf_leaf_435_clk (.X(clknet_leaf_435_clk),
    .A(clknet_8_105_0_clk));
 sg13g2_nand2_1 _14955_ (.Y(_08498_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[16] ),
    .B(net9808));
 sg13g2_o21ai_1 _14956_ (.B1(_08498_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[16] ),
    .A1(net9808),
    .A2(_08495_));
 sg13g2_buf_16 clkbuf_leaf_434_clk (.X(clknet_leaf_434_clk),
    .A(clknet_8_107_0_clk));
 sg13g2_inv_2 _14958_ (.Y(_08500_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[16] ));
 sg13g2_buf_16 clkbuf_leaf_433_clk (.X(clknet_leaf_433_clk),
    .A(clknet_8_103_0_clk));
 sg13g2_buf_16 clkbuf_leaf_432_clk (.X(clknet_leaf_432_clk),
    .A(clknet_8_108_0_clk));
 sg13g2_nand2_1 _14961_ (.Y(_08503_),
    .A(net9700),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[16] ));
 sg13g2_o21ai_1 _14962_ (.B1(_08503_),
    .Y(_00039_),
    .A1(_08500_),
    .A2(net9701));
 sg13g2_inv_2 _14963_ (.Y(_08504_),
    .A(\u_ac_controller_soc_inst.io_rdata[17] ));
 sg13g2_a22oi_1 _14964_ (.Y(_08505_),
    .B1(net10245),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[17] ),
    .A2(net10233),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[17] ));
 sg13g2_o21ai_1 _14965_ (.B1(_08505_),
    .Y(_08506_),
    .A1(_08504_),
    .A2(_08408_));
 sg13g2_mux2_1 _14966_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[17] ),
    .A1(_08506_),
    .S(net9805),
    .X(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[17] ));
 sg13g2_buf_16 clkbuf_leaf_430_clk (.X(clknet_leaf_430_clk),
    .A(clknet_8_103_0_clk));
 sg13g2_mux2_1 _14968_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[17] ),
    .S(net9701),
    .X(_00040_));
 sg13g2_buf_16 clkbuf_leaf_429_clk (.X(clknet_leaf_429_clk),
    .A(clknet_8_102_0_clk));
 sg13g2_and2_1 _14970_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[18] ),
    .B(net10233),
    .X(_08509_));
 sg13g2_a221oi_1 _14971_ (.B2(\u_ac_controller_soc_inst.io_rdata[18] ),
    .C1(_08509_),
    .B1(net10185),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[18] ),
    .Y(_08510_),
    .A2(net10245));
 sg13g2_buf_16 clkbuf_leaf_428_clk (.X(clknet_leaf_428_clk),
    .A(clknet_8_102_0_clk));
 sg13g2_nand2_1 _14973_ (.Y(_08512_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[18] ),
    .B(net9808));
 sg13g2_o21ai_1 _14974_ (.B1(_08512_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[18] ),
    .A1(net9808),
    .A2(_08510_));
 sg13g2_buf_16 clkbuf_leaf_427_clk (.X(clknet_leaf_427_clk),
    .A(clknet_8_102_0_clk));
 sg13g2_mux2_1 _14976_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[18] ),
    .S(net9701),
    .X(_00041_));
 sg13g2_and2_1 _14977_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[19] ),
    .B(net10233),
    .X(_08514_));
 sg13g2_a221oi_1 _14978_ (.B2(\u_ac_controller_soc_inst.io_rdata[19] ),
    .C1(_08514_),
    .B1(net10185),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[19] ),
    .Y(_08515_),
    .A2(net10245));
 sg13g2_buf_16 clkbuf_leaf_426_clk (.X(clknet_leaf_426_clk),
    .A(clknet_8_102_0_clk));
 sg13g2_nand2_1 _14980_ (.Y(_08517_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[19] ),
    .B(net9808));
 sg13g2_o21ai_1 _14981_ (.B1(_08517_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[19] ),
    .A1(net9808),
    .A2(_08515_));
 sg13g2_inv_1 _14982_ (.Y(_08518_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[19] ));
 sg13g2_nand2_1 _14983_ (.Y(_08519_),
    .A(net9701),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[19] ));
 sg13g2_o21ai_1 _14984_ (.B1(_08519_),
    .Y(_00042_),
    .A1(_08518_),
    .A2(net9701));
 sg13g2_a22oi_1 _14985_ (.Y(_08520_),
    .B1(net10245),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[20] ),
    .A2(net10233),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[20] ));
 sg13g2_nand2_1 _14986_ (.Y(_08521_),
    .A(\u_ac_controller_soc_inst.io_rdata[20] ),
    .B(net10183));
 sg13g2_and2_1 _14987_ (.A(_08520_),
    .B(_08521_),
    .X(_08522_));
 sg13g2_buf_16 clkbuf_leaf_425_clk (.X(clknet_leaf_425_clk),
    .A(clknet_8_99_0_clk));
 sg13g2_buf_16 clkbuf_leaf_424_clk (.X(clknet_leaf_424_clk),
    .A(clknet_8_79_0_clk));
 sg13g2_nand2_1 _14990_ (.Y(_08525_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[20] ),
    .B(net9808));
 sg13g2_o21ai_1 _14991_ (.B1(_08525_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[20] ),
    .A1(net9808),
    .A2(_08522_));
 sg13g2_buf_16 clkbuf_leaf_422_clk (.X(clknet_leaf_422_clk),
    .A(clknet_8_103_0_clk));
 sg13g2_inv_2 _14993_ (.Y(_08527_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11] ));
 sg13g2_nand2_1 _14994_ (.Y(_08528_),
    .A(net9700),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[20] ));
 sg13g2_o21ai_1 _14995_ (.B1(_08528_),
    .Y(_00033_),
    .A1(_08527_),
    .A2(net9702));
 sg13g2_a22oi_1 _14996_ (.Y(_08529_),
    .B1(net10243),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[21] ),
    .A2(net10230),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[21] ));
 sg13g2_nand2_1 _14997_ (.Y(_08530_),
    .A(\u_ac_controller_soc_inst.io_rdata[21] ),
    .B(net10183));
 sg13g2_and2_1 _14998_ (.A(_08529_),
    .B(_08530_),
    .X(_08531_));
 sg13g2_buf_16 clkbuf_leaf_421_clk (.X(clknet_leaf_421_clk),
    .A(clknet_8_101_0_clk));
 sg13g2_buf_16 clkbuf_leaf_420_clk (.X(clknet_leaf_420_clk),
    .A(clknet_8_101_0_clk));
 sg13g2_nand2_1 _15001_ (.Y(_08534_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[21] ),
    .B(net9807));
 sg13g2_o21ai_1 _15002_ (.B1(_08534_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[21] ),
    .A1(net9807),
    .A2(_08531_));
 sg13g2_buf_16 clkbuf_leaf_419_clk (.X(clknet_leaf_419_clk),
    .A(clknet_8_90_0_clk));
 sg13g2_mux2_1 _15004_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[21] ),
    .S(net9702),
    .X(_00034_));
 sg13g2_and2_1 _15005_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[22] ),
    .B(net10233),
    .X(_08536_));
 sg13g2_a221oi_1 _15006_ (.B2(\u_ac_controller_soc_inst.io_rdata[22] ),
    .C1(_08536_),
    .B1(net10185),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[22] ),
    .Y(_08537_),
    .A2(net10245));
 sg13g2_buf_16 clkbuf_leaf_417_clk (.X(clknet_leaf_417_clk),
    .A(clknet_8_90_0_clk));
 sg13g2_buf_2 place9645 (.A(_10033_),
    .X(net9645));
 sg13g2_nand2_1 _15009_ (.Y(_08540_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[22] ),
    .B(net9809));
 sg13g2_o21ai_1 _15010_ (.B1(_08540_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[22] ),
    .A1(net9809),
    .A2(_08537_));
 sg13g2_buf_2 place9648 (.A(net9647),
    .X(net9648));
 sg13g2_mux2_1 _15012_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[22] ),
    .S(net9704),
    .X(_00035_));
 sg13g2_and2_1 _15013_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[23] ),
    .B(net10233),
    .X(_08542_));
 sg13g2_a221oi_1 _15014_ (.B2(\u_ac_controller_soc_inst.io_rdata[23] ),
    .C1(_08542_),
    .B1(_08420_),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[23] ),
    .Y(_08543_),
    .A2(net10244));
 sg13g2_buf_2 place9679 (.A(net9678),
    .X(net9679));
 sg13g2_buf_2 place9646 (.A(net9645),
    .X(net9646));
 sg13g2_nand2_1 _15017_ (.Y(_08546_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[23] ),
    .B(net9806));
 sg13g2_o21ai_1 _15018_ (.B1(_08546_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[23] ),
    .A1(net9806),
    .A2(_08543_));
 sg13g2_buf_2 place9670 (.A(net9665),
    .X(net9670));
 sg13g2_inv_2 _15020_ (.Y(_08548_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3] ));
 sg13g2_nand2_1 _15021_ (.Y(_08549_),
    .A(net9704),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[23] ));
 sg13g2_o21ai_1 _15022_ (.B1(_08549_),
    .Y(_00036_),
    .A1(_08548_),
    .A2(net9704));
 sg13g2_buf_2 place9636 (.A(net9635),
    .X(net9636));
 sg13g2_inv_2 _15024_ (.Y(_08551_),
    .A(\u_ac_controller_soc_inst.io_rdata[24] ));
 sg13g2_a22oi_1 _15025_ (.Y(_08552_),
    .B1(net10243),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[24] ),
    .A2(net10230),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[24] ));
 sg13g2_o21ai_1 _15026_ (.B1(_08552_),
    .Y(_08553_),
    .A1(_08551_),
    .A2(net10186));
 sg13g2_mux2_1 _15027_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[24] ),
    .A1(_08553_),
    .S(_08417_),
    .X(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[24] ));
 sg13g2_buf_2 place10827 (.A(_00000_),
    .X(net10827));
 sg13g2_mux2_1 _15029_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[24] ),
    .S(net9704),
    .X(_00037_));
 sg13g2_buf_2 place10845 (.A(_00000_),
    .X(net10845));
 sg13g2_buf_2 place9644 (.A(net9643),
    .X(net9644));
 sg13g2_nor2b_1 _15032_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[4] ),
    .B_N(net10464),
    .Y(_08557_));
 sg13g2_buf_2 place9642 (.A(net9641),
    .X(net9642));
 sg13g2_inv_1 _15034_ (.Y(_08559_),
    .A(_00124_));
 sg13g2_nor2_2 _15035_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr ),
    .Y(_08560_));
 sg13g2_a221oi_1 _15036_ (.B2(_08560_),
    .C1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_qspi ),
    .B1(_08559_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi ),
    .Y(_08561_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[6] ));
 sg13g2_nor3_2 _15037_ (.A(_08204_),
    .B(_08557_),
    .C(_08561_),
    .Y(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io0_do ));
 sg13g2_nor2_1 _15038_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi ),
    .B(net10465),
    .Y(_08562_));
 sg13g2_nor4_2 _15039_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[0] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[1] ),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[3] ),
    .Y(_08563_),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[2] ));
 sg13g2_nand2b_2 _15040_ (.Y(_08564_),
    .B(_08563_),
    .A_N(_08562_));
 sg13g2_buf_2 place9643 (.A(_10041_),
    .X(net9643));
 sg13g2_nor2b_1 _15042_ (.A(net10464),
    .B_N(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[7] ),
    .Y(_08566_));
 sg13g2_a21oi_2 _15043_ (.B1(_08566_),
    .Y(_08567_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[5] ),
    .A1(net10464));
 sg13g2_nor2_1 _15044_ (.A(_08564_),
    .B(_08567_),
    .Y(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io1_do ));
 sg13g2_buf_2 place9641 (.A(_10041_),
    .X(net9641));
 sg13g2_and3_2 _15046_ (.X(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io2_do ),
    .A(net10464),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[6] ),
    .C(_08563_));
 sg13g2_nand2_1 _15047_ (.Y(_08569_),
    .A(net10464),
    .B(_08563_));
 sg13g2_nor2_1 _15048_ (.A(_00124_),
    .B(_08569_),
    .Y(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io3_do ));
 sg13g2_inv_1 _15049_ (.Y(_08570_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[0] ));
 sg13g2_a21oi_2 _15050_ (.B1(_08204_),
    .Y(_08571_),
    .A2(_08562_),
    .A1(net10466));
 sg13g2_buf_16 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_8_1_0_clk));
 sg13g2_buf_2 place9934 (.A(net9933),
    .X(net9934));
 sg13g2_o21ai_1 _15053_ (.B1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_rd ),
    .Y(_08574_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi ),
    .A2(net10465));
 sg13g2_nand3_1 _15054_ (.B(_08571_),
    .C(_08574_),
    .A(net10485),
    .Y(_08575_));
 sg13g2_o21ai_1 _15055_ (.B1(_08575_),
    .Y(spi_flash_io0_oe),
    .A1(net10486),
    .A2(_08570_));
 sg13g2_nor2_1 _15056_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_rd ),
    .B(_08564_),
    .Y(_08576_));
 sg13g2_mux2_1 _15057_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[1] ),
    .A1(_08576_),
    .S(net10486),
    .X(spi_flash_io1_oe));
 sg13g2_inv_1 _15058_ (.Y(_08577_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[2] ));
 sg13g2_inv_1 _15059_ (.Y(_08578_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_rd ));
 sg13g2_nand4_1 _15060_ (.B(_08578_),
    .C(net10485),
    .A(net10465),
    .Y(_08579_),
    .D(_08563_));
 sg13g2_o21ai_1 _15061_ (.B1(_08579_),
    .Y(spi_flash_io2_oe),
    .A1(net10485),
    .A2(_08577_));
 sg13g2_inv_1 _15062_ (.Y(_08580_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[3] ));
 sg13g2_o21ai_1 _15063_ (.B1(_08579_),
    .Y(spi_flash_io3_oe),
    .A1(net10485),
    .A2(_08580_));
 sg13g2_a21o_2 _15064_ (.A2(_08488_),
    .A1(_08487_),
    .B1(_08489_),
    .X(_08581_));
 sg13g2_buf_2 place9725 (.A(net9723),
    .X(net9725));
 sg13g2_buf_2 place11054 (.A(net11037),
    .X(net11054));
 sg13g2_inv_1 _15067_ (.Y(_08584_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_slti_blt_slt ));
 sg13g2_buf_2 place10944 (.A(net10939),
    .X(net10944));
 sg13g2_inv_8 _15069_ (.Y(_08586_),
    .A(net10533));
 sg13g2_buf_2 place9708 (.A(_04607_),
    .X(net9708));
 sg13g2_buf_2 place9771 (.A(_04955_),
    .X(net9771));
 sg13g2_nor2b_1 _15072_ (.A(net10537),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[30] ),
    .Y(_08589_));
 sg13g2_nand2b_2 _15073_ (.Y(_08590_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[30] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[30] ));
 sg13g2_nand2b_2 _15074_ (.Y(_08591_),
    .B(_08590_),
    .A_N(_08589_));
 sg13g2_buf_2 place9703 (.A(net9702),
    .X(net9703));
 sg13g2_xor2_1 _15076_ (.B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[31] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[31] ),
    .X(_08593_));
 sg13g2_buf_2 place10937 (.A(net10936),
    .X(net10937));
 sg13g2_buf_2 place10938 (.A(net10937),
    .X(net10938));
 sg13g2_buf_2 place10943 (.A(net10942),
    .X(net10943));
 sg13g2_xor2_1 _15080_ (.B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[28] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[28] ),
    .X(_08597_));
 sg13g2_buf_2 place10936 (.A(net10935),
    .X(net10936));
 sg13g2_buf_2 place10974 (.A(net10973),
    .X(net10974));
 sg13g2_xor2_1 _15083_ (.B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[29] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[29] ),
    .X(_08600_));
 sg13g2_or4_1 _15084_ (.A(_08591_),
    .B(_08593_),
    .C(_08597_),
    .D(_08600_),
    .X(_08601_));
 sg13g2_buf_2 place10957 (.A(net10953),
    .X(net10957));
 sg13g2_buf_2 place10891 (.A(net10890),
    .X(net10891));
 sg13g2_buf_2 place10955 (.A(net10954),
    .X(net10955));
 sg13g2_inv_4 _15088_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[26] ),
    .Y(_08605_));
 sg13g2_nor2_2 _15089_ (.A(net10509),
    .B(_08605_),
    .Y(_08606_));
 sg13g2_nand2_2 _15090_ (.Y(_08607_),
    .A(net10509),
    .B(_08605_));
 sg13g2_nand2b_2 _15091_ (.Y(_08608_),
    .B(_08607_),
    .A_N(_08606_));
 sg13g2_buf_2 place10942 (.A(net10940),
    .X(net10942));
 sg13g2_inv_2 _15093_ (.Y(_08610_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[25] ));
 sg13g2_nor2_2 _15094_ (.A(net10510),
    .B(_08610_),
    .Y(_08611_));
 sg13g2_buf_2 place10879 (.A(net10878),
    .X(net10879));
 sg13g2_buf_2 place10966 (.A(net10965),
    .X(net10966));
 sg13g2_nand2_2 _15097_ (.Y(_08614_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[25] ),
    .B(_08610_));
 sg13g2_nand2b_2 _15098_ (.Y(_08615_),
    .B(_08614_),
    .A_N(_08611_));
 sg13g2_buf_2 place10878 (.A(_00008_),
    .X(net10878));
 sg13g2_buf_2 place10890 (.A(net10888),
    .X(net10890));
 sg13g2_buf_16 clkbuf_leaf_130_clk (.X(clknet_leaf_130_clk),
    .A(clknet_8_15_0_clk));
 sg13g2_nor2b_2 _15102_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[24] ),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[24] ),
    .Y(_08619_));
 sg13g2_inv_4 _15103_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[24] ),
    .Y(_08620_));
 sg13g2_nor2_1 _15104_ (.A(_08620_),
    .B(net10555),
    .Y(_08621_));
 sg13g2_or2_1 _15105_ (.X(_08622_),
    .B(_08621_),
    .A(_08619_));
 sg13g2_buf_16 clkbuf_leaf_124_clk (.X(clknet_leaf_124_clk),
    .A(clknet_8_26_0_clk));
 sg13g2_nor3_1 _15107_ (.A(_08608_),
    .B(_08615_),
    .C(_08622_),
    .Y(_08624_));
 sg13g2_buf_2 place9627 (.A(_04222_),
    .X(net9627));
 sg13g2_buf_2 place9647 (.A(net9645),
    .X(net9647));
 sg13g2_xnor2_1 _15110_ (.Y(_08627_),
    .A(net10511),
    .B(net10558));
 sg13g2_nand2_1 _15111_ (.Y(_08628_),
    .A(_08624_),
    .B(_08627_));
 sg13g2_buf_2 place9678 (.A(_10005_),
    .X(net9678));
 sg13g2_buf_2 place9797 (.A(net9795),
    .X(net9797));
 sg13g2_xnor2_1 _15114_ (.Y(_08631_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[21] ),
    .B(net10564));
 sg13g2_buf_2 place10436 (.A(net10435),
    .X(net10436));
 sg13g2_buf_2 place9798 (.A(_09902_),
    .X(net9798));
 sg13g2_nor2b_2 _15117_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[22] ),
    .B_N(net10561),
    .Y(_08634_));
 sg13g2_buf_2 place10111 (.A(_10253_),
    .X(net10111));
 sg13g2_nor2b_2 _15119_ (.A(net10561),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[22] ),
    .Y(_08636_));
 sg13g2_buf_2 place10160 (.A(_03922_),
    .X(net10160));
 sg13g2_nor2_2 _15121_ (.A(_08634_),
    .B(_08636_),
    .Y(_08638_));
 sg13g2_buf_2 place10129 (.A(net10126),
    .X(net10129));
 sg13g2_buf_2 place9665 (.A(_11943_),
    .X(net9665));
 sg13g2_xnor2_1 _15124_ (.Y(_08641_),
    .A(net10512),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[20] ));
 sg13g2_nand3_1 _15125_ (.B(_08638_),
    .C(_08641_),
    .A(_08631_),
    .Y(_08642_));
 sg13g2_buf_2 place9688 (.A(_09997_),
    .X(net9688));
 sg13g2_buf_2 place9667 (.A(net9666),
    .X(net9667));
 sg13g2_nor2b_1 _15128_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[27] ),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[27] ),
    .Y(_08645_));
 sg13g2_nand2b_1 _15129_ (.Y(_08646_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[27] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[27] ));
 sg13g2_nand2b_2 _15130_ (.Y(_08647_),
    .B(_08646_),
    .A_N(_08645_));
 sg13g2_buf_2 place9666 (.A(net9665),
    .X(net9666));
 sg13g2_nor3_2 _15132_ (.A(_08628_),
    .B(_08642_),
    .C(_08647_),
    .Y(_08649_));
 sg13g2_buf_2 place9691 (.A(net9690),
    .X(net9691));
 sg13g2_buf_2 place9662 (.A(net9661),
    .X(net9662));
 sg13g2_nor2b_2 _15135_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[17] ),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[17] ),
    .Y(_08652_));
 sg13g2_inv_4 _15136_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[17] ),
    .Y(_08653_));
 sg13g2_nand2_1 _15137_ (.Y(_08654_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[17] ),
    .B(_08653_));
 sg13g2_nand2b_2 _15138_ (.Y(_08655_),
    .B(_08654_),
    .A_N(_08652_));
 sg13g2_buf_2 place9638 (.A(net9637),
    .X(net9638));
 sg13g2_buf_2 place9658 (.A(net9656),
    .X(net9658));
 sg13g2_buf_2 place9661 (.A(net9658),
    .X(net9661));
 sg13g2_nor2b_1 _15142_ (.A(net10574),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[19] ),
    .Y(_08659_));
 sg13g2_nand2b_2 _15143_ (.Y(_08660_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[19] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[19] ));
 sg13g2_nand2b_2 _15144_ (.Y(_08661_),
    .B(_08660_),
    .A_N(_08659_));
 sg13g2_buf_2 place9856 (.A(net9853),
    .X(net9856));
 sg13g2_buf_2 place10097 (.A(_10335_),
    .X(net10097));
 sg13g2_xor2_1 _15147_ (.B(net10576),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[18] ),
    .X(_08664_));
 sg13g2_buf_2 place9639 (.A(_10056_),
    .X(net9639));
 sg13g2_buf_2 place9640 (.A(net9639),
    .X(net9640));
 sg13g2_buf_2 place10811 (.A(_00001_),
    .X(net10811));
 sg13g2_xor2_1 _15151_ (.B(net10580),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[16] ),
    .X(_08668_));
 sg13g2_nor4_2 _15152_ (.A(_08655_),
    .B(_08661_),
    .C(_08664_),
    .Y(_08669_),
    .D(_08668_));
 sg13g2_buf_2 place9847 (.A(_11204_),
    .X(net9847));
 sg13g2_buf_2 place9852 (.A(net9849),
    .X(net9852));
 sg13g2_buf_2 place9659 (.A(net9658),
    .X(net9659));
 sg13g2_nand3b_1 _15156_ (.B(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[0] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[1] ),
    .Y(_08673_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[0] ));
 sg13g2_buf_2 place10022 (.A(net10020),
    .X(net10022));
 sg13g2_buf_2 place9660 (.A(net9658),
    .X(net9660));
 sg13g2_buf_2 place9631 (.A(net9629),
    .X(net9631));
 sg13g2_nand2b_1 _15160_ (.Y(_08677_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[2] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[2] ));
 sg13g2_nand3_1 _15161_ (.B(_08673_),
    .C(_08677_),
    .A(net10532),
    .Y(_08678_));
 sg13g2_buf_2 place9851 (.A(net9849),
    .X(net9851));
 sg13g2_inv_4 _15163_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[3] ),
    .Y(_08680_));
 sg13g2_nand3_1 _15164_ (.B(_08673_),
    .C(_08677_),
    .A(_08680_),
    .Y(_08681_));
 sg13g2_inv_1 _15165_ (.Y(_08682_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[1] ));
 sg13g2_nand2b_1 _15166_ (.Y(_08683_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[0] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[0] ));
 sg13g2_a21oi_1 _15167_ (.A1(_08682_),
    .A2(_08683_),
    .Y(_08684_),
    .B1(net10572));
 sg13g2_a21o_2 _15168_ (.A2(_08681_),
    .A1(_08678_),
    .B1(_08684_),
    .X(_08685_));
 sg13g2_buf_16 clkbuf_leaf_123_clk (.X(clknet_leaf_123_clk),
    .A(clknet_8_27_0_clk));
 sg13g2_nand2_1 _15170_ (.Y(_08687_),
    .A(_08680_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[3] ));
 sg13g2_nor2b_1 _15171_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[2] ),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[2] ),
    .Y(_08688_));
 sg13g2_o21ai_1 _15172_ (.B1(_08688_),
    .Y(_08689_),
    .A1(_08680_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[3] ));
 sg13g2_and2_1 _15173_ (.A(_08687_),
    .B(_08689_),
    .X(_08690_));
 sg13g2_buf_2 place9629 (.A(_04222_),
    .X(net9629));
 sg13g2_buf_2 place9935 (.A(net9933),
    .X(net9935));
 sg13g2_nand2b_2 _15176_ (.Y(_08693_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[5] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[5] ));
 sg13g2_buf_2 place9628 (.A(net9627),
    .X(net9628));
 sg13g2_nand2_1 _15178_ (.Y(_08695_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[4] ),
    .B(_08693_));
 sg13g2_buf_16 clkbuf_leaf_122_clk (.X(clknet_leaf_122_clk),
    .A(clknet_8_25_0_clk));
 sg13g2_nand2b_1 _15180_ (.Y(_08697_),
    .B(_08693_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[4] ));
 sg13g2_a22oi_1 _15181_ (.Y(_08698_),
    .B1(_08695_),
    .B2(_08697_),
    .A2(_08690_),
    .A1(_08685_));
 sg13g2_buf_2 place10159 (.A(net10152),
    .X(net10159));
 sg13g2_buf_16 clkbuf_leaf_94_clk (.X(clknet_leaf_94_clk),
    .A(clknet_8_59_0_clk));
 sg13g2_inv_4 _15184_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[4] ),
    .Y(_08701_));
 sg13g2_nor2_1 _15185_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[4] ),
    .B(_08701_),
    .Y(_08702_));
 sg13g2_buf_16 clkbuf_leaf_87_clk (.X(clknet_leaf_87_clk),
    .A(clknet_8_10_0_clk));
 sg13g2_nor2b_2 _15187_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[5] ),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[5] ),
    .Y(_08704_));
 sg13g2_a21oi_2 _15188_ (.B1(_08704_),
    .Y(_08705_),
    .A2(_08702_),
    .A1(_08693_));
 sg13g2_inv_4 _15189_ (.A(_08705_),
    .Y(_08706_));
 sg13g2_buf_2 place9630 (.A(net9629),
    .X(net9630));
 sg13g2_buf_16 clkbuf_leaf_121_clk (.X(clknet_leaf_121_clk),
    .A(clknet_8_24_0_clk));
 sg13g2_inv_4 _15192_ (.A(net10522),
    .Y(_08709_));
 sg13g2_buf_16 clkbuf_leaf_120_clk (.X(clknet_leaf_120_clk),
    .A(clknet_8_24_0_clk));
 sg13g2_buf_16 clkbuf_leaf_116_clk (.X(clknet_leaf_116_clk),
    .A(clknet_8_12_0_clk));
 sg13g2_nand2b_2 _15195_ (.Y(_08712_),
    .B(net10523),
    .A_N(net10500));
 sg13g2_buf_2 place10826 (.A(net10823),
    .X(net10826));
 sg13g2_nand2b_1 _15197_ (.Y(_08714_),
    .B(net10500),
    .A_N(net10523));
 sg13g2_buf_16 clkbuf_leaf_90_clk (.X(clknet_leaf_90_clk),
    .A(clknet_8_8_0_clk));
 sg13g2_inv_2 _15199_ (.Y(_08716_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[7] ));
 sg13g2_buf_2 place10245 (.A(net10244),
    .X(net10245));
 sg13g2_buf_2 place10809 (.A(net10808),
    .X(net10809));
 sg13g2_nor2b_2 _15202_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[6] ),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[6] ),
    .Y(_08719_));
 sg13g2_nand2_1 _15203_ (.Y(_08720_),
    .A(_08716_),
    .B(_08719_));
 sg13g2_buf_2 place10805 (.A(net10803),
    .X(net10805));
 sg13g2_o21ai_1 _15205_ (.B1(net10501),
    .Y(_08722_),
    .A1(_08716_),
    .A2(_08719_));
 sg13g2_nand3_1 _15206_ (.B(_08720_),
    .C(_08722_),
    .A(_08714_),
    .Y(_08723_));
 sg13g2_buf_2 place10808 (.A(_00001_),
    .X(net10808));
 sg13g2_buf_16 clkbuf_leaf_114_clk (.X(clknet_leaf_114_clk),
    .A(clknet_8_12_0_clk));
 sg13g2_buf_16 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_8_59_0_clk));
 sg13g2_xnor2_1 _15210_ (.Y(_08727_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[13] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[13] ));
 sg13g2_buf_16 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_8_58_0_clk));
 sg13g2_buf_16 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_8_2_0_clk));
 sg13g2_nand2b_2 _15213_ (.Y(_08730_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[14] ),
    .A_N(net10516));
 sg13g2_buf_16 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_8_8_0_clk));
 sg13g2_nand2b_1 _15215_ (.Y(_08732_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[14] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[14] ));
 sg13g2_and2_1 _15216_ (.A(_08730_),
    .B(_08732_),
    .X(_08733_));
 sg13g2_buf_16 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_8_51_0_clk));
 sg13g2_buf_16 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_8_49_0_clk));
 sg13g2_buf_16 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_8_2_0_clk));
 sg13g2_xor2_1 _15220_ (.B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[15] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[15] ),
    .X(_08737_));
 sg13g2_buf_16 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_8_55_0_clk));
 sg13g2_buf_16 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_8_51_0_clk));
 sg13g2_xor2_1 _15223_ (.B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[10] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[10] ),
    .X(_08740_));
 sg13g2_buf_16 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_8_57_0_clk));
 sg13g2_buf_16 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_8_51_0_clk));
 sg13g2_xor2_1 _15226_ (.B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[11] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[11] ),
    .X(_08743_));
 sg13g2_buf_16 clkbuf_leaf_113_clk (.X(clknet_leaf_113_clk),
    .A(clknet_8_26_0_clk));
 sg13g2_buf_16 clkbuf_leaf_107_clk (.X(clknet_leaf_107_clk),
    .A(clknet_8_14_0_clk));
 sg13g2_xor2_1 _15229_ (.B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[12] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[12] ),
    .X(_08746_));
 sg13g2_nor4_1 _15230_ (.A(_08737_),
    .B(_08740_),
    .C(_08743_),
    .D(_08746_),
    .Y(_08747_));
 sg13g2_nand3_1 _15231_ (.B(_08733_),
    .C(_08747_),
    .A(_08727_),
    .Y(_08748_));
 sg13g2_buf_16 clkbuf_leaf_102_clk (.X(clknet_leaf_102_clk),
    .A(clknet_8_11_0_clk));
 sg13g2_a221oi_1 _15233_ (.B2(_08723_),
    .C1(_08748_),
    .B1(_08712_),
    .A1(net10499),
    .Y(_08750_),
    .A2(_08709_));
 sg13g2_o21ai_1 _15234_ (.B1(_08750_),
    .Y(_08751_),
    .A1(_08698_),
    .A2(_08706_));
 sg13g2_inv_2 _15235_ (.Y(_08752_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[13] ));
 sg13g2_buf_16 clkbuf_leaf_106_clk (.X(clknet_leaf_106_clk),
    .A(clknet_8_61_0_clk));
 sg13g2_inv_4 _15237_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[11] ),
    .Y(_08754_));
 sg13g2_nand2b_1 _15238_ (.Y(_08755_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[10] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[10] ));
 sg13g2_o21ai_1 _15239_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[11] ),
    .Y(_08756_),
    .A1(_08754_),
    .A2(_08755_));
 sg13g2_nand2_1 _15240_ (.Y(_08757_),
    .A(_08754_),
    .B(_08755_));
 sg13g2_inv_4 _15241_ (.A(net10590),
    .Y(_08758_));
 sg13g2_nor2_1 _15242_ (.A(net10518),
    .B(_08758_),
    .Y(_08759_));
 sg13g2_a221oi_1 _15243_ (.B2(_08757_),
    .C1(_08759_),
    .B1(_08756_),
    .A1(_08752_),
    .Y(_08760_),
    .A2(net10586));
 sg13g2_inv_2 _15244_ (.Y(_08761_),
    .A(net10586));
 sg13g2_nor2b_1 _15245_ (.A(net10590),
    .B_N(net10518),
    .Y(_08762_));
 sg13g2_o21ai_1 _15246_ (.B1(_08762_),
    .Y(_08763_),
    .A1(net10517),
    .A2(_08761_));
 sg13g2_o21ai_1 _15247_ (.B1(_08763_),
    .Y(_08764_),
    .A1(_08752_),
    .A2(net10586));
 sg13g2_inv_1 _15248_ (.Y(_08765_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[15] ));
 sg13g2_and2_1 _15249_ (.A(_08765_),
    .B(_08730_),
    .X(_08766_));
 sg13g2_o21ai_1 _15250_ (.B1(_08766_),
    .Y(_08767_),
    .A1(_08760_),
    .A2(_08764_));
 sg13g2_and2_1 _15251_ (.A(net10515),
    .B(_08730_),
    .X(_08768_));
 sg13g2_o21ai_1 _15252_ (.B1(_08768_),
    .Y(_08769_),
    .A1(_08760_),
    .A2(_08764_));
 sg13g2_inv_2 _15253_ (.Y(_08770_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[15] ));
 sg13g2_a21oi_1 _15254_ (.A1(_08770_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[15] ),
    .Y(_08771_),
    .B1(_08732_));
 sg13g2_a21oi_1 _15255_ (.A1(net10515),
    .A2(_08765_),
    .Y(_08772_),
    .B1(_08771_));
 sg13g2_nand3_1 _15256_ (.B(_08769_),
    .C(_08772_),
    .A(_08767_),
    .Y(_08773_));
 sg13g2_buf_16 clkbuf_leaf_104_clk (.X(clknet_leaf_104_clk),
    .A(clknet_8_14_0_clk));
 sg13g2_nand2b_2 _15258_ (.Y(_08775_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[6] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[6] ));
 sg13g2_a21oi_1 _15259_ (.A1(_08716_),
    .A2(_08775_),
    .Y(_08776_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[7] ));
 sg13g2_o21ai_1 _15260_ (.B1(_08712_),
    .Y(_08777_),
    .A1(_08716_),
    .A2(_08775_));
 sg13g2_o21ai_1 _15261_ (.B1(net10522),
    .Y(_08778_),
    .A1(_08776_),
    .A2(_08777_));
 sg13g2_inv_4 _15262_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[9] ),
    .Y(_08779_));
 sg13g2_o21ai_1 _15263_ (.B1(_08779_),
    .Y(_08780_),
    .A1(_08776_),
    .A2(_08777_));
 sg13g2_a221oi_1 _15264_ (.B2(_08780_),
    .C1(_08748_),
    .B1(_08778_),
    .A1(_08712_),
    .Y(_08781_),
    .A2(_08723_));
 sg13g2_nor3_1 _15265_ (.A(net10499),
    .B(_08709_),
    .C(_08748_),
    .Y(_08782_));
 sg13g2_nor2_2 _15266_ (.A(_08781_),
    .B(_08782_),
    .Y(_08783_));
 sg13g2_nand3_1 _15267_ (.B(_08773_),
    .C(_08783_),
    .A(_08751_),
    .Y(_08784_));
 sg13g2_buf_16 clkbuf_leaf_105_clk (.X(clknet_leaf_105_clk),
    .A(clknet_8_62_0_clk));
 sg13g2_inv_8 _15269_ (.Y(_08786_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[18] ));
 sg13g2_nor2_1 _15270_ (.A(_08786_),
    .B(net10576),
    .Y(_08787_));
 sg13g2_nand2b_1 _15271_ (.Y(_08788_),
    .B(net10580),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[16] ));
 sg13g2_nor2_1 _15272_ (.A(_08653_),
    .B(_08788_),
    .Y(_08789_));
 sg13g2_a21oi_1 _15273_ (.A1(_08653_),
    .A2(_08788_),
    .Y(_08790_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[17] ));
 sg13g2_nor2_1 _15274_ (.A(_08789_),
    .B(_08790_),
    .Y(_08791_));
 sg13g2_nand2_1 _15275_ (.Y(_08792_),
    .A(_08786_),
    .B(net10576));
 sg13g2_o21ai_1 _15276_ (.B1(_08792_),
    .Y(_08793_),
    .A1(_08787_),
    .A2(_08791_));
 sg13g2_nand2_1 _15277_ (.Y(_08794_),
    .A(net10574),
    .B(_08793_));
 sg13g2_nor2_1 _15278_ (.A(net10574),
    .B(_08793_),
    .Y(_08795_));
 sg13g2_a21oi_1 _15279_ (.A1(net10514),
    .A2(_08794_),
    .Y(_08796_),
    .B1(_08795_));
 sg13g2_a21o_2 _15280_ (.A2(_08784_),
    .A1(_08669_),
    .B1(_08796_),
    .X(_08797_));
 sg13g2_inv_4 _15281_ (.A(net10546),
    .Y(_08798_));
 sg13g2_nor2b_2 _15282_ (.A(net10512),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[20] ),
    .Y(_08799_));
 sg13g2_nand2_1 _15283_ (.Y(_08800_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[21] ),
    .B(_08799_));
 sg13g2_inv_8 _15284_ (.Y(_08801_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[21] ));
 sg13g2_o21ai_1 _15285_ (.B1(_08801_),
    .Y(_08802_),
    .A1(net10564),
    .A2(_08799_));
 sg13g2_a21oi_1 _15286_ (.A1(_08800_),
    .A2(_08802_),
    .Y(_08803_),
    .B1(_08636_));
 sg13g2_nor3_1 _15287_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[23] ),
    .B(_08634_),
    .C(_08803_),
    .Y(_08804_));
 sg13g2_o21ai_1 _15288_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[23] ),
    .Y(_08805_),
    .A1(_08634_),
    .A2(_08803_));
 sg13g2_o21ai_1 _15289_ (.B1(_08805_),
    .Y(_08806_),
    .A1(net10511),
    .A2(_08804_));
 sg13g2_buf_16 clkbuf_leaf_111_clk (.X(clknet_leaf_111_clk),
    .A(clknet_8_15_0_clk));
 sg13g2_nor2_1 _15291_ (.A(net10553),
    .B(_08619_),
    .Y(_08808_));
 sg13g2_nand2_1 _15292_ (.Y(_08809_),
    .A(net10552),
    .B(_08619_));
 sg13g2_o21ai_1 _15293_ (.B1(_08809_),
    .Y(_08810_),
    .A1(net10510),
    .A2(_08808_));
 sg13g2_a221oi_1 _15294_ (.B2(_08607_),
    .C1(_08606_),
    .B1(_08810_),
    .A1(_08624_),
    .Y(_08811_),
    .A2(_08806_));
 sg13g2_buf_16 clkbuf_leaf_110_clk (.X(clknet_leaf_110_clk),
    .A(clknet_8_15_0_clk));
 sg13g2_o21ai_1 _15296_ (.B1(net10508),
    .Y(_08813_),
    .A1(_08798_),
    .A2(_08811_));
 sg13g2_nand2_1 _15297_ (.Y(_08814_),
    .A(_08798_),
    .B(_08811_));
 sg13g2_a22oi_1 _15298_ (.Y(_08815_),
    .B1(_08813_),
    .B2(_08814_),
    .A2(_08797_),
    .A1(_08649_));
 sg13g2_buf_16 clkbuf_leaf_108_clk (.X(clknet_leaf_108_clk),
    .A(clknet_8_14_0_clk));
 sg13g2_nor2b_2 _15300_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[28] ),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[28] ),
    .Y(_08817_));
 sg13g2_nand2_1 _15301_ (.Y(_08818_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[29] ),
    .B(_08817_));
 sg13g2_nand2_1 _15302_ (.Y(_08819_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[29] ),
    .B(_08818_));
 sg13g2_o21ai_1 _15303_ (.B1(_08819_),
    .Y(_08820_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[29] ),
    .A2(_08817_));
 sg13g2_o21ai_1 _15304_ (.B1(_08590_),
    .Y(_08821_),
    .A1(_08589_),
    .A2(_08820_));
 sg13g2_inv_1 _15305_ (.Y(_08822_),
    .A(_08821_));
 sg13g2_o21ai_1 _15306_ (.B1(_08822_),
    .Y(_08823_),
    .A1(_08601_),
    .A2(_08815_));
 sg13g2_nand2_1 _15307_ (.Y(_08824_),
    .A(_08586_),
    .B(_08823_));
 sg13g2_o21ai_1 _15308_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[31] ),
    .Y(_08825_),
    .A1(_08586_),
    .A2(_08823_));
 sg13g2_and3_1 _15309_ (.X(_08826_),
    .A(_08584_),
    .B(_08824_),
    .C(_08825_));
 sg13g2_a21oi_1 _15310_ (.A1(_08824_),
    .A2(_08825_),
    .Y(_08827_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.instr_bge ));
 sg13g2_nor2_1 _15311_ (.A(\u_ac_controller_soc_inst.u_picorv32.is_slti_blt_slt ),
    .B(\u_ac_controller_soc_inst.u_picorv32.is_sltiu_bltu_sltu ),
    .Y(_08828_));
 sg13g2_inv_1 _15312_ (.Y(_08829_),
    .A(_08748_));
 sg13g2_xor2_1 _15313_ (.B(net10522),
    .A(net10499),
    .X(_08830_));
 sg13g2_buf_16 clkbuf_leaf_119_clk (.X(clknet_leaf_119_clk),
    .A(clknet_8_24_0_clk));
 sg13g2_xor2_1 _15315_ (.B(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[1] ),
    .A(net10572),
    .X(_08832_));
 sg13g2_nand2_1 _15316_ (.Y(_08833_),
    .A(_08712_),
    .B(_08714_));
 sg13g2_xor2_1 _15317_ (.B(net10524),
    .A(net10501),
    .X(_08834_));
 sg13g2_nor4_1 _15318_ (.A(_08830_),
    .B(_08832_),
    .C(_08833_),
    .D(_08834_),
    .Y(_08835_));
 sg13g2_nor2b_2 _15319_ (.A(_08719_),
    .B_N(_08775_),
    .Y(_08836_));
 sg13g2_nor2b_2 _15320_ (.A(_08704_),
    .B_N(_08693_),
    .Y(_08837_));
 sg13g2_nand3_1 _15321_ (.B(_08836_),
    .C(_08837_),
    .A(_08835_),
    .Y(_08838_));
 sg13g2_xnor2_1 _15322_ (.Y(_08839_),
    .A(net10504),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[4] ));
 sg13g2_xnor2_1 _15323_ (.Y(_08840_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[3] ),
    .B(net10532));
 sg13g2_buf_16 clkbuf_leaf_118_clk (.X(clknet_leaf_118_clk),
    .A(clknet_8_26_0_clk));
 sg13g2_xnor2_1 _15325_ (.Y(_08842_),
    .A(net10505),
    .B(net10540));
 sg13g2_buf_16 clkbuf_leaf_117_clk (.X(clknet_leaf_117_clk),
    .A(clknet_8_24_0_clk));
 sg13g2_nor2_2 _15327_ (.A(net10599),
    .B(net10520),
    .Y(_08844_));
 sg13g2_nand2_2 _15328_ (.Y(_08845_),
    .A(net10599),
    .B(net10520));
 sg13g2_nand2b_1 _15329_ (.Y(_08846_),
    .B(_08845_),
    .A_N(_08844_));
 sg13g2_nand4_1 _15330_ (.B(_08840_),
    .C(_08842_),
    .A(_08839_),
    .Y(_08847_),
    .D(_08846_));
 sg13g2_nor3_2 _15331_ (.A(_08601_),
    .B(_08838_),
    .C(_08847_),
    .Y(_08848_));
 sg13g2_nand4_1 _15332_ (.B(_08669_),
    .C(_08829_),
    .A(_08649_),
    .Y(_08849_),
    .D(_08848_));
 sg13g2_inv_2 _15333_ (.Y(_08850_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_bgeu ));
 sg13g2_buf_2 place10911 (.A(_00006_),
    .X(net10911));
 sg13g2_a21oi_1 _15335_ (.A1(_08586_),
    .A2(_08822_),
    .Y(_08852_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[31] ));
 sg13g2_a21oi_1 _15336_ (.A1(net10533),
    .A2(_08821_),
    .Y(_08853_),
    .B1(_08852_));
 sg13g2_o21ai_1 _15337_ (.B1(_08853_),
    .Y(_08854_),
    .A1(_08601_),
    .A2(_08815_));
 sg13g2_nor2b_1 _15338_ (.A(\u_ac_controller_soc_inst.u_picorv32.is_sltiu_bltu_sltu ),
    .B_N(_08853_),
    .Y(_08855_));
 sg13g2_or2_1 _15339_ (.X(_08856_),
    .B(_08815_),
    .A(_08601_));
 sg13g2_a22oi_1 _15340_ (.Y(_08857_),
    .B1(_08855_),
    .B2(_08856_),
    .A2(_08854_),
    .A1(_08850_));
 sg13g2_a221oi_1 _15341_ (.B2(\u_ac_controller_soc_inst.u_picorv32.instr_bne ),
    .C1(_08857_),
    .B1(_08849_),
    .A1(_08303_),
    .Y(_08858_),
    .A2(_08828_));
 sg13g2_o21ai_1 _15342_ (.B1(_08858_),
    .Y(_08859_),
    .A1(_08826_),
    .A2(_08827_));
 sg13g2_buf_2 place10914 (.A(_00006_),
    .X(net10914));
 sg13g2_inv_4 _15344_ (.A(\u_ac_controller_soc_inst.u_picorv32.is_beq_bne_blt_bge_bltu_bgeu ),
    .Y(_08861_));
 sg13g2_buf_2 place9673 (.A(net9671),
    .X(net9673));
 sg13g2_and2_1 _15346_ (.A(_08303_),
    .B(_08828_),
    .X(_08863_));
 sg13g2_nand2_2 _15347_ (.Y(_08864_),
    .A(_08863_),
    .B(_08849_));
 sg13g2_inv_2 _15348_ (.Y(_08865_),
    .A(_08864_));
 sg13g2_nor4_1 _15349_ (.A(_08395_),
    .B(_08861_),
    .C(_07972_),
    .D(_08865_),
    .Y(_08866_));
 sg13g2_a22oi_1 _15350_ (.Y(_00044_),
    .B1(_08859_),
    .B2(_08866_),
    .A2(_08581_),
    .A1(_08387_));
 sg13g2_buf_2 place10908 (.A(net10906),
    .X(net10908));
 sg13g2_buf_16 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_8_55_0_clk));
 sg13g2_a21oi_1 _15353_ (.A1(_00134_),
    .A2(net10406),
    .Y(_08869_),
    .B1(_08365_));
 sg13g2_buf_2 place10913 (.A(net10912),
    .X(net10913));
 sg13g2_nor4_2 _15355_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3] ),
    .Y(_08871_),
    .D(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2] ));
 sg13g2_nand2_2 _15356_ (.Y(_08872_),
    .A(_00131_),
    .B(_08871_));
 sg13g2_buf_2 place9635 (.A(net9634),
    .X(net9635));
 sg13g2_buf_2 place10754 (.A(net10753),
    .X(net10754));
 sg13g2_buf_2 place10756 (.A(net10755),
    .X(net10756));
 sg13g2_buf_2 place9664 (.A(net9663),
    .X(net9664));
 sg13g2_buf_2 place10749 (.A(net10748),
    .X(net10749));
 sg13g2_buf_2 place9633 (.A(net9632),
    .X(net9633));
 sg13g2_mux4_1 _15363_ (.S0(net10840),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][2] ),
    .S1(net10823),
    .X(_08879_));
 sg13g2_buf_2 place10411 (.A(net10410),
    .X(net10411));
 sg13g2_mux4_1 _15365_ (.S0(net10844),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][2] ),
    .S1(net10823),
    .X(_08881_));
 sg13g2_buf_2 place10916 (.A(net10915),
    .X(net10916));
 sg13g2_buf_2 place9759 (.A(net9758),
    .X(net9759));
 sg13g2_buf_2 place9757 (.A(net9756),
    .X(net9757));
 sg13g2_mux4_1 _15369_ (.S0(net10844),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][2] ),
    .S1(net10826),
    .X(_08885_));
 sg13g2_mux4_1 _15370_ (.S0(net10842),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][2] ),
    .S1(net10824),
    .X(_08886_));
 sg13g2_buf_2 place10856 (.A(net10855),
    .X(net10856));
 sg13g2_buf_2 place10861 (.A(net10857),
    .X(net10861));
 sg13g2_buf_2 place9760 (.A(net9759),
    .X(net9760));
 sg13g2_mux4_1 _15374_ (.S0(net10780),
    .A0(_08879_),
    .A1(_08881_),
    .A2(_08885_),
    .A3(_08886_),
    .S1(net10770),
    .X(_08890_));
 sg13g2_buf_2 place9632 (.A(_10065_),
    .X(net9632));
 sg13g2_mux4_1 _15376_ (.S0(net10840),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][2] ),
    .S1(net10823),
    .X(_08892_));
 sg13g2_mux4_1 _15377_ (.S0(net10844),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][2] ),
    .S1(net10826),
    .X(_08893_));
 sg13g2_buf_2 place10740 (.A(net10739),
    .X(net10740));
 sg13g2_mux4_1 _15379_ (.S0(net10842),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][2] ),
    .S1(net10824),
    .X(_08895_));
 sg13g2_mux4_1 _15380_ (.S0(net10844),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][2] ),
    .S1(net10826),
    .X(_08896_));
 sg13g2_mux4_1 _15381_ (.S0(net10780),
    .A0(_08892_),
    .A1(_08893_),
    .A2(_08895_),
    .A3(_08896_),
    .S1(net10770),
    .X(_08897_));
 sg13g2_buf_2 place9758 (.A(net9757),
    .X(net9758));
 sg13g2_buf_2 place10829 (.A(net10827),
    .X(net10829));
 sg13g2_mux2_1 _15384_ (.A0(_08890_),
    .A1(_08897_),
    .S(net10762),
    .X(_08900_));
 sg13g2_nand2_2 _15385_ (.Y(_08901_),
    .A(_08872_),
    .B(_08900_));
 sg13g2_nand2_1 _15386_ (.Y(_08902_),
    .A(net10632),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2] ));
 sg13g2_o21ai_1 _15387_ (.B1(_08902_),
    .Y(_08903_),
    .A1(net10632),
    .A2(_08901_));
 sg13g2_nor2_1 _15388_ (.A(net10705),
    .B(_08903_),
    .Y(_08904_));
 sg13g2_a21oi_1 _15389_ (.A1(net10705),
    .A2(_08869_),
    .Y(_00048_),
    .B1(_08904_));
 sg13g2_inv_1 _15390_ (.Y(_08905_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_sh[1] ));
 sg13g2_inv_1 _15391_ (.Y(_08906_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_sh[0] ));
 sg13g2_a21oi_1 _15392_ (.A1(_08905_),
    .A2(_08906_),
    .Y(_08907_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.reg_sh[4] ));
 sg13g2_nor3_1 _15393_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_sh[2] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_sh[3] ),
    .C(_08907_),
    .Y(_08908_));
 sg13g2_a21oi_1 _15394_ (.A1(\u_ac_controller_soc_inst.u_picorv32.reg_sh[2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_sh[3] ),
    .Y(_08909_),
    .B1(_08908_));
 sg13g2_mux4_1 _15395_ (.S0(net10829),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][3] ),
    .S1(net10813),
    .X(_08910_));
 sg13g2_mux4_1 _15396_ (.S0(net10829),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][3] ),
    .S1(net10813),
    .X(_08911_));
 sg13g2_mux4_1 _15397_ (.S0(net10830),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][3] ),
    .S1(net10814),
    .X(_08912_));
 sg13g2_mux4_1 _15398_ (.S0(net10829),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][3] ),
    .S1(net10813),
    .X(_08913_));
 sg13g2_buf_2 place10828 (.A(net10827),
    .X(net10828));
 sg13g2_mux4_1 _15400_ (.S0(net10780),
    .A0(_08910_),
    .A1(_08911_),
    .A2(_08912_),
    .A3(_08913_),
    .S1(net10772),
    .X(_08915_));
 sg13g2_mux4_1 _15401_ (.S0(net10832),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][3] ),
    .S1(net10809),
    .X(_08916_));
 sg13g2_mux4_1 _15402_ (.S0(net10831),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][3] ),
    .S1(net10808),
    .X(_08917_));
 sg13g2_mux4_1 _15403_ (.S0(net10831),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][3] ),
    .S1(net10808),
    .X(_08918_));
 sg13g2_mux4_1 _15404_ (.S0(net10827),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][3] ),
    .S1(net10811),
    .X(_08919_));
 sg13g2_mux4_1 _15405_ (.S0(net10779),
    .A0(_08916_),
    .A1(_08917_),
    .A2(_08918_),
    .A3(_08919_),
    .S1(net10772),
    .X(_08920_));
 sg13g2_mux2_1 _15406_ (.A0(_08915_),
    .A1(_08920_),
    .S(net10768),
    .X(_08921_));
 sg13g2_nand2_2 _15407_ (.Y(_08922_),
    .A(_08872_),
    .B(_08921_));
 sg13g2_nand2_1 _15408_ (.Y(_08923_),
    .A(net10632),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3] ));
 sg13g2_o21ai_1 _15409_ (.B1(_08923_),
    .Y(_08924_),
    .A1(net10632),
    .A2(_08922_));
 sg13g2_nor2_1 _15410_ (.A(net10705),
    .B(_08924_),
    .Y(_08925_));
 sg13g2_a21oi_1 _15411_ (.A1(net10705),
    .A2(_08909_),
    .Y(_00049_),
    .B1(_08925_));
 sg13g2_o21ai_1 _15412_ (.B1(\u_ac_controller_soc_inst.u_picorv32.reg_sh[4] ),
    .Y(_08926_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_sh[2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_sh[3] ));
 sg13g2_nor2b_1 _15413_ (.A(_08365_),
    .B_N(_08926_),
    .Y(_08927_));
 sg13g2_mux4_1 _15414_ (.S0(net10851),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][4] ),
    .S1(net10810),
    .X(_08928_));
 sg13g2_mux4_1 _15415_ (.S0(net10851),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][4] ),
    .S1(net10810),
    .X(_08929_));
 sg13g2_mux4_1 _15416_ (.S0(net10851),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][4] ),
    .S1(net10810),
    .X(_08930_));
 sg13g2_mux4_1 _15417_ (.S0(net10851),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][4] ),
    .S1(net10810),
    .X(_08931_));
 sg13g2_mux4_1 _15418_ (.S0(net10779),
    .A0(_08928_),
    .A1(_08929_),
    .A2(_08930_),
    .A3(_08931_),
    .S1(net10772),
    .X(_08932_));
 sg13g2_mux4_1 _15419_ (.S0(net10851),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][4] ),
    .S1(net10810),
    .X(_08933_));
 sg13g2_mux4_1 _15420_ (.S0(net10851),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][4] ),
    .S1(net10810),
    .X(_08934_));
 sg13g2_mux4_1 _15421_ (.S0(net10851),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][4] ),
    .S1(net10810),
    .X(_08935_));
 sg13g2_mux4_1 _15422_ (.S0(net10851),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][4] ),
    .S1(net10810),
    .X(_08936_));
 sg13g2_mux4_1 _15423_ (.S0(net10779),
    .A0(_08933_),
    .A1(_08934_),
    .A2(_08935_),
    .A3(_08936_),
    .S1(net10772),
    .X(_08937_));
 sg13g2_mux2_1 _15424_ (.A0(_08932_),
    .A1(_08937_),
    .S(net10768),
    .X(_08938_));
 sg13g2_nand2_2 _15425_ (.Y(_08939_),
    .A(_08872_),
    .B(_08938_));
 sg13g2_nand2_1 _15426_ (.Y(_08940_),
    .A(net10632),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[4] ));
 sg13g2_o21ai_1 _15427_ (.B1(_08940_),
    .Y(_08941_),
    .A1(net10632),
    .A2(_08939_));
 sg13g2_nor2_1 _15428_ (.A(net10705),
    .B(_08941_),
    .Y(_08942_));
 sg13g2_a21oi_1 _15429_ (.A1(net10705),
    .A2(_08927_),
    .Y(_00050_),
    .B1(_08942_));
 sg13g2_buf_2 place10844 (.A(net10840),
    .X(net10844));
 sg13g2_nor2_1 _15431_ (.A(net10695),
    .B(net10708),
    .Y(_08944_));
 sg13g2_and2_1 _15432_ (.A(_00110_),
    .B(_08944_),
    .X(_08945_));
 sg13g2_buf_2 place10931 (.A(net10930),
    .X(net10931));
 sg13g2_buf_2 place10761 (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[4] ),
    .X(net10761));
 sg13g2_buf_2 place10869 (.A(_00009_),
    .X(net10869));
 sg13g2_buf_2 place10751 (.A(net10750),
    .X(net10751));
 sg13g2_buf_2 place10854 (.A(net10845),
    .X(net10854));
 sg13g2_buf_2 place10855 (.A(net10854),
    .X(net10855));
 sg13g2_buf_16 clkbuf_leaf_58_clk (.X(clknet_leaf_58_clk),
    .A(clknet_8_6_0_clk));
 sg13g2_buf_2 place10932 (.A(net10923),
    .X(net10932));
 sg13g2_buf_2 place9668 (.A(net9665),
    .X(net9668));
 sg13g2_nand2_1 _15442_ (.Y(_08955_),
    .A(net10650),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[32] ));
 sg13g2_buf_2 place9637 (.A(_10056_),
    .X(net9637));
 sg13g2_buf_2 place9634 (.A(_10065_),
    .X(net9634));
 sg13g2_buf_2 place10930 (.A(net10929),
    .X(net10930));
 sg13g2_buf_2 place10912 (.A(net10911),
    .X(net10912));
 sg13g2_a22oi_1 _15447_ (.Y(_08960_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[0] ),
    .B2(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstr ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[32] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh ));
 sg13g2_nand3_1 _15448_ (.B(_08955_),
    .C(_08960_),
    .A(net10435),
    .Y(_08961_));
 sg13g2_o21ai_1 _15449_ (.B1(_08961_),
    .Y(_08962_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[0] ),
    .A2(net10436));
 sg13g2_or2_1 _15450_ (.X(_08963_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[1] ),
    .A(net10601));
 sg13g2_buf_2 place10927 (.A(net10925),
    .X(net10927));
 sg13g2_buf_2 place10819 (.A(net10818),
    .X(net10819));
 sg13g2_o21ai_1 _15453_ (.B1(net10696),
    .Y(_08966_),
    .A1(_08415_),
    .A2(net10403));
 sg13g2_buf_2 place10764 (.A(_00004_),
    .X(net10764));
 sg13g2_inv_1 _15455_ (.Y(_08968_),
    .A(net10603));
 sg13g2_inv_2 _15456_ (.Y(_08969_),
    .A(net10568));
 sg13g2_buf_2 place10815 (.A(_00001_),
    .X(net10815));
 sg13g2_nor2_2 _15458_ (.A(net10601),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[1] ),
    .Y(_08971_));
 sg13g2_buf_16 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_8_8_0_clk));
 sg13g2_nor2_1 _15460_ (.A(_08969_),
    .B(_08971_),
    .Y(_08973_));
 sg13g2_nor2_1 _15461_ (.A(net10568),
    .B(_08415_),
    .Y(_08974_));
 sg13g2_a21oi_1 _15462_ (.A1(_08495_),
    .A2(_08973_),
    .Y(_08975_),
    .B1(_08974_));
 sg13g2_nand2_1 _15463_ (.Y(_08976_),
    .A(\u_ac_controller_soc_inst.io_rdata[8] ),
    .B(net10184));
 sg13g2_nand2_1 _15464_ (.Y(_08977_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[8] ),
    .B(_08425_));
 sg13g2_a22oi_1 _15465_ (.Y(_08978_),
    .B1(net10242),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[8] ),
    .A2(net10231),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[8] ));
 sg13g2_nand3_1 _15466_ (.B(_08977_),
    .C(_08978_),
    .A(_08976_),
    .Y(_08979_));
 sg13g2_mux2_1 _15467_ (.A0(_08553_),
    .A1(_08979_),
    .S(net10400),
    .X(_08980_));
 sg13g2_buf_2 place10813 (.A(net10811),
    .X(net10813));
 sg13g2_buf_2 place10817 (.A(net10816),
    .X(net10817));
 sg13g2_mux2_1 _15470_ (.A0(_08975_),
    .A1(_08980_),
    .S(net10597),
    .X(_08983_));
 sg13g2_buf_2 place10812 (.A(net10811),
    .X(net10812));
 sg13g2_nand2_1 _15472_ (.Y(_08985_),
    .A(_00052_),
    .B(net10403));
 sg13g2_a22oi_1 _15473_ (.Y(_08986_),
    .B1(_08985_),
    .B2(_08975_),
    .A2(_08983_),
    .A1(_08968_));
 sg13g2_inv_1 _15474_ (.Y(_08987_),
    .A(_00054_));
 sg13g2_a22oi_1 _15475_ (.Y(_08988_),
    .B1(_08987_),
    .B2(net10711),
    .A2(net10699),
    .A1(net10597));
 sg13g2_o21ai_1 _15476_ (.B1(_08988_),
    .Y(_08989_),
    .A1(_08966_),
    .A2(_08986_));
 sg13g2_nor2_1 _15477_ (.A(_08989_),
    .B(_08945_),
    .Y(_08990_));
 sg13g2_a21oi_1 _15478_ (.A1(_08945_),
    .A2(_08962_),
    .Y(_02144_),
    .B1(_08990_));
 sg13g2_buf_2 place10915 (.A(_00006_),
    .X(net10915));
 sg13g2_nand2_1 _15480_ (.Y(_08992_),
    .A(net10650),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[33] ));
 sg13g2_buf_2 place10919 (.A(_00006_),
    .X(net10919));
 sg13g2_a22oi_1 _15482_ (.Y(_08994_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[1] ),
    .B2(net10645),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[33] ),
    .A1(net10641));
 sg13g2_nand3_1 _15483_ (.B(_08992_),
    .C(_08994_),
    .A(net10434),
    .Y(_08995_));
 sg13g2_o21ai_1 _15484_ (.B1(_08995_),
    .Y(_08996_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[1] ),
    .A2(net10436));
 sg13g2_nand2_2 _15485_ (.Y(_08997_),
    .A(_00110_),
    .B(_08944_));
 sg13g2_buf_2 place10840 (.A(net10833),
    .X(net10840));
 sg13g2_buf_16 clkbuf_leaf_86_clk (.X(clknet_leaf_86_clk),
    .A(clknet_8_9_0_clk));
 sg13g2_buf_16 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_8_4_0_clk));
 sg13g2_buf_16 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_8_6_0_clk));
 sg13g2_xor2_1 _15490_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[1] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[1] ),
    .X(_09002_));
 sg13g2_buf_2 place10843 (.A(net10842),
    .X(net10843));
 sg13g2_a22oi_1 _15492_ (.Y(_09004_),
    .B1(_09002_),
    .B2(net10711),
    .A2(net10699),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[1] ));
 sg13g2_buf_2 place10810 (.A(net10808),
    .X(net10810));
 sg13g2_o21ai_1 _15494_ (.B1(_00052_),
    .Y(_09006_),
    .A1(net10595),
    .A2(_00129_));
 sg13g2_inv_1 _15495_ (.Y(_09007_),
    .A(_09006_));
 sg13g2_nor2_1 _15496_ (.A(net10400),
    .B(_09007_),
    .Y(_09008_));
 sg13g2_nor2b_2 _15497_ (.A(_00129_),
    .B_N(net10595),
    .Y(_09009_));
 sg13g2_inv_2 _15498_ (.Y(_09010_),
    .A(\u_ac_controller_soc_inst.io_rdata[25] ));
 sg13g2_a22oi_1 _15499_ (.Y(_09011_),
    .B1(net10243),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[25] ),
    .A2(net10230),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[25] ));
 sg13g2_o21ai_1 _15500_ (.B1(_09011_),
    .Y(_09012_),
    .A1(_09010_),
    .A2(net10186));
 sg13g2_buf_16 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_8_5_0_clk));
 sg13g2_inv_1 _15502_ (.Y(_09014_),
    .A(\u_ac_controller_soc_inst.io_rdata[9] ));
 sg13g2_a22oi_1 _15503_ (.Y(_09015_),
    .B1(net10242),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[9] ),
    .A2(net10231),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[9] ));
 sg13g2_o21ai_1 _15504_ (.B1(_09015_),
    .Y(_09016_),
    .A1(_09014_),
    .A2(net10186));
 sg13g2_mux2_1 _15505_ (.A0(_09012_),
    .A1(_09016_),
    .S(net10400),
    .X(_09017_));
 sg13g2_a22oi_1 _15506_ (.Y(_09018_),
    .B1(_09009_),
    .B2(_09017_),
    .A2(_09008_),
    .A1(_08506_));
 sg13g2_o21ai_1 _15507_ (.B1(net10403),
    .Y(_09019_),
    .A1(net10568),
    .A2(_09007_));
 sg13g2_nand2_1 _15508_ (.Y(_09020_),
    .A(_08428_),
    .B(_09019_));
 sg13g2_o21ai_1 _15509_ (.B1(_09020_),
    .Y(_09021_),
    .A1(_08971_),
    .A2(_09018_));
 sg13g2_nand2_1 _15510_ (.Y(_09022_),
    .A(net10696),
    .B(_09021_));
 sg13g2_and3_1 _15511_ (.X(_09023_),
    .A(net10281),
    .B(_09004_),
    .C(_09022_));
 sg13g2_a21oi_2 _15512_ (.B1(_09023_),
    .Y(_02155_),
    .A2(_08996_),
    .A1(net10285));
 sg13g2_buf_16 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_8_4_0_clk));
 sg13g2_buf_2 place10807 (.A(net10805),
    .X(net10807));
 sg13g2_nand2_1 _15515_ (.Y(_09026_),
    .A(net10651),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[34] ));
 sg13g2_buf_2 place10806 (.A(net10805),
    .X(net10806));
 sg13g2_buf_16 clkbuf_leaf_101_clk (.X(clknet_leaf_101_clk),
    .A(clknet_8_10_0_clk));
 sg13g2_a22oi_1 _15518_ (.Y(_09029_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[2] ),
    .B2(net10645),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[34] ),
    .A1(net10641));
 sg13g2_nand3_1 _15519_ (.B(_09026_),
    .C(_09029_),
    .A(net10437),
    .Y(_09030_));
 sg13g2_o21ai_1 _15520_ (.B1(_09030_),
    .Y(_09031_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[2] ),
    .A2(net10436));
 sg13g2_buf_2 place10929 (.A(net10924),
    .X(net10929));
 sg13g2_buf_16 clkbuf_leaf_85_clk (.X(clknet_leaf_85_clk),
    .A(clknet_8_9_0_clk));
 sg13g2_nand2_1 _15523_ (.Y(_09034_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[1] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[1] ));
 sg13g2_buf_16 clkbuf_leaf_88_clk (.X(clknet_leaf_88_clk),
    .A(clknet_8_10_0_clk));
 sg13g2_buf_16 clkbuf_leaf_69_clk (.X(clknet_leaf_69_clk),
    .A(clknet_8_18_0_clk));
 sg13g2_buf_2 place10835 (.A(net10834),
    .X(net10835));
 sg13g2_xor2_1 _15527_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[2] ),
    .A(net10491),
    .X(_09038_));
 sg13g2_xnor2_1 _15528_ (.Y(_09039_),
    .A(_09034_),
    .B(_09038_));
 sg13g2_a22oi_1 _15529_ (.Y(_09040_),
    .B1(_09039_),
    .B2(net10711),
    .A2(net10540),
    .A1(net10699));
 sg13g2_and2_1 _15530_ (.A(\u_ac_controller_soc_inst.spi_sensor_rdata[26] ),
    .B(net10243),
    .X(_09041_));
 sg13g2_a221oi_1 _15531_ (.B2(\u_ac_controller_soc_inst.io_rdata[26] ),
    .C1(_09041_),
    .B1(_08420_),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[26] ),
    .Y(_09042_),
    .A2(net10232));
 sg13g2_buf_2 place10830 (.A(net10829),
    .X(net10830));
 sg13g2_mux2_1 _15533_ (.A0(_08510_),
    .A1(_09042_),
    .S(net10596),
    .X(_09044_));
 sg13g2_and2_1 _15534_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[10] ),
    .B(net10231),
    .X(_09045_));
 sg13g2_a221oi_1 _15535_ (.B2(\u_ac_controller_soc_inst.io_rdata[10] ),
    .C1(_09045_),
    .B1(net10184),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[10] ),
    .Y(_09046_),
    .A2(net10242));
 sg13g2_buf_2 place10832 (.A(net10831),
    .X(net10832));
 sg13g2_nor2b_2 _15537_ (.A(net10571),
    .B_N(net10596),
    .Y(_09048_));
 sg13g2_buf_2 place10831 (.A(net10827),
    .X(net10831));
 sg13g2_a221oi_1 _15539_ (.B2(_09048_),
    .C1(net10603),
    .B1(_09046_),
    .A1(net10570),
    .Y(_09050_),
    .A2(_09044_));
 sg13g2_a21oi_1 _15540_ (.A1(net10597),
    .A2(_09050_),
    .Y(_09051_),
    .B1(net10569));
 sg13g2_o21ai_1 _15541_ (.B1(_08434_),
    .Y(_09052_),
    .A1(net10396),
    .A2(_09051_));
 sg13g2_buf_2 place10839 (.A(net10835),
    .X(net10839));
 sg13g2_a21oi_1 _15543_ (.A1(net10569),
    .A2(_08510_),
    .Y(_09054_),
    .B1(_00052_));
 sg13g2_or3_1 _15544_ (.A(net10396),
    .B(_09050_),
    .C(_09054_),
    .X(_09055_));
 sg13g2_nand3_1 _15545_ (.B(_09052_),
    .C(_09055_),
    .A(net10696),
    .Y(_09056_));
 sg13g2_and3_1 _15546_ (.X(_09057_),
    .A(net10281),
    .B(_09040_),
    .C(_09056_));
 sg13g2_a21oi_2 _15547_ (.B1(_09057_),
    .Y(_02166_),
    .A2(_09031_),
    .A1(net10285));
 sg13g2_buf_2 place10838 (.A(net10835),
    .X(net10838));
 sg13g2_nand2_1 _15549_ (.Y(_09059_),
    .A(net10651),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[35] ));
 sg13g2_buf_2 place10842 (.A(net10840),
    .X(net10842));
 sg13g2_a22oi_1 _15551_ (.Y(_09061_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[3] ),
    .B2(net10645),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[35] ),
    .A1(net10641));
 sg13g2_nand3_1 _15552_ (.B(_09059_),
    .C(_09061_),
    .A(net10437),
    .Y(_09062_));
 sg13g2_o21ai_1 _15553_ (.B1(_09062_),
    .Y(_09063_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[3] ),
    .A2(net10436));
 sg13g2_nor2_2 _15554_ (.A(net10491),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[2] ),
    .Y(_09064_));
 sg13g2_a22oi_1 _15555_ (.Y(_09065_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[2] ),
    .B2(net10491),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[1] ));
 sg13g2_buf_2 place10837 (.A(net10836),
    .X(net10837));
 sg13g2_nor2_2 _15557_ (.A(_09064_),
    .B(_09065_),
    .Y(_09067_));
 sg13g2_buf_2 place10918 (.A(net10915),
    .X(net10918));
 sg13g2_buf_16 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_8_4_0_clk));
 sg13g2_xnor2_1 _15560_ (.Y(_09070_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[3] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[3] ));
 sg13g2_xnor2_1 _15561_ (.Y(_09071_),
    .A(_09067_),
    .B(_09070_));
 sg13g2_a22oi_1 _15562_ (.Y(_09072_),
    .B1(_09071_),
    .B2(net10711),
    .A2(net10532),
    .A1(net10699));
 sg13g2_and2_1 _15563_ (.A(\u_ac_controller_soc_inst.spi_sensor_rdata[27] ),
    .B(net10245),
    .X(_09073_));
 sg13g2_a221oi_1 _15564_ (.B2(\u_ac_controller_soc_inst.io_rdata[27] ),
    .C1(_09073_),
    .B1(net10185),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[27] ),
    .Y(_09074_),
    .A2(net10233));
 sg13g2_buf_16 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_8_0_0_clk));
 sg13g2_mux2_1 _15566_ (.A0(_08515_),
    .A1(_09074_),
    .S(net10596),
    .X(_09076_));
 sg13g2_and2_1 _15567_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[11] ),
    .B(net10232),
    .X(_09077_));
 sg13g2_a221oi_1 _15568_ (.B2(\u_ac_controller_soc_inst.io_rdata[11] ),
    .C1(_09077_),
    .B1(net10183),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[11] ),
    .Y(_09078_),
    .A2(net10242));
 sg13g2_buf_2 place10841 (.A(net10840),
    .X(net10841));
 sg13g2_a221oi_1 _15570_ (.B2(_09048_),
    .C1(net10603),
    .B1(_09078_),
    .A1(net10570),
    .Y(_09080_),
    .A2(_09076_));
 sg13g2_a21oi_1 _15571_ (.A1(net10597),
    .A2(_09080_),
    .Y(_09081_),
    .B1(net10569));
 sg13g2_o21ai_1 _15572_ (.B1(_08439_),
    .Y(_09082_),
    .A1(net10396),
    .A2(_09081_));
 sg13g2_a21oi_1 _15573_ (.A1(net10569),
    .A2(_08515_),
    .Y(_09083_),
    .B1(_00052_));
 sg13g2_or3_1 _15574_ (.A(net10396),
    .B(_09080_),
    .C(_09083_),
    .X(_09084_));
 sg13g2_nand3_1 _15575_ (.B(_09082_),
    .C(_09084_),
    .A(net10696),
    .Y(_09085_));
 sg13g2_and3_1 _15576_ (.X(_09086_),
    .A(net10281),
    .B(_09072_),
    .C(_09085_));
 sg13g2_a21oi_2 _15577_ (.B1(_09086_),
    .Y(_02169_),
    .A2(_09063_),
    .A1(net10285));
 sg13g2_buf_2 place10834 (.A(net10833),
    .X(net10834));
 sg13g2_buf_16 clkbuf_leaf_96_clk (.X(clknet_leaf_96_clk),
    .A(clknet_8_59_0_clk));
 sg13g2_buf_16 clkbuf_leaf_75_clk (.X(clknet_leaf_75_clk),
    .A(clknet_8_12_0_clk));
 sg13g2_nor2_1 _15581_ (.A(net10490),
    .B(net10673),
    .Y(_09090_));
 sg13g2_inv_1 _15582_ (.Y(_09091_),
    .A(_09090_));
 sg13g2_nand2_1 _15583_ (.Y(_09092_),
    .A(net10490),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[3] ));
 sg13g2_o21ai_1 _15584_ (.B1(_09092_),
    .Y(_09093_),
    .A1(_09064_),
    .A2(_09065_));
 sg13g2_and2_1 _15585_ (.A(_09091_),
    .B(_09093_),
    .X(_09094_));
 sg13g2_buf_2 place10836 (.A(net10835),
    .X(net10836));
 sg13g2_buf_16 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_8_4_0_clk));
 sg13g2_buf_2 place10833 (.A(_00000_),
    .X(net10833));
 sg13g2_xnor2_1 _15589_ (.Y(_09098_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[4] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[4] ));
 sg13g2_xnor2_1 _15590_ (.Y(_09099_),
    .A(_09094_),
    .B(_09098_));
 sg13g2_buf_16 clkbuf_leaf_68_clk (.X(clknet_leaf_68_clk),
    .A(clknet_8_13_0_clk));
 sg13g2_a21oi_1 _15592_ (.A1(_08470_),
    .A2(_09048_),
    .Y(_09101_),
    .B1(net10603));
 sg13g2_a21o_1 _15593_ (.A2(_09101_),
    .A1(net10598),
    .B1(net10570),
    .X(_09102_));
 sg13g2_a21oi_1 _15594_ (.A1(net10403),
    .A2(_09102_),
    .Y(_09103_),
    .B1(_08448_));
 sg13g2_nand2_1 _15595_ (.Y(_09104_),
    .A(_08520_),
    .B(_08521_));
 sg13g2_and2_1 _15596_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[28] ),
    .B(net10232),
    .X(_09105_));
 sg13g2_a221oi_1 _15597_ (.B2(\u_ac_controller_soc_inst.io_rdata[28] ),
    .C1(_09105_),
    .B1(net10185),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[28] ),
    .Y(_09106_),
    .A2(net10244));
 sg13g2_buf_2 place10909 (.A(net10905),
    .X(net10909));
 sg13g2_nand2_1 _15599_ (.Y(_09108_),
    .A(net10598),
    .B(_09106_));
 sg13g2_o21ai_1 _15600_ (.B1(_09108_),
    .Y(_09109_),
    .A1(net10598),
    .A2(_09104_));
 sg13g2_inv_1 _15601_ (.Y(_09110_),
    .A(_09101_));
 sg13g2_a21oi_1 _15602_ (.A1(net10570),
    .A2(_09109_),
    .Y(_09111_),
    .B1(_09110_));
 sg13g2_a21oi_1 _15603_ (.A1(net10569),
    .A2(_08522_),
    .Y(_09112_),
    .B1(_00052_));
 sg13g2_nor3_1 _15604_ (.A(net10396),
    .B(_09111_),
    .C(_09112_),
    .Y(_09113_));
 sg13g2_nor3_2 _15605_ (.A(net10460),
    .B(_09103_),
    .C(_09113_),
    .Y(_09114_));
 sg13g2_a221oi_1 _15606_ (.B2(net10711),
    .C1(_09114_),
    .B1(_09099_),
    .A1(net10699),
    .Y(_09115_),
    .A2(net10530));
 sg13g2_buf_2 place10910 (.A(net10905),
    .X(net10910));
 sg13g2_nor3_2 _15608_ (.A(net10639),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstr ),
    .C(net10647),
    .Y(_09117_));
 sg13g2_buf_16 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_8_2_0_clk));
 sg13g2_nand2b_1 _15610_ (.Y(_09119_),
    .B(net10395),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.count_cycle[4] ));
 sg13g2_buf_16 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_8_3_0_clk));
 sg13g2_buf_16 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_8_53_0_clk));
 sg13g2_buf_16 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_8_54_0_clk));
 sg13g2_buf_16 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_8_54_0_clk));
 sg13g2_nand2_1 _15615_ (.Y(_09124_),
    .A(net10651),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[36] ));
 sg13g2_buf_16 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_8_54_0_clk));
 sg13g2_buf_16 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_8_0_0_clk));
 sg13g2_buf_16 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_8_2_0_clk));
 sg13g2_buf_2 place10824 (.A(net10823),
    .X(net10824));
 sg13g2_a22oi_1 _15620_ (.Y(_09129_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[4] ),
    .B2(net10645),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[36] ),
    .A1(net10641));
 sg13g2_nand3_1 _15621_ (.B(_09124_),
    .C(_09129_),
    .A(net10437),
    .Y(_09130_));
 sg13g2_a21oi_2 _15622_ (.B1(net10282),
    .Y(_09131_),
    .A2(_09130_),
    .A1(_09119_));
 sg13g2_a21oi_2 _15623_ (.B1(_09131_),
    .Y(_02170_),
    .A2(_09115_),
    .A1(net10281));
 sg13g2_buf_2 place10825 (.A(net10824),
    .X(net10825));
 sg13g2_or2_1 _15625_ (.X(_09133_),
    .B(net10672),
    .A(net10489));
 sg13g2_and2_1 _15626_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[4] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[4] ),
    .X(_09134_));
 sg13g2_a21o_1 _15627_ (.A2(_09133_),
    .A1(_09094_),
    .B1(_09134_),
    .X(_09135_));
 sg13g2_buf_16 clkbuf_leaf_84_clk (.X(clknet_leaf_84_clk),
    .A(clknet_8_9_0_clk));
 sg13g2_buf_2 place10933 (.A(net10932),
    .X(net10933));
 sg13g2_buf_2 place10818 (.A(net10817),
    .X(net10818));
 sg13g2_xnor2_1 _15631_ (.Y(_09139_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[5] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[5] ));
 sg13g2_xnor2_1 _15632_ (.Y(_09140_),
    .A(_09135_),
    .B(_09139_));
 sg13g2_a21oi_1 _15633_ (.A1(_08464_),
    .A2(_09048_),
    .Y(_09141_),
    .B1(net10603));
 sg13g2_a21o_1 _15634_ (.A2(_09141_),
    .A1(net10598),
    .B1(net10570),
    .X(_09142_));
 sg13g2_a21oi_1 _15635_ (.A1(net10403),
    .A2(_09142_),
    .Y(_09143_),
    .B1(_08454_));
 sg13g2_nand2_1 _15636_ (.Y(_09144_),
    .A(_08529_),
    .B(_08530_));
 sg13g2_buf_2 place11032 (.A(net11003),
    .X(net11032));
 sg13g2_and2_1 _15638_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[29] ),
    .B(net10230),
    .X(_09146_));
 sg13g2_a221oi_1 _15639_ (.B2(\u_ac_controller_soc_inst.io_rdata[29] ),
    .C1(_09146_),
    .B1(net10183),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[29] ),
    .Y(_09147_),
    .A2(_07887_));
 sg13g2_nand2_1 _15640_ (.Y(_09148_),
    .A(net10598),
    .B(_09147_));
 sg13g2_o21ai_1 _15641_ (.B1(_09148_),
    .Y(_09149_),
    .A1(net10598),
    .A2(_09144_));
 sg13g2_inv_1 _15642_ (.Y(_09150_),
    .A(_09141_));
 sg13g2_a21oi_1 _15643_ (.A1(net10570),
    .A2(_09149_),
    .Y(_09151_),
    .B1(_09150_));
 sg13g2_a21oi_1 _15644_ (.A1(net10569),
    .A2(_08531_),
    .Y(_09152_),
    .B1(_00052_));
 sg13g2_nor3_1 _15645_ (.A(net10396),
    .B(_09151_),
    .C(_09152_),
    .Y(_09153_));
 sg13g2_nor3_2 _15646_ (.A(net10460),
    .B(_09143_),
    .C(_09153_),
    .Y(_09154_));
 sg13g2_a221oi_1 _15647_ (.B2(net10711),
    .C1(_09154_),
    .B1(_09140_),
    .A1(net10699),
    .Y(_09155_),
    .A2(net10529));
 sg13g2_buf_2 place11020 (.A(net11018),
    .X(net11020));
 sg13g2_nand2b_1 _15649_ (.Y(_09157_),
    .B(net10395),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.count_cycle[5] ));
 sg13g2_nand2_1 _15650_ (.Y(_09158_),
    .A(net10651),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[37] ));
 sg13g2_buf_2 place11024 (.A(net11023),
    .X(net11024));
 sg13g2_a22oi_1 _15652_ (.Y(_09160_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[5] ),
    .B2(net10646),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[37] ),
    .A1(net10642));
 sg13g2_nand3_1 _15653_ (.B(_09158_),
    .C(_09160_),
    .A(net10437),
    .Y(_09161_));
 sg13g2_a21oi_2 _15654_ (.B1(net10282),
    .Y(_09162_),
    .A2(_09161_),
    .A1(_09157_));
 sg13g2_a21oi_2 _15655_ (.B1(_09162_),
    .Y(_02171_),
    .A2(_09155_),
    .A1(net10281));
 sg13g2_buf_2 place10821 (.A(net10817),
    .X(net10821));
 sg13g2_a221oi_1 _15657_ (.B2(_09093_),
    .C1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[5] ),
    .B1(_09091_),
    .A1(net10489),
    .Y(_09164_),
    .A2(net10672));
 sg13g2_buf_2 place10820 (.A(net10818),
    .X(net10820));
 sg13g2_o21ai_1 _15659_ (.B1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[5] ),
    .Y(_09166_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[5] ),
    .A2(_09133_));
 sg13g2_or2_1 _15660_ (.X(_09167_),
    .B(_09166_),
    .A(_09164_));
 sg13g2_nand2_1 _15661_ (.Y(_09168_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[5] ),
    .B(_09135_));
 sg13g2_nand2_1 _15662_ (.Y(_09169_),
    .A(_09167_),
    .B(_09168_));
 sg13g2_buf_16 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_8_1_0_clk));
 sg13g2_buf_16 clkbuf_leaf_81_clk (.X(clknet_leaf_81_clk),
    .A(clknet_8_13_0_clk));
 sg13g2_xnor2_1 _15665_ (.Y(_09172_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[6] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[6] ));
 sg13g2_xnor2_1 _15666_ (.Y(_09173_),
    .A(_09169_),
    .B(_09172_));
 sg13g2_a21oi_1 _15667_ (.A1(_08476_),
    .A2(_09048_),
    .Y(_09174_),
    .B1(net10603));
 sg13g2_a21o_1 _15668_ (.A2(_09174_),
    .A1(net10598),
    .B1(net10570),
    .X(_09175_));
 sg13g2_a21oi_1 _15669_ (.A1(net10403),
    .A2(_09175_),
    .Y(_09176_),
    .B1(_08459_));
 sg13g2_and2_1 _15670_ (.A(\u_ac_controller_soc_inst.spi_flash_rdata[30] ),
    .B(net10232),
    .X(_09177_));
 sg13g2_a221oi_1 _15671_ (.B2(\u_ac_controller_soc_inst.io_rdata[30] ),
    .C1(_09177_),
    .B1(net10185),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[30] ),
    .Y(_09178_),
    .A2(net10244));
 sg13g2_buf_2 place11053 (.A(net11052),
    .X(net11053));
 sg13g2_mux2_1 _15673_ (.A0(_08537_),
    .A1(_09178_),
    .S(net10598),
    .X(_09180_));
 sg13g2_inv_1 _15674_ (.Y(_09181_),
    .A(_09174_));
 sg13g2_a21oi_1 _15675_ (.A1(net10570),
    .A2(_09180_),
    .Y(_09182_),
    .B1(_09181_));
 sg13g2_a21oi_1 _15676_ (.A1(net10569),
    .A2(_08537_),
    .Y(_09183_),
    .B1(_00052_));
 sg13g2_nor3_1 _15677_ (.A(net10396),
    .B(_09182_),
    .C(_09183_),
    .Y(_09184_));
 sg13g2_nor3_2 _15678_ (.A(net10460),
    .B(_09176_),
    .C(_09184_),
    .Y(_09185_));
 sg13g2_a221oi_1 _15679_ (.B2(net10711),
    .C1(_09185_),
    .B1(_09173_),
    .A1(net10699),
    .Y(_09186_),
    .A2(net10527));
 sg13g2_buf_16 clkbuf_leaf_60_clk (.X(clknet_leaf_60_clk),
    .A(clknet_8_3_0_clk));
 sg13g2_nand2b_1 _15681_ (.Y(_09188_),
    .B(net10395),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.count_cycle[6] ));
 sg13g2_nand2_1 _15682_ (.Y(_09189_),
    .A(net10651),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[38] ));
 sg13g2_buf_16 clkbuf_leaf_77_clk (.X(clknet_leaf_77_clk),
    .A(clknet_8_11_0_clk));
 sg13g2_a22oi_1 _15684_ (.Y(_09191_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[6] ),
    .B2(net10646),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[38] ),
    .A1(net10642));
 sg13g2_nand3_1 _15685_ (.B(_09189_),
    .C(_09191_),
    .A(net10437),
    .Y(_09192_));
 sg13g2_a21oi_2 _15686_ (.B1(net10282),
    .Y(_09193_),
    .A2(_09192_),
    .A1(_09188_));
 sg13g2_a21oi_1 _15687_ (.A1(net10281),
    .A2(_09186_),
    .Y(_02172_),
    .B1(_09193_));
 sg13g2_buf_2 place10934 (.A(net10932),
    .X(net10934));
 sg13g2_buf_2 place11030 (.A(net11029),
    .X(net11030));
 sg13g2_nand2_1 _15690_ (.Y(_09196_),
    .A(net10651),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[39] ));
 sg13g2_buf_2 place11017 (.A(net11016),
    .X(net11017));
 sg13g2_buf_2 place11028 (.A(net11027),
    .X(net11028));
 sg13g2_a22oi_1 _15693_ (.Y(_09199_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[7] ),
    .B2(net10646),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[39] ),
    .A1(net10642));
 sg13g2_nand3_1 _15694_ (.B(_09196_),
    .C(_09199_),
    .A(net10435),
    .Y(_09200_));
 sg13g2_o21ai_1 _15695_ (.B1(_09200_),
    .Y(_09201_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[7] ),
    .A2(net10437));
 sg13g2_nand3_1 _15696_ (.B(_08483_),
    .C(_09009_),
    .A(_08969_),
    .Y(_09202_));
 sg13g2_nor2_1 _15697_ (.A(_08543_),
    .B(_09007_),
    .Y(_09203_));
 sg13g2_nand2b_1 _15698_ (.Y(_09204_),
    .B(\u_ac_controller_soc_inst.io_rdata[31] ),
    .A_N(net10245));
 sg13g2_inv_1 _15699_ (.Y(_09205_),
    .A(_00127_));
 sg13g2_inv_1 _15700_ (.Y(_09206_),
    .A(_00128_));
 sg13g2_a22oi_1 _15701_ (.Y(_09207_),
    .B1(net10244),
    .B2(_09206_),
    .A2(net10231),
    .A1(_09205_));
 sg13g2_o21ai_1 _15702_ (.B1(_09207_),
    .Y(_09208_),
    .A1(_08408_),
    .A2(_09204_));
 sg13g2_buf_2 place11052 (.A(net11051),
    .X(net11052));
 sg13g2_and2_1 _15704_ (.A(_09009_),
    .B(_09208_),
    .X(_09210_));
 sg13g2_o21ai_1 _15705_ (.B1(net10568),
    .Y(_09211_),
    .A1(_09203_),
    .A2(_09210_));
 sg13g2_a21oi_1 _15706_ (.A1(_09202_),
    .A2(_09211_),
    .Y(_09212_),
    .B1(_08971_));
 sg13g2_buf_2 place10996 (.A(net10993),
    .X(net10996));
 sg13g2_a22oi_1 _15708_ (.Y(_09214_),
    .B1(_07927_),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[7] ),
    .A2(net10247),
    .A1(\u_ac_controller_soc_inst.io_rdata[7] ));
 sg13g2_inv_1 _15709_ (.Y(_09215_),
    .A(_00126_));
 sg13g2_a22oi_1 _15710_ (.Y(_09216_),
    .B1(net10243),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[7] ),
    .A2(net10230),
    .A1(_09215_));
 sg13g2_o21ai_1 _15711_ (.B1(_09216_),
    .Y(_09217_),
    .A1(_00086_),
    .A2(_09214_));
 sg13g2_and2_1 _15712_ (.A(_09019_),
    .B(_09217_),
    .X(_09218_));
 sg13g2_nor2_1 _15713_ (.A(_09212_),
    .B(_09218_),
    .Y(_09219_));
 sg13g2_buf_2 place11040 (.A(net11039),
    .X(net11040));
 sg13g2_buf_16 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_8_5_0_clk));
 sg13g2_buf_2 place11051 (.A(net11050),
    .X(net11051));
 sg13g2_xor2_1 _15717_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[7] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[7] ),
    .X(_09223_));
 sg13g2_nor2_1 _15718_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[6] ),
    .B(net10670),
    .Y(_09224_));
 sg13g2_a21oi_1 _15719_ (.A1(_09167_),
    .A2(_09168_),
    .Y(_09225_),
    .B1(_09224_));
 sg13g2_a21oi_1 _15720_ (.A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[6] ),
    .Y(_09226_),
    .B1(_09225_));
 sg13g2_xnor2_1 _15721_ (.Y(_09227_),
    .A(_09223_),
    .B(_09226_));
 sg13g2_a22oi_1 _15722_ (.Y(_09228_),
    .B1(_09227_),
    .B2(net10712),
    .A2(net10524),
    .A1(net10700));
 sg13g2_o21ai_1 _15723_ (.B1(_09228_),
    .Y(_09229_),
    .A1(net10460),
    .A2(_09219_));
 sg13g2_nor2_1 _15724_ (.A(net10285),
    .B(_09229_),
    .Y(_09230_));
 sg13g2_a21oi_2 _15725_ (.B1(_09230_),
    .Y(_02173_),
    .A2(_09201_),
    .A1(net10285));
 sg13g2_buf_2 place10983 (.A(net10982),
    .X(net10983));
 sg13g2_nand2_1 _15727_ (.Y(_09232_),
    .A(net10651),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[40] ));
 sg13g2_buf_2 place10982 (.A(net10981),
    .X(net10982));
 sg13g2_a22oi_1 _15729_ (.Y(_09234_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[8] ),
    .B2(net10646),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[40] ),
    .A1(net10642));
 sg13g2_nand3_1 _15730_ (.B(_09232_),
    .C(_09234_),
    .A(net10435),
    .Y(_09235_));
 sg13g2_o21ai_1 _15731_ (.B1(_09235_),
    .Y(_09236_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[8] ),
    .A2(net10436));
 sg13g2_buf_2 place10920 (.A(net10919),
    .X(net10920));
 sg13g2_nor2_1 _15733_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[7] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[7] ),
    .Y(_09238_));
 sg13g2_nand2_2 _15734_ (.Y(_09239_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[7] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[7] ));
 sg13g2_o21ai_1 _15735_ (.B1(_09239_),
    .Y(_09240_),
    .A1(_09226_),
    .A2(_09238_));
 sg13g2_buf_2 place10922 (.A(net10921),
    .X(net10922));
 sg13g2_buf_2 place10975 (.A(net10974),
    .X(net10975));
 sg13g2_xnor2_1 _15738_ (.Y(_09243_),
    .A(net10488),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[8] ));
 sg13g2_xnor2_1 _15739_ (.Y(_09244_),
    .A(_09240_),
    .B(_09243_));
 sg13g2_a22oi_1 _15740_ (.Y(_09245_),
    .B1(_09244_),
    .B2(net10712),
    .A2(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[8] ),
    .A1(net10700));
 sg13g2_buf_2 place10993 (.A(net10990),
    .X(net10993));
 sg13g2_nor2b_2 _15742_ (.A(_09219_),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.latched_is_lb ),
    .Y(_09247_));
 sg13g2_buf_2 place10997 (.A(net10996),
    .X(net10997));
 sg13g2_buf_2 place10947 (.A(net10935),
    .X(net10947));
 sg13g2_nor2b_2 _15745_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_is_lh ),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.latched_is_lb ),
    .Y(_09250_));
 sg13g2_a22oi_1 _15746_ (.Y(_09251_),
    .B1(_08980_),
    .B2(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[2] ),
    .A2(_08979_),
    .A1(net10399));
 sg13g2_nor2_1 _15747_ (.A(_09250_),
    .B(_09251_),
    .Y(_09252_));
 sg13g2_o21ai_1 _15748_ (.B1(net10696),
    .Y(_09253_),
    .A1(_09247_),
    .A2(_09252_));
 sg13g2_and3_1 _15749_ (.X(_09254_),
    .A(net10281),
    .B(_09245_),
    .C(_09253_));
 sg13g2_a21oi_2 _15750_ (.B1(_09254_),
    .Y(_02174_),
    .A2(_09236_),
    .A1(net10285));
 sg13g2_buf_2 place11029 (.A(net11027),
    .X(net11029));
 sg13g2_nand2_1 _15752_ (.Y(_09256_),
    .A(net10651),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[41] ));
 sg13g2_buf_2 place10994 (.A(net10993),
    .X(net10994));
 sg13g2_a22oi_1 _15754_ (.Y(_09258_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[9] ),
    .B2(net10646),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[41] ),
    .A1(net10642));
 sg13g2_nand3_1 _15755_ (.B(_09256_),
    .C(_09258_),
    .A(net10435),
    .Y(_09259_));
 sg13g2_o21ai_1 _15756_ (.B1(_09259_),
    .Y(_09260_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[9] ),
    .A2(net10436));
 sg13g2_and2_1 _15757_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[2] ),
    .B(net10568),
    .X(_09261_));
 sg13g2_nand2_2 _15758_ (.Y(_09262_),
    .A(net10601),
    .B(net10571));
 sg13g2_nand2b_1 _15759_ (.Y(_09263_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[1] ),
    .A_N(net10601));
 sg13g2_buf_2 place10949 (.A(net10935),
    .X(net10949));
 sg13g2_and2_1 _15761_ (.A(_09262_),
    .B(_09263_),
    .X(_09265_));
 sg13g2_buf_2 place10988 (.A(net10987),
    .X(net10988));
 sg13g2_a22oi_1 _15763_ (.Y(_09267_),
    .B1(_09265_),
    .B2(_09016_),
    .A2(_09261_),
    .A1(_09012_));
 sg13g2_nor2_1 _15764_ (.A(_09250_),
    .B(_09267_),
    .Y(_09268_));
 sg13g2_o21ai_1 _15765_ (.B1(net10696),
    .Y(_09269_),
    .A1(_09247_),
    .A2(_09268_));
 sg13g2_buf_2 place10995 (.A(net10993),
    .X(net10995));
 sg13g2_buf_2 place10973 (.A(net10964),
    .X(net10973));
 sg13g2_buf_2 place10948 (.A(net10935),
    .X(net10948));
 sg13g2_xnor2_1 _15769_ (.Y(_09273_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[9] ),
    .B(net10668));
 sg13g2_nand2_1 _15770_ (.Y(_09274_),
    .A(net10672),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[5] ));
 sg13g2_nor4_1 _15771_ (.A(_09064_),
    .B(_09065_),
    .C(_09090_),
    .D(_09274_),
    .Y(_09275_));
 sg13g2_nand2_1 _15772_ (.Y(_09276_),
    .A(net10489),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[5] ));
 sg13g2_nor4_1 _15773_ (.A(_09064_),
    .B(_09065_),
    .C(_09090_),
    .D(_09276_),
    .Y(_09277_));
 sg13g2_nand3_1 _15774_ (.B(net10672),
    .C(net10671),
    .A(net10489),
    .Y(_09278_));
 sg13g2_nand4_1 _15775_ (.B(net10673),
    .C(net10672),
    .A(net10490),
    .Y(_09279_),
    .D(net10671));
 sg13g2_nand4_1 _15776_ (.B(net10489),
    .C(net10673),
    .A(net10490),
    .Y(_09280_),
    .D(net10671));
 sg13g2_nand3_1 _15777_ (.B(_09279_),
    .C(_09280_),
    .A(_09278_),
    .Y(_09281_));
 sg13g2_nand2b_1 _15778_ (.Y(_09282_),
    .B(_09239_),
    .A_N(net10670));
 sg13g2_nor4_1 _15779_ (.A(_09275_),
    .B(_09277_),
    .C(_09281_),
    .D(_09282_),
    .Y(_09283_));
 sg13g2_o21ai_1 _15780_ (.B1(_09283_),
    .Y(_09284_),
    .A1(_09164_),
    .A2(_09166_));
 sg13g2_inv_4 _15781_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[6] ),
    .Y(_09285_));
 sg13g2_nand2_1 _15782_ (.Y(_09286_),
    .A(_09285_),
    .B(_09239_));
 sg13g2_nor4_1 _15783_ (.A(_09275_),
    .B(_09277_),
    .C(_09281_),
    .D(_09286_),
    .Y(_09287_));
 sg13g2_o21ai_1 _15784_ (.B1(_09287_),
    .Y(_09288_),
    .A1(_09164_),
    .A2(_09166_));
 sg13g2_a21oi_1 _15785_ (.A1(_09224_),
    .A2(_09239_),
    .Y(_09289_),
    .B1(_09238_));
 sg13g2_or2_1 _15786_ (.X(_09290_),
    .B(net10669),
    .A(net10488));
 sg13g2_nand4_1 _15787_ (.B(_09288_),
    .C(_09289_),
    .A(_09284_),
    .Y(_09291_),
    .D(_09290_));
 sg13g2_nand2_1 _15788_ (.Y(_09292_),
    .A(net10488),
    .B(net10669));
 sg13g2_nand2_1 _15789_ (.Y(_09293_),
    .A(_09291_),
    .B(_09292_));
 sg13g2_xnor2_1 _15790_ (.Y(_09294_),
    .A(_09273_),
    .B(_09293_));
 sg13g2_a22oi_1 _15791_ (.Y(_09295_),
    .B1(_09294_),
    .B2(net10712),
    .A2(net10521),
    .A1(net10700));
 sg13g2_and3_1 _15792_ (.X(_09296_),
    .A(net10281),
    .B(_09269_),
    .C(_09295_));
 sg13g2_a21oi_2 _15793_ (.B1(_09296_),
    .Y(_02175_),
    .A2(_09260_),
    .A1(net10285));
 sg13g2_buf_2 place10816 (.A(net10815),
    .X(net10816));
 sg13g2_buf_2 place11033 (.A(net11032),
    .X(net11033));
 sg13g2_buf_2 place10823 (.A(net10822),
    .X(net10823));
 sg13g2_nand2_1 _15797_ (.Y(_09300_),
    .A(net10650),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[42] ));
 sg13g2_buf_16 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_8_52_0_clk));
 sg13g2_a22oi_1 _15799_ (.Y(_09302_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[10] ),
    .B2(net10646),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[42] ),
    .A1(net10642));
 sg13g2_nand3_1 _15800_ (.B(_09300_),
    .C(_09302_),
    .A(net10434),
    .Y(_09303_));
 sg13g2_o21ai_1 _15801_ (.B1(_09303_),
    .Y(_09304_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[10] ),
    .A2(net10435));
 sg13g2_nand2b_2 _15802_ (.Y(_09305_),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_is_lb ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.latched_is_lh ));
 sg13g2_buf_2 place11019 (.A(net11018),
    .X(net11019));
 sg13g2_nand2b_1 _15804_ (.Y(_09307_),
    .B(_09265_),
    .A_N(_09046_));
 sg13g2_o21ai_1 _15805_ (.B1(_09307_),
    .Y(_09308_),
    .A1(_09042_),
    .A2(_09262_));
 sg13g2_and2_1 _15806_ (.A(_09305_),
    .B(_09308_),
    .X(_09309_));
 sg13g2_o21ai_1 _15807_ (.B1(net10696),
    .Y(_09310_),
    .A1(_09247_),
    .A2(_09309_));
 sg13g2_buf_2 place11018 (.A(net11014),
    .X(net11018));
 sg13g2_and2_1 _15809_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[9] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[9] ),
    .X(_09312_));
 sg13g2_buf_2 place11026 (.A(net11025),
    .X(net11026));
 sg13g2_nor2_1 _15811_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[9] ),
    .B(net10668),
    .Y(_09314_));
 sg13g2_a21oi_2 _15812_ (.B1(_09314_),
    .Y(_09315_),
    .A2(_09292_),
    .A1(_09291_));
 sg13g2_or2_1 _15813_ (.X(_09316_),
    .B(_09315_),
    .A(_09312_));
 sg13g2_buf_2 place11034 (.A(net11033),
    .X(net11034));
 sg13g2_buf_16 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_8_48_0_clk));
 sg13g2_buf_2 place11031 (.A(net11030),
    .X(net11031));
 sg13g2_buf_16 clkbuf_leaf_83_clk (.X(clknet_leaf_83_clk),
    .A(clknet_8_3_0_clk));
 sg13g2_xnor2_1 _15818_ (.Y(_09321_),
    .A(net10498),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[10] ));
 sg13g2_xnor2_1 _15819_ (.Y(_09322_),
    .A(_09316_),
    .B(_09321_));
 sg13g2_a22oi_1 _15820_ (.Y(_09323_),
    .B1(_09322_),
    .B2(net10710),
    .A2(net10594),
    .A1(net10700));
 sg13g2_and3_1 _15821_ (.X(_09324_),
    .A(_08997_),
    .B(_09310_),
    .C(_09323_));
 sg13g2_a21oi_1 _15822_ (.A1(net10285),
    .A2(_09304_),
    .Y(_02145_),
    .B1(_09324_));
 sg13g2_buf_2 place11027 (.A(net11026),
    .X(net11027));
 sg13g2_nor2_1 _15824_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[10] ),
    .B(_09316_),
    .Y(_09326_));
 sg13g2_a21oi_1 _15825_ (.A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[10] ),
    .A2(_09316_),
    .Y(_09327_),
    .B1(net10498));
 sg13g2_nor2_2 _15826_ (.A(_09326_),
    .B(_09327_),
    .Y(_09328_));
 sg13g2_buf_2 place10814 (.A(net10813),
    .X(net10814));
 sg13g2_buf_2 place11021 (.A(net11020),
    .X(net11021));
 sg13g2_xnor2_1 _15829_ (.Y(_09331_),
    .A(net10497),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[11] ));
 sg13g2_xnor2_1 _15830_ (.Y(_09332_),
    .A(_09328_),
    .B(_09331_));
 sg13g2_nand2b_1 _15831_ (.Y(_09333_),
    .B(_09265_),
    .A_N(_09078_));
 sg13g2_o21ai_1 _15832_ (.B1(_09333_),
    .Y(_09334_),
    .A1(_09074_),
    .A2(_09262_));
 sg13g2_and2_1 _15833_ (.A(_09305_),
    .B(_09334_),
    .X(_09335_));
 sg13g2_o21ai_1 _15834_ (.B1(\u_ac_controller_soc_inst.u_picorv32.cpu_state[6] ),
    .Y(_09336_),
    .A1(_09247_),
    .A2(_09335_));
 sg13g2_inv_1 _15835_ (.Y(_09337_),
    .A(_09336_));
 sg13g2_a221oi_1 _15836_ (.B2(net10711),
    .C1(_09337_),
    .B1(_09332_),
    .A1(net10699),
    .Y(_09338_),
    .A2(net10592));
 sg13g2_buf_2 place11036 (.A(net11035),
    .X(net11036));
 sg13g2_nand2b_1 _15838_ (.Y(_09340_),
    .B(net10395),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.count_cycle[11] ));
 sg13g2_buf_16 clkbuf_leaf_82_clk (.X(clknet_leaf_82_clk),
    .A(clknet_8_3_0_clk));
 sg13g2_nand2_1 _15840_ (.Y(_09342_),
    .A(net10650),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[43] ));
 sg13g2_buf_2 place10822 (.A(net10816),
    .X(net10822));
 sg13g2_a22oi_1 _15842_ (.Y(_09344_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[11] ),
    .B2(net10645),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[43] ),
    .A1(net10641));
 sg13g2_nand3_1 _15843_ (.B(_09342_),
    .C(_09344_),
    .A(net10434),
    .Y(_09345_));
 sg13g2_a21oi_2 _15844_ (.B1(net10282),
    .Y(_09346_),
    .A2(_09345_),
    .A1(_09340_));
 sg13g2_a21oi_1 _15845_ (.A1(_08997_),
    .A2(_09338_),
    .Y(_02146_),
    .B1(_09346_));
 sg13g2_buf_2 place11025 (.A(net11018),
    .X(net11025));
 sg13g2_inv_1 _16345__11058 (.Y(net11058),
    .A(clknet_leaf_284_clk));
 sg13g2_a21o_1 _15848_ (.A2(_09328_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[11] ),
    .B1(net10497),
    .X(_09349_));
 sg13g2_o21ai_1 _15849_ (.B1(_09349_),
    .Y(_09350_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[11] ),
    .A2(_09328_));
 sg13g2_buf_16 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_8_49_0_clk));
 sg13g2_buf_2 place11022 (.A(net11020),
    .X(net11022));
 sg13g2_buf_2 place11023 (.A(net11022),
    .X(net11023));
 sg13g2_xnor2_1 _15853_ (.Y(_09354_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[12] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[12] ));
 sg13g2_xor2_1 _15854_ (.B(_09354_),
    .A(_09350_),
    .X(_09355_));
 sg13g2_nand2b_1 _15855_ (.Y(_09356_),
    .B(_09265_),
    .A_N(_08470_));
 sg13g2_o21ai_1 _15856_ (.B1(_09356_),
    .Y(_09357_),
    .A1(_09106_),
    .A2(_09262_));
 sg13g2_a21oi_1 _15857_ (.A1(_09305_),
    .A2(_09357_),
    .Y(_09358_),
    .B1(_09247_));
 sg13g2_nor2_1 _15858_ (.A(net10460),
    .B(_09358_),
    .Y(_09359_));
 sg13g2_a221oi_1 _15859_ (.B2(net10710),
    .C1(_09359_),
    .B1(_09355_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpu_state[4] ),
    .Y(_09360_),
    .A2(net10590));
 sg13g2_inv_1 _16345__11059 (.Y(net11059),
    .A(clknet_8_68_0_clk));
 sg13g2_nand2b_1 _15861_ (.Y(_09362_),
    .B(net10395),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.count_cycle[12] ));
 sg13g2_nand2_1 _15862_ (.Y(_09363_),
    .A(net10650),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[44] ));
 sg13g2_buf_2 place10924 (.A(net10923),
    .X(net10924));
 sg13g2_buf_2 place10917 (.A(net10916),
    .X(net10917));
 sg13g2_a22oi_1 _15865_ (.Y(_09366_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[12] ),
    .B2(net10646),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[44] ),
    .A1(net10642));
 sg13g2_nand3_1 _15866_ (.B(_09363_),
    .C(_09366_),
    .A(net10434),
    .Y(_09367_));
 sg13g2_a21oi_2 _15867_ (.B1(net10282),
    .Y(_09368_),
    .A2(_09367_),
    .A1(_09362_));
 sg13g2_a21oi_2 _15868_ (.B1(_09368_),
    .Y(_02147_),
    .A2(_09360_),
    .A1(_08997_));
 sg13g2_buf_2 place10926 (.A(net10925),
    .X(net10926));
 sg13g2_inv_1 _16345__11061 (.Y(net11061),
    .A(clknet_leaf_235_clk));
 sg13g2_xor2_1 _15871_ (.B(net10691),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[13] ),
    .X(_09371_));
 sg13g2_nor2_1 _15872_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[12] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[12] ),
    .Y(_09372_));
 sg13g2_nand2_1 _15873_ (.Y(_09373_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[12] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[12] ));
 sg13g2_o21ai_1 _15874_ (.B1(_09373_),
    .Y(_09374_),
    .A1(_09350_),
    .A2(_09372_));
 sg13g2_xnor2_1 _15875_ (.Y(_09375_),
    .A(_09371_),
    .B(_09374_));
 sg13g2_nand2_2 _15876_ (.Y(_09376_),
    .A(net10713),
    .B(net10283));
 sg13g2_buf_2 place11035 (.A(net11034),
    .X(net11035));
 sg13g2_a221oi_1 _15878_ (.B2(\u_ac_controller_soc_inst.io_rdata[29] ),
    .C1(_09146_),
    .B1(net10183),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[29] ),
    .Y(_09378_),
    .A2(net10243));
 sg13g2_nand2b_1 _15879_ (.Y(_09379_),
    .B(_09265_),
    .A_N(_08464_));
 sg13g2_o21ai_1 _15880_ (.B1(_09379_),
    .Y(_09380_),
    .A1(_09378_),
    .A2(_09262_));
 sg13g2_a21o_1 _15881_ (.A2(_09380_),
    .A1(_09305_),
    .B1(_09247_),
    .X(_09381_));
 sg13g2_buf_2 place10921 (.A(net10920),
    .X(net10921));
 sg13g2_nand2_1 _15883_ (.Y(_09383_),
    .A(net10650),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[45] ));
 sg13g2_a22oi_1 _15884_ (.Y(_09384_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[13] ),
    .B2(net10646),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[45] ),
    .A1(net10642));
 sg13g2_nand3_1 _15885_ (.B(_09383_),
    .C(_09384_),
    .A(net10434),
    .Y(_09385_));
 sg13g2_o21ai_1 _15886_ (.B1(_09385_),
    .Y(_09386_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[13] ),
    .A2(net10434));
 sg13g2_nor2_2 _15887_ (.A(net10282),
    .B(_09386_),
    .Y(_09387_));
 sg13g2_a221oi_1 _15888_ (.B2(\u_ac_controller_soc_inst.u_picorv32.cpu_state[6] ),
    .C1(_09387_),
    .B1(_09381_),
    .A1(net10708),
    .Y(_09388_),
    .A2(net10587));
 sg13g2_o21ai_1 _15889_ (.B1(_09388_),
    .Y(_02148_),
    .A1(_09375_),
    .A2(_09376_));
 sg13g2_buf_2 place10925 (.A(net10924),
    .X(net10925));
 sg13g2_inv_1 _16345__11060 (.Y(net11060),
    .A(clknet_leaf_235_clk));
 sg13g2_nand2_1 _15892_ (.Y(_09391_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycleh ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[46] ));
 sg13g2_buf_16 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_8_48_0_clk));
 sg13g2_a22oi_1 _15894_ (.Y(_09393_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[14] ),
    .B2(net10645),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[46] ),
    .A1(net10641));
 sg13g2_nand3_1 _15895_ (.B(_09391_),
    .C(_09393_),
    .A(net10433),
    .Y(_09394_));
 sg13g2_o21ai_1 _15896_ (.B1(_09394_),
    .Y(_09395_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[14] ),
    .A2(net10433));
 sg13g2_nand2b_1 _15897_ (.Y(_09396_),
    .B(_09261_),
    .A_N(_09178_));
 sg13g2_nand2b_1 _15898_ (.Y(_09397_),
    .B(_09265_),
    .A_N(_08476_));
 sg13g2_a21oi_1 _15899_ (.A1(_09396_),
    .A2(_09397_),
    .Y(_09398_),
    .B1(_09250_));
 sg13g2_o21ai_1 _15900_ (.B1(net10696),
    .Y(_09399_),
    .A1(_09247_),
    .A2(_09398_));
 sg13g2_buf_16 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_8_50_0_clk));
 sg13g2_nor2_1 _15902_ (.A(_09331_),
    .B(_09354_),
    .Y(_09401_));
 sg13g2_nand2_2 _15903_ (.Y(_09402_),
    .A(_09371_),
    .B(_09401_));
 sg13g2_nor4_1 _15904_ (.A(_09243_),
    .B(_09273_),
    .C(_09321_),
    .D(_09402_),
    .Y(_09403_));
 sg13g2_nor2_1 _15905_ (.A(net10498),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[10] ),
    .Y(_09404_));
 sg13g2_a21oi_1 _15906_ (.A1(net10488),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[8] ),
    .Y(_09405_),
    .B1(_09312_));
 sg13g2_nand2_1 _15907_ (.Y(_09406_),
    .A(net10498),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[10] ));
 sg13g2_o21ai_1 _15908_ (.B1(_09406_),
    .Y(_09407_),
    .A1(_09314_),
    .A2(_09405_));
 sg13g2_nor2b_1 _15909_ (.A(_09404_),
    .B_N(_09407_),
    .Y(_09408_));
 sg13g2_a21o_1 _15910_ (.A2(_09408_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[11] ),
    .B1(net10497),
    .X(_09409_));
 sg13g2_o21ai_1 _15911_ (.B1(_09409_),
    .Y(_09410_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[11] ),
    .A2(_09408_));
 sg13g2_o21ai_1 _15912_ (.B1(_09373_),
    .Y(_09411_),
    .A1(_09372_),
    .A2(_09410_));
 sg13g2_a21o_1 _15913_ (.A2(_09411_),
    .A1(net10691),
    .B1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[13] ),
    .X(_09412_));
 sg13g2_or2_1 _15914_ (.X(_09413_),
    .B(_09411_),
    .A(net10691));
 sg13g2_a22oi_1 _15915_ (.Y(_09414_),
    .B1(_09412_),
    .B2(_09413_),
    .A2(_09403_),
    .A1(_09240_));
 sg13g2_buf_16 clkbuf_leaf_137_clk (.X(clknet_leaf_137_clk),
    .A(clknet_8_30_0_clk));
 sg13g2_buf_16 clkbuf_leaf_136_clk (.X(clknet_leaf_136_clk),
    .A(clknet_8_244_0_clk));
 sg13g2_xor2_1 _15918_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[14] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[14] ),
    .X(_09417_));
 sg13g2_xnor2_1 _15919_ (.Y(_09418_),
    .A(_09414_),
    .B(_09417_));
 sg13g2_a22oi_1 _15920_ (.Y(_09419_),
    .B1(_09418_),
    .B2(net10710),
    .A2(net10585),
    .A1(net10700));
 sg13g2_and3_1 _15921_ (.X(_09420_),
    .A(_08997_),
    .B(_09399_),
    .C(_09419_));
 sg13g2_a21oi_1 _15922_ (.A1(_08945_),
    .A2(_09395_),
    .Y(_02149_),
    .B1(_09420_));
 sg13g2_buf_16 clkbuf_leaf_62_clk (.X(clknet_leaf_62_clk),
    .A(clknet_8_7_0_clk));
 sg13g2_nand2_1 _15924_ (.Y(_09422_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycleh ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[47] ));
 sg13g2_buf_2 place10952 (.A(net10950),
    .X(net10952));
 sg13g2_a22oi_1 _15926_ (.Y(_09424_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[15] ),
    .B2(net10645),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[47] ),
    .A1(net10641));
 sg13g2_nand3_1 _15927_ (.B(_09422_),
    .C(_09424_),
    .A(net10433),
    .Y(_09425_));
 sg13g2_o21ai_1 _15928_ (.B1(_09425_),
    .Y(_09426_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[15] ),
    .A2(net10433));
 sg13g2_nand2_1 _15929_ (.Y(_09427_),
    .A(net10497),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[11] ));
 sg13g2_o21ai_1 _15930_ (.B1(_09373_),
    .Y(_09428_),
    .A1(_09372_),
    .A2(_09427_));
 sg13g2_a21oi_1 _15931_ (.A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[13] ),
    .A2(_09428_),
    .Y(_09429_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[13] ));
 sg13g2_nor2_1 _15932_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[13] ),
    .B(_09428_),
    .Y(_09430_));
 sg13g2_nand2_1 _15933_ (.Y(_09431_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[14] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[14] ));
 sg13g2_o21ai_1 _15934_ (.B1(_09431_),
    .Y(_09432_),
    .A1(_09429_),
    .A2(_09430_));
 sg13g2_inv_1 _15935_ (.Y(_09433_),
    .A(_09432_));
 sg13g2_nand2b_2 _15936_ (.Y(_09434_),
    .B(_09406_),
    .A_N(_09312_));
 sg13g2_nor2_2 _15937_ (.A(_09402_),
    .B(_09404_),
    .Y(_09435_));
 sg13g2_o21ai_1 _15938_ (.B1(_09435_),
    .Y(_09436_),
    .A1(_09315_),
    .A2(_09434_));
 sg13g2_nor2_1 _15939_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[14] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[14] ),
    .Y(_09437_));
 sg13g2_a21oi_2 _15940_ (.B1(_09437_),
    .Y(_09438_),
    .A2(_09436_),
    .A1(_09433_));
 sg13g2_buf_2 place11037 (.A(resetn),
    .X(net11037));
 sg13g2_buf_2 place10972 (.A(net10970),
    .X(net10972));
 sg13g2_xnor2_1 _15943_ (.Y(_09441_),
    .A(net10496),
    .B(net10690));
 sg13g2_xnor2_1 _15944_ (.Y(_09442_),
    .A(_09438_),
    .B(_09441_));
 sg13g2_nand2_1 _15945_ (.Y(_09443_),
    .A(net10709),
    .B(_09442_));
 sg13g2_buf_2 place10951 (.A(net10950),
    .X(net10951));
 sg13g2_o21ai_1 _15947_ (.B1(\u_ac_controller_soc_inst.u_picorv32.latched_is_lb ),
    .Y(_09445_),
    .A1(_09212_),
    .A2(_09218_));
 sg13g2_a22oi_1 _15948_ (.Y(_09446_),
    .B1(_08973_),
    .B2(_09208_),
    .A2(_08483_),
    .A1(_08969_));
 sg13g2_nor2_1 _15949_ (.A(_00052_),
    .B(_09446_),
    .Y(_09447_));
 sg13g2_a21oi_1 _15950_ (.A1(_08483_),
    .A2(net10399),
    .Y(_09448_),
    .B1(_09447_));
 sg13g2_mux2_1 _15951_ (.A0(\u_ac_controller_soc_inst.u_picorv32.latched_is_lb ),
    .A1(_09448_),
    .S(\u_ac_controller_soc_inst.u_picorv32.latched_is_lh ),
    .X(_09449_));
 sg13g2_a21oi_2 _15952_ (.B1(_07949_),
    .Y(_09450_),
    .A2(_09449_),
    .A1(_09445_));
 sg13g2_buf_2 place10901 (.A(net10900),
    .X(net10901));
 sg13g2_buf_2 place11043 (.A(net11041),
    .X(net11043));
 sg13g2_nor2_2 _15955_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_is_lh ),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_is_lb ),
    .Y(_09453_));
 sg13g2_buf_2 place10900 (.A(net10893),
    .X(net10900));
 sg13g2_nand2_1 _15957_ (.Y(_09455_),
    .A(_09453_),
    .B(_09448_));
 sg13g2_a22oi_1 _15958_ (.Y(_09456_),
    .B1(_09450_),
    .B2(_09455_),
    .A2(net10583),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpu_state[4] ));
 sg13g2_and3_1 _15959_ (.X(_09457_),
    .A(net10283),
    .B(_09443_),
    .C(_09456_));
 sg13g2_a21oi_1 _15960_ (.A1(net10286),
    .A2(_09426_),
    .Y(_02150_),
    .B1(_09457_));
 sg13g2_buf_2 place11000 (.A(net10997),
    .X(net11000));
 sg13g2_nand2_1 _15962_ (.Y(_09459_),
    .A(net10648),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[48] ));
 sg13g2_buf_2 place11039 (.A(net11038),
    .X(net11039));
 sg13g2_buf_2 place10971 (.A(net10970),
    .X(net10971));
 sg13g2_a22oi_1 _15965_ (.Y(_09462_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[16] ),
    .B2(net10643),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[48] ),
    .A1(net10639));
 sg13g2_nand3_1 _15966_ (.B(_09459_),
    .C(_09462_),
    .A(_08320_),
    .Y(_09463_));
 sg13g2_o21ai_1 _15967_ (.B1(_09463_),
    .Y(_09464_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[16] ),
    .A2(net10433));
 sg13g2_nor2_1 _15968_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[15] ),
    .B(_09438_),
    .Y(_09465_));
 sg13g2_a21oi_1 _15969_ (.A1(net10690),
    .A2(_09438_),
    .Y(_09466_),
    .B1(net10496));
 sg13g2_nor2_1 _15970_ (.A(_09465_),
    .B(_09466_),
    .Y(_09467_));
 sg13g2_buf_16 clkbuf_leaf_134_clk (.X(clknet_leaf_134_clk),
    .A(clknet_8_30_0_clk));
 sg13g2_buf_2 place11042 (.A(net11041),
    .X(net11042));
 sg13g2_xnor2_1 _15973_ (.Y(_09470_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[16] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[16] ));
 sg13g2_xor2_1 _15974_ (.B(_09470_),
    .A(_09467_),
    .X(_09471_));
 sg13g2_buf_2 place10999 (.A(net10998),
    .X(net10999));
 sg13g2_buf_2 place10998 (.A(net10997),
    .X(net10998));
 sg13g2_o21ai_1 _15977_ (.B1(net10393),
    .Y(_09474_),
    .A1(_08495_),
    .A2(net10405));
 sg13g2_a22oi_1 _15978_ (.Y(_09475_),
    .B1(_09450_),
    .B2(_09474_),
    .A2(net10581),
    .A1(net10697));
 sg13g2_o21ai_1 _15979_ (.B1(_09475_),
    .Y(_09476_),
    .A1(_08395_),
    .A2(_09471_));
 sg13g2_nor2_1 _15980_ (.A(net10286),
    .B(_09476_),
    .Y(_09477_));
 sg13g2_a21oi_1 _15981_ (.A1(net10286),
    .A2(_09464_),
    .Y(_02151_),
    .B1(_09477_));
 sg13g2_buf_2 place10895 (.A(net10894),
    .X(net10895));
 sg13g2_buf_2 place11057 (.A(net11056),
    .X(net11057));
 sg13g2_buf_2 place10950 (.A(_00005_),
    .X(net10950));
 sg13g2_buf_2 place10899 (.A(net10897),
    .X(net10899));
 sg13g2_xor2_1 _15986_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[17] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[17] ),
    .X(_09482_));
 sg13g2_or2_1 _15987_ (.X(_09483_),
    .B(net10689),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[16] ));
 sg13g2_and2_1 _15988_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[16] ),
    .B(net10689),
    .X(_09484_));
 sg13g2_a21oi_1 _15989_ (.A1(_09467_),
    .A2(_09483_),
    .Y(_09485_),
    .B1(_09484_));
 sg13g2_xnor2_1 _15990_ (.Y(_09486_),
    .A(_09482_),
    .B(_09485_));
 sg13g2_nand2_1 _15991_ (.Y(_09487_),
    .A(net10709),
    .B(_09486_));
 sg13g2_buf_16 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_8_0_0_clk));
 sg13g2_buf_2 place11048 (.A(net11037),
    .X(net11048));
 sg13g2_or2_1 _15994_ (.X(_09490_),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_is_lb ),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_is_lh ));
 sg13g2_buf_2 place11050 (.A(net11048),
    .X(net11050));
 sg13g2_a21o_1 _15996_ (.A2(net10399),
    .A1(_08506_),
    .B1(_09490_),
    .X(_09492_));
 sg13g2_a221oi_1 _15997_ (.B2(_09492_),
    .C1(net10286),
    .B1(_09450_),
    .A1(net10697),
    .Y(_09493_),
    .A2(net10578));
 sg13g2_buf_2 place11055 (.A(net11054),
    .X(net11055));
 sg13g2_buf_16 clkbuf_leaf_131_clk (.X(clknet_leaf_131_clk),
    .A(clknet_8_149_0_clk));
 sg13g2_nand2_1 _16000_ (.Y(_09496_),
    .A(net10648),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[49] ));
 sg13g2_buf_2 place11056 (.A(net11037),
    .X(net11056));
 sg13g2_a22oi_1 _16002_ (.Y(_09498_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[17] ),
    .B2(net10643),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[49] ),
    .A1(net10639));
 sg13g2_nand3_1 _16003_ (.B(_09496_),
    .C(_09498_),
    .A(net10430),
    .Y(_09499_));
 sg13g2_o21ai_1 _16004_ (.B1(_09499_),
    .Y(_09500_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[17] ),
    .A2(net10430));
 sg13g2_a22oi_1 _16005_ (.Y(_02152_),
    .B1(_09500_),
    .B2(net10286),
    .A2(_09493_),
    .A1(_09487_));
 sg13g2_buf_2 place11041 (.A(net11040),
    .X(net11041));
 sg13g2_nand2b_1 _16007_ (.Y(_09502_),
    .B(_09117_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.count_cycle[18] ));
 sg13g2_buf_16 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_8_5_0_clk));
 sg13g2_nand2_1 _16009_ (.Y(_09504_),
    .A(net10647),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[50] ));
 sg13g2_buf_2 place11046 (.A(net11041),
    .X(net11046));
 sg13g2_buf_2 place11047 (.A(net11046),
    .X(net11047));
 sg13g2_a22oi_1 _16012_ (.Y(_09507_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[18] ),
    .B2(net10643),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[50] ),
    .A1(net10639));
 sg13g2_nand3_1 _16013_ (.B(_09504_),
    .C(_09507_),
    .A(net10430),
    .Y(_09508_));
 sg13g2_a21oi_2 _16014_ (.B1(net10284),
    .Y(_09509_),
    .A2(_09508_),
    .A1(_09502_));
 sg13g2_o21ai_1 _16015_ (.B1(net10393),
    .Y(_09510_),
    .A1(_08510_),
    .A2(net10405));
 sg13g2_nand2_1 _16016_ (.Y(_09511_),
    .A(net9697),
    .B(_09510_));
 sg13g2_buf_16 clkbuf_leaf_78_clk (.X(clknet_leaf_78_clk),
    .A(clknet_8_11_0_clk));
 sg13g2_nand2_1 _16018_ (.Y(_09513_),
    .A(net10697),
    .B(net10576));
 sg13g2_and2_1 _16019_ (.A(_09511_),
    .B(_09513_),
    .X(_09514_));
 sg13g2_nor2_1 _16020_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[17] ),
    .B(net10688),
    .Y(_09515_));
 sg13g2_nand2_1 _16021_ (.Y(_09516_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[17] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[17] ));
 sg13g2_o21ai_1 _16022_ (.B1(_09516_),
    .Y(_09517_),
    .A1(_09485_),
    .A2(_09515_));
 sg13g2_buf_2 place11049 (.A(net11048),
    .X(net11049));
 sg13g2_buf_16 clkbuf_leaf_72_clk (.X(clknet_leaf_72_clk),
    .A(clknet_8_18_0_clk));
 sg13g2_xor2_1 _16025_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[18] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[18] ),
    .X(_09520_));
 sg13g2_and4_1 _16026_ (.A(net10283),
    .B(_09514_),
    .C(_09517_),
    .D(_09520_),
    .X(_09521_));
 sg13g2_nand2_1 _16027_ (.Y(_09522_),
    .A(_09511_),
    .B(_09513_));
 sg13g2_nor4_1 _16028_ (.A(net10286),
    .B(_09522_),
    .C(_09517_),
    .D(_09520_),
    .Y(_09523_));
 sg13g2_nor3_1 _16029_ (.A(net10709),
    .B(net10286),
    .C(_09522_),
    .Y(_09524_));
 sg13g2_nor4_1 _16030_ (.A(_09509_),
    .B(_09521_),
    .C(_09523_),
    .D(_09524_),
    .Y(_02153_));
 sg13g2_nand2_1 _16031_ (.Y(_09525_),
    .A(net10647),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[51] ));
 sg13g2_buf_16 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_8_0_0_clk));
 sg13g2_buf_2 place11038 (.A(net11037),
    .X(net11038));
 sg13g2_a22oi_1 _16034_ (.Y(_09528_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[19] ),
    .B2(net10643),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[51] ),
    .A1(net10639));
 sg13g2_nand3_1 _16035_ (.B(_09525_),
    .C(_09528_),
    .A(net10430),
    .Y(_09529_));
 sg13g2_o21ai_1 _16036_ (.B1(_09529_),
    .Y(_09530_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[19] ),
    .A2(net10430));
 sg13g2_and2_1 _16037_ (.A(net10496),
    .B(net10690),
    .X(_09531_));
 sg13g2_a221oi_1 _16038_ (.B2(_09531_),
    .C1(_09484_),
    .B1(_09483_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[17] ),
    .Y(_09532_),
    .A2(net10688));
 sg13g2_nor2_1 _16039_ (.A(_09515_),
    .B(_09532_),
    .Y(_09533_));
 sg13g2_a21o_1 _16040_ (.A2(_09533_),
    .A1(net10687),
    .B1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[18] ),
    .X(_09534_));
 sg13g2_or2_1 _16041_ (.X(_09535_),
    .B(_09533_),
    .A(net10687));
 sg13g2_nand2_1 _16042_ (.Y(_09536_),
    .A(_09482_),
    .B(_09520_));
 sg13g2_nor4_1 _16043_ (.A(_09437_),
    .B(_09441_),
    .C(_09470_),
    .D(_09536_),
    .Y(_09537_));
 sg13g2_a22oi_1 _16044_ (.Y(_09538_),
    .B1(_09537_),
    .B2(_09432_),
    .A2(_09535_),
    .A1(_09534_));
 sg13g2_and2_1 _16045_ (.A(_09435_),
    .B(_09537_),
    .X(_09539_));
 sg13g2_o21ai_1 _16046_ (.B1(_09539_),
    .Y(_09540_),
    .A1(_09315_),
    .A2(_09434_));
 sg13g2_nand2_2 _16047_ (.Y(_09541_),
    .A(_09538_),
    .B(_09540_));
 sg13g2_buf_2 place10928 (.A(net10927),
    .X(net10928));
 sg13g2_buf_2 place10923 (.A(net10919),
    .X(net10923));
 sg13g2_xnor2_1 _16050_ (.Y(_09544_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[19] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[19] ));
 sg13g2_xnor2_1 _16051_ (.Y(_09545_),
    .A(_09541_),
    .B(_09544_));
 sg13g2_nand2_1 _16052_ (.Y(_09546_),
    .A(net10713),
    .B(_09545_));
 sg13g2_buf_2 place11044 (.A(net11043),
    .X(net11044));
 sg13g2_o21ai_1 _16054_ (.B1(net10393),
    .Y(_09548_),
    .A1(_08515_),
    .A2(net10405));
 sg13g2_a22oi_1 _16055_ (.Y(_09549_),
    .B1(net9697),
    .B2(_09548_),
    .A2(net10574),
    .A1(net10697));
 sg13g2_and3_2 _16056_ (.X(_09550_),
    .A(net10284),
    .B(_09546_),
    .C(_09549_));
 sg13g2_a21oi_1 _16057_ (.A1(net10288),
    .A2(_09530_),
    .Y(_02154_),
    .B1(_09550_));
 sg13g2_buf_16 clkbuf_leaf_61_clk (.X(clknet_leaf_61_clk),
    .A(clknet_8_6_0_clk));
 sg13g2_nand2_1 _16059_ (.Y(_09552_),
    .A(net10649),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[52] ));
 sg13g2_buf_2 place11045 (.A(net11044),
    .X(net11045));
 sg13g2_a22oi_1 _16061_ (.Y(_09554_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[20] ),
    .B2(net10643),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[52] ),
    .A1(net10639));
 sg13g2_nand3_1 _16062_ (.B(_09552_),
    .C(_09554_),
    .A(net10432),
    .Y(_09555_));
 sg13g2_o21ai_1 _16063_ (.B1(_09555_),
    .Y(_09556_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[20] ),
    .A2(net10431));
 sg13g2_buf_16 clkbuf_leaf_65_clk (.X(clknet_leaf_65_clk),
    .A(clknet_8_7_0_clk));
 sg13g2_nand2_1 _16065_ (.Y(_09558_),
    .A(net10698),
    .B(net10567));
 sg13g2_buf_16 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_8_53_0_clk));
 sg13g2_buf_16 clkbuf_leaf_70_clk (.X(clknet_leaf_70_clk),
    .A(clknet_8_18_0_clk));
 sg13g2_and2_1 _16068_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[20] ),
    .B(net10685),
    .X(_09561_));
 sg13g2_buf_16 clkbuf_leaf_71_clk (.X(clknet_leaf_71_clk),
    .A(clknet_8_18_0_clk));
 sg13g2_buf_16 clkbuf_leaf_63_clk (.X(clknet_leaf_63_clk),
    .A(clknet_8_7_0_clk));
 sg13g2_nor2_2 _16071_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[20] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[20] ),
    .Y(_09564_));
 sg13g2_nor2_1 _16072_ (.A(_09561_),
    .B(_09564_),
    .Y(_09565_));
 sg13g2_or2_1 _16073_ (.X(_09566_),
    .B(net10686),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[19] ));
 sg13g2_buf_16 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_8_1_0_clk));
 sg13g2_and2_1 _16075_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[19] ),
    .B(net10686),
    .X(_09568_));
 sg13g2_buf_2 place10893 (.A(_00006_),
    .X(net10893));
 sg13g2_a21oi_1 _16077_ (.A1(_09541_),
    .A2(_09566_),
    .Y(_09570_),
    .B1(_09568_));
 sg13g2_xnor2_1 _16078_ (.Y(_09571_),
    .A(_09565_),
    .B(_09570_));
 sg13g2_o21ai_1 _16079_ (.B1(net10393),
    .Y(_09572_),
    .A1(_08522_),
    .A2(net10405));
 sg13g2_a22oi_1 _16080_ (.Y(_09573_),
    .B1(_09572_),
    .B2(net9697),
    .A2(_09571_),
    .A1(net10709));
 sg13g2_and3_2 _16081_ (.X(_09574_),
    .A(net10283),
    .B(_09558_),
    .C(_09573_));
 sg13g2_a21oi_1 _16082_ (.A1(net10288),
    .A2(_09556_),
    .Y(_02156_),
    .B1(_09574_));
 sg13g2_buf_2 place11003 (.A(_08213_),
    .X(net11003));
 sg13g2_nand2_1 _16084_ (.Y(_09576_),
    .A(net10649),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[53] ));
 sg13g2_buf_16 clkbuf_leaf_73_clk (.X(clknet_leaf_73_clk),
    .A(clknet_8_18_0_clk));
 sg13g2_a22oi_1 _16086_ (.Y(_09578_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[21] ),
    .B2(net10644),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[53] ),
    .A1(net10640));
 sg13g2_nand3_1 _16087_ (.B(_09576_),
    .C(_09578_),
    .A(net10432),
    .Y(_09579_));
 sg13g2_o21ai_1 _16088_ (.B1(_09579_),
    .Y(_09580_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[21] ),
    .A2(net10431));
 sg13g2_a221oi_1 _16089_ (.B2(_09566_),
    .C1(_09568_),
    .B1(_09541_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[20] ),
    .Y(_09581_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[20] ));
 sg13g2_nor2_1 _16090_ (.A(_09564_),
    .B(_09581_),
    .Y(_09582_));
 sg13g2_buf_2 place11014 (.A(net11013),
    .X(net11014));
 sg13g2_buf_2 place10978 (.A(net10977),
    .X(net10978));
 sg13g2_buf_2 place11016 (.A(net11015),
    .X(net11016));
 sg13g2_xnor2_1 _16094_ (.Y(_09586_),
    .A(net10495),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[21] ));
 sg13g2_xor2_1 _16095_ (.B(_09586_),
    .A(_09582_),
    .X(_09587_));
 sg13g2_buf_2 place11013 (.A(net11004),
    .X(net11013));
 sg13g2_buf_2 place11012 (.A(net11009),
    .X(net11012));
 sg13g2_o21ai_1 _16098_ (.B1(net10393),
    .Y(_09590_),
    .A1(_08531_),
    .A2(net10405));
 sg13g2_a22oi_1 _16099_ (.Y(_09591_),
    .B1(net9697),
    .B2(_09590_),
    .A2(net10565),
    .A1(net10697));
 sg13g2_o21ai_1 _16100_ (.B1(_09591_),
    .Y(_09592_),
    .A1(_08395_),
    .A2(_09587_));
 sg13g2_nor2_1 _16101_ (.A(net10287),
    .B(_09592_),
    .Y(_09593_));
 sg13g2_a21oi_1 _16102_ (.A1(net10288),
    .A2(_09580_),
    .Y(_02157_),
    .B1(_09593_));
 sg13g2_buf_2 place11015 (.A(net11014),
    .X(net11015));
 sg13g2_nand2_1 _16104_ (.Y(_09595_),
    .A(net10649),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[54] ));
 sg13g2_buf_2 place10970 (.A(net10964),
    .X(net10970));
 sg13g2_a22oi_1 _16106_ (.Y(_09597_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[22] ),
    .B2(net10644),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[54] ),
    .A1(net10640));
 sg13g2_nand3_1 _16107_ (.B(_09595_),
    .C(_09597_),
    .A(net10432),
    .Y(_09598_));
 sg13g2_o21ai_1 _16108_ (.B1(_09598_),
    .Y(_09599_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[22] ),
    .A2(net10431));
 sg13g2_nand2b_1 _16109_ (.Y(_09600_),
    .B(_09566_),
    .A_N(_09564_));
 sg13g2_nand2b_1 _16110_ (.Y(_09601_),
    .B(_09600_),
    .A_N(_09561_));
 sg13g2_o21ai_1 _16111_ (.B1(_09601_),
    .Y(_09602_),
    .A1(net10495),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[21] ));
 sg13g2_a21oi_1 _16112_ (.A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[21] ),
    .A2(_09561_),
    .Y(_09603_),
    .B1(_09568_));
 sg13g2_nor2b_1 _16113_ (.A(_09541_),
    .B_N(_09603_),
    .Y(_09604_));
 sg13g2_o21ai_1 _16114_ (.B1(net10495),
    .Y(_09605_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[21] ),
    .A2(_09561_));
 sg13g2_o21ai_1 _16115_ (.B1(_09605_),
    .Y(_09606_),
    .A1(_09602_),
    .A2(_09604_));
 sg13g2_buf_2 place10969 (.A(net10967),
    .X(net10969));
 sg13g2_buf_2 place10958 (.A(_00005_),
    .X(net10958));
 sg13g2_buf_2 place10935 (.A(_00005_),
    .X(net10935));
 sg13g2_xor2_1 _16119_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[22] ),
    .A(net10494),
    .X(_09610_));
 sg13g2_xnor2_1 _16120_ (.Y(_09611_),
    .A(_09606_),
    .B(_09610_));
 sg13g2_buf_2 place10953 (.A(_00005_),
    .X(net10953));
 sg13g2_o21ai_1 _16122_ (.B1(net10393),
    .Y(_09613_),
    .A1(_08537_),
    .A2(net10405));
 sg13g2_a22oi_1 _16123_ (.Y(_09614_),
    .B1(net9697),
    .B2(_09613_),
    .A2(net10561),
    .A1(net10697));
 sg13g2_o21ai_1 _16124_ (.B1(_09614_),
    .Y(_09615_),
    .A1(_08395_),
    .A2(_09611_));
 sg13g2_nor2_1 _16125_ (.A(net10287),
    .B(_09615_),
    .Y(_09616_));
 sg13g2_a21oi_1 _16126_ (.A1(net10288),
    .A2(_09599_),
    .Y(_02158_),
    .B1(_09616_));
 sg13g2_buf_16 clkbuf_leaf_76_clk (.X(clknet_leaf_76_clk),
    .A(clknet_8_12_0_clk));
 sg13g2_buf_2 place10968 (.A(net10967),
    .X(net10968));
 sg13g2_nand2_1 _16129_ (.Y(_09619_),
    .A(net10649),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[55] ));
 sg13g2_buf_2 place10976 (.A(_08213_),
    .X(net10976));
 sg13g2_a22oi_1 _16131_ (.Y(_09621_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[23] ),
    .B2(net10644),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[55] ),
    .A1(net10640));
 sg13g2_nand3_1 _16132_ (.B(_09619_),
    .C(_09621_),
    .A(net10432),
    .Y(_09622_));
 sg13g2_o21ai_1 _16133_ (.B1(_09622_),
    .Y(_09623_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[23] ),
    .A2(net10431));
 sg13g2_buf_2 place10874 (.A(net10872),
    .X(net10874));
 sg13g2_buf_2 place10873 (.A(net10872),
    .X(net10873));
 sg13g2_xor2_1 _16136_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[23] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[23] ),
    .X(_09626_));
 sg13g2_nand3_1 _16137_ (.B(_09540_),
    .C(_09603_),
    .A(_09538_),
    .Y(_09627_));
 sg13g2_nand2_1 _16138_ (.Y(_09628_),
    .A(net10494),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[22] ));
 sg13g2_nand2_1 _16139_ (.Y(_09629_),
    .A(_09605_),
    .B(_09628_));
 sg13g2_nand2_1 _16140_ (.Y(_09630_),
    .A(_09605_),
    .B(_09602_));
 sg13g2_o21ai_1 _16141_ (.B1(_09630_),
    .Y(_09631_),
    .A1(net10494),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[22] ));
 sg13g2_nand2_1 _16142_ (.Y(_09632_),
    .A(_09628_),
    .B(_09631_));
 sg13g2_o21ai_1 _16143_ (.B1(_09632_),
    .Y(_09633_),
    .A1(_09627_),
    .A2(_09629_));
 sg13g2_buf_2 place10872 (.A(_00009_),
    .X(net10872));
 sg13g2_xor2_1 _16145_ (.B(_09633_),
    .A(_09626_),
    .X(_09635_));
 sg13g2_buf_2 place10906 (.A(net10905),
    .X(net10906));
 sg13g2_buf_2 place10984 (.A(net10981),
    .X(net10984));
 sg13g2_o21ai_1 _16148_ (.B1(net10393),
    .Y(_09638_),
    .A1(_08543_),
    .A2(net10405));
 sg13g2_a22oi_1 _16149_ (.Y(_09639_),
    .B1(net9697),
    .B2(_09638_),
    .A2(net10559),
    .A1(net10697));
 sg13g2_o21ai_1 _16150_ (.B1(_09639_),
    .Y(_09640_),
    .A1(_08395_),
    .A2(_09635_));
 sg13g2_nor2_1 _16151_ (.A(net10287),
    .B(_09640_),
    .Y(_09641_));
 sg13g2_a21oi_1 _16152_ (.A1(net10288),
    .A2(_09623_),
    .Y(_02159_),
    .B1(_09641_));
 sg13g2_buf_2 place10992 (.A(net10991),
    .X(net10992));
 sg13g2_buf_2 place10941 (.A(net10940),
    .X(net10941));
 sg13g2_buf_2 place10889 (.A(net10888),
    .X(net10889));
 sg13g2_buf_2 place10875 (.A(net10874),
    .X(net10875));
 sg13g2_buf_2 place10954 (.A(net10953),
    .X(net10954));
 sg13g2_buf_2 place10987 (.A(net10986),
    .X(net10987));
 sg13g2_xnor2_1 _16159_ (.Y(_09648_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[24] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[24] ));
 sg13g2_nand2_1 _16160_ (.Y(_09649_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[23] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[23] ));
 sg13g2_nor2_1 _16161_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[23] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[23] ),
    .Y(_09650_));
 sg13g2_a21oi_1 _16162_ (.A1(_09633_),
    .A2(_09649_),
    .Y(_09651_),
    .B1(_09650_));
 sg13g2_xnor2_1 _16163_ (.Y(_09652_),
    .A(_09648_),
    .B(_09651_));
 sg13g2_a21oi_2 _16164_ (.B1(_09490_),
    .Y(_09653_),
    .A2(net10399),
    .A1(_08553_));
 sg13g2_nor2b_1 _16165_ (.A(_09653_),
    .B_N(net9697),
    .Y(_09654_));
 sg13g2_a221oi_1 _16166_ (.B2(net10713),
    .C1(_09654_),
    .B1(_09652_),
    .A1(net10698),
    .Y(_09655_),
    .A2(net10556));
 sg13g2_buf_2 place10991 (.A(net10990),
    .X(net10991));
 sg13g2_nand2b_1 _16168_ (.Y(_09657_),
    .B(_09117_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.count_cycle[24] ));
 sg13g2_buf_2 place10986 (.A(net10979),
    .X(net10986));
 sg13g2_nand2_1 _16170_ (.Y(_09659_),
    .A(net10649),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[56] ));
 sg13g2_buf_2 place10989 (.A(net10979),
    .X(net10989));
 sg13g2_buf_2 place10853 (.A(net10845),
    .X(net10853));
 sg13g2_a22oi_1 _16173_ (.Y(_09662_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[24] ),
    .B2(net10644),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[56] ),
    .A1(net10640));
 sg13g2_nand3_1 _16174_ (.B(_09659_),
    .C(_09662_),
    .A(net10432),
    .Y(_09663_));
 sg13g2_a21oi_1 _16175_ (.A1(_09657_),
    .A2(_09663_),
    .Y(_09664_),
    .B1(net10284));
 sg13g2_a21oi_1 _16176_ (.A1(net10284),
    .A2(_09655_),
    .Y(_02160_),
    .B1(_09664_));
 sg13g2_buf_2 place10979 (.A(net10976),
    .X(net10979));
 sg13g2_buf_2 place10877 (.A(_00009_),
    .X(net10877));
 sg13g2_buf_2 place10852 (.A(net10850),
    .X(net10852));
 sg13g2_xor2_1 _16180_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[25] ),
    .A(net10493),
    .X(_09668_));
 sg13g2_nor2_1 _16181_ (.A(_09586_),
    .B(_09648_),
    .Y(_09669_));
 sg13g2_nand3_1 _16182_ (.B(_09626_),
    .C(_09669_),
    .A(_09610_),
    .Y(_09670_));
 sg13g2_inv_1 _16183_ (.Y(_09671_),
    .A(_09670_));
 sg13g2_nor2_1 _16184_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[24] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[24] ),
    .Y(_09672_));
 sg13g2_nor2_1 _16185_ (.A(net10494),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[22] ),
    .Y(_09673_));
 sg13g2_a22oi_1 _16186_ (.Y(_09674_),
    .B1(net10682),
    .B2(net10494),
    .A2(net10683),
    .A1(net10495));
 sg13g2_inv_2 _16187_ (.Y(_09675_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[23] ));
 sg13g2_o21ai_1 _16188_ (.B1(_09675_),
    .Y(_09676_),
    .A1(_09673_),
    .A2(_09674_));
 sg13g2_nor3_1 _16189_ (.A(_09675_),
    .B(_09673_),
    .C(_09674_),
    .Y(_09677_));
 sg13g2_a221oi_1 _16190_ (.B2(\u_ac_controller_soc_inst.u_picorv32.reg_pc[23] ),
    .C1(_09677_),
    .B1(_09676_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[24] ),
    .Y(_09678_),
    .A2(net10681));
 sg13g2_nor2_2 _16191_ (.A(_09672_),
    .B(_09678_),
    .Y(_09679_));
 sg13g2_a21oi_1 _16192_ (.A1(_09582_),
    .A2(_09671_),
    .Y(_09680_),
    .B1(_09679_));
 sg13g2_xnor2_1 _16193_ (.Y(_09681_),
    .A(_09668_),
    .B(_09680_));
 sg13g2_nand2_1 _16194_ (.Y(_09682_),
    .A(net10713),
    .B(_09681_));
 sg13g2_buf_2 place10977 (.A(net10976),
    .X(net10977));
 sg13g2_a21o_2 _16196_ (.A2(_09012_),
    .A1(net10399),
    .B1(_09490_),
    .X(_09684_));
 sg13g2_a221oi_1 _16197_ (.B2(_09684_),
    .C1(net10287),
    .B1(net9698),
    .A1(net10698),
    .Y(_09685_),
    .A2(net10553));
 sg13g2_buf_2 place10848 (.A(net10846),
    .X(net10848));
 sg13g2_nand2_1 _16199_ (.Y(_09687_),
    .A(net10649),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[57] ));
 sg13g2_a22oi_1 _16200_ (.Y(_09688_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[25] ),
    .B2(net10644),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[57] ),
    .A1(net10640));
 sg13g2_nand3_1 _16201_ (.B(_09687_),
    .C(_09688_),
    .A(net10432),
    .Y(_09689_));
 sg13g2_o21ai_1 _16202_ (.B1(_09689_),
    .Y(_09690_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[25] ),
    .A2(net10431));
 sg13g2_a22oi_1 _16203_ (.Y(_02161_),
    .B1(_09690_),
    .B2(net10288),
    .A2(_09685_),
    .A1(_09682_));
 sg13g2_buf_16 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_8_6_0_clk));
 sg13g2_buf_2 place10990 (.A(net10989),
    .X(net10990));
 sg13g2_xor2_1 _16206_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[26] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[26] ),
    .X(_09693_));
 sg13g2_nor2_1 _16207_ (.A(net10493),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[25] ),
    .Y(_09694_));
 sg13g2_nand2_1 _16208_ (.Y(_09695_),
    .A(net10493),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[25] ));
 sg13g2_nand2_1 _16209_ (.Y(_09696_),
    .A(_09650_),
    .B(_09695_));
 sg13g2_a21oi_1 _16210_ (.A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[24] ),
    .Y(_09697_),
    .B1(_09696_));
 sg13g2_a21oi_1 _16211_ (.A1(_09672_),
    .A2(_09695_),
    .Y(_09698_),
    .B1(_09697_));
 sg13g2_nand2_1 _16212_ (.Y(_09699_),
    .A(_09649_),
    .B(_09695_));
 sg13g2_nor2_1 _16213_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[24] ),
    .B(_09699_),
    .Y(_09700_));
 sg13g2_nor2_1 _16214_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[24] ),
    .B(_09699_),
    .Y(_09701_));
 sg13g2_o21ai_1 _16215_ (.B1(_09633_),
    .Y(_09702_),
    .A1(_09700_),
    .A2(_09701_));
 sg13g2_nand3b_1 _16216_ (.B(_09698_),
    .C(_09702_),
    .Y(_09703_),
    .A_N(_09694_));
 sg13g2_xnor2_1 _16217_ (.Y(_09704_),
    .A(_09693_),
    .B(_09703_));
 sg13g2_nand2_1 _16218_ (.Y(_09705_),
    .A(net10713),
    .B(_09704_));
 sg13g2_buf_2 place10981 (.A(net10980),
    .X(net10981));
 sg13g2_buf_2 place10980 (.A(net10979),
    .X(net10980));
 sg13g2_buf_2 place10867 (.A(net10866),
    .X(net10867));
 sg13g2_o21ai_1 _16222_ (.B1(_09453_),
    .Y(_09709_),
    .A1(net10404),
    .A2(_09042_));
 sg13g2_a221oi_1 _16223_ (.B2(_09709_),
    .C1(net10287),
    .B1(net9698),
    .A1(net10698),
    .Y(_09710_),
    .A2(net10550));
 sg13g2_buf_2 place10850 (.A(net10846),
    .X(net10850));
 sg13g2_nand2_1 _16225_ (.Y(_09712_),
    .A(net10649),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[58] ));
 sg13g2_buf_2 place10849 (.A(net10846),
    .X(net10849));
 sg13g2_buf_2 place10985 (.A(net10984),
    .X(net10985));
 sg13g2_a22oi_1 _16228_ (.Y(_09715_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[26] ),
    .B2(net10644),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[58] ),
    .A1(net10640));
 sg13g2_nand3_1 _16229_ (.B(_09712_),
    .C(_09715_),
    .A(net10432),
    .Y(_09716_));
 sg13g2_o21ai_1 _16230_ (.B1(_09716_),
    .Y(_09717_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[26] ),
    .A2(net10431));
 sg13g2_a22oi_1 _16231_ (.Y(_02162_),
    .B1(_09717_),
    .B2(net10288),
    .A2(_09710_),
    .A1(_09705_));
 sg13g2_buf_2 place10793 (.A(net10784),
    .X(net10793));
 sg13g2_nand2_1 _16233_ (.Y(_09719_),
    .A(net10649),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[59] ));
 sg13g2_a22oi_1 _16234_ (.Y(_09720_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[27] ),
    .B2(net10644),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[59] ),
    .A1(net10640));
 sg13g2_nand3_1 _16235_ (.B(_09719_),
    .C(_09720_),
    .A(net10432),
    .Y(_09721_));
 sg13g2_o21ai_1 _16236_ (.B1(_09721_),
    .Y(_09722_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[27] ),
    .A2(net10431));
 sg13g2_buf_2 place10791 (.A(net10790),
    .X(net10791));
 sg13g2_buf_2 place10876 (.A(_00009_),
    .X(net10876));
 sg13g2_buf_2 place10965 (.A(net10964),
    .X(net10965));
 sg13g2_xor2_1 _16240_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[27] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[27] ),
    .X(_09726_));
 sg13g2_nor2_1 _16241_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[26] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[26] ),
    .Y(_09727_));
 sg13g2_nor2_1 _16242_ (.A(_09726_),
    .B(_09727_),
    .Y(_09728_));
 sg13g2_nand2_2 _16243_ (.Y(_09729_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[26] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[26] ));
 sg13g2_and2_1 _16244_ (.A(_09726_),
    .B(_09729_),
    .X(_09730_));
 sg13g2_mux2_1 _16245_ (.A0(_09728_),
    .A1(_09730_),
    .S(_09703_),
    .X(_09731_));
 sg13g2_nand2_1 _16246_ (.Y(_09732_),
    .A(_09726_),
    .B(_09727_));
 sg13g2_o21ai_1 _16247_ (.B1(_09732_),
    .Y(_09733_),
    .A1(_09726_),
    .A2(_09729_));
 sg13g2_o21ai_1 _16248_ (.B1(net10713),
    .Y(_09734_),
    .A1(_09731_),
    .A2(_09733_));
 sg13g2_buf_2 place10964 (.A(net10958),
    .X(net10964));
 sg13g2_o21ai_1 _16250_ (.B1(_09453_),
    .Y(_09736_),
    .A1(net10404),
    .A2(_09074_));
 sg13g2_a221oi_1 _16251_ (.B2(_09736_),
    .C1(net10287),
    .B1(net9698),
    .A1(net10698),
    .Y(_09737_),
    .A2(net10547));
 sg13g2_a22oi_1 _16252_ (.Y(_02163_),
    .B1(_09734_),
    .B2(_09737_),
    .A2(_09722_),
    .A1(net10288));
 sg13g2_nor2_1 _16253_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[27] ),
    .B(net10678),
    .Y(_09738_));
 sg13g2_nor2_1 _16254_ (.A(_09694_),
    .B(_09738_),
    .Y(_09739_));
 sg13g2_nand4_1 _16255_ (.B(_09702_),
    .C(_09698_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[26] ),
    .Y(_09740_),
    .D(_09739_));
 sg13g2_nand4_1 _16256_ (.B(_09702_),
    .C(_09698_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[26] ),
    .Y(_09741_),
    .D(_09739_));
 sg13g2_nor2_1 _16257_ (.A(_09729_),
    .B(_09738_),
    .Y(_09742_));
 sg13g2_a21oi_1 _16258_ (.A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[27] ),
    .Y(_09743_),
    .B1(_09742_));
 sg13g2_nand3_1 _16259_ (.B(_09741_),
    .C(_09743_),
    .A(_09740_),
    .Y(_09744_));
 sg13g2_buf_2 place10851 (.A(net10850),
    .X(net10851));
 sg13g2_buf_2 place10956 (.A(net10954),
    .X(net10956));
 sg13g2_buf_2 place10788 (.A(net10787),
    .X(net10788));
 sg13g2_xor2_1 _16263_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[28] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[28] ),
    .X(_09748_));
 sg13g2_xnor2_1 _16264_ (.Y(_09749_),
    .A(_09744_),
    .B(_09748_));
 sg13g2_buf_2 place10786 (.A(net10784),
    .X(net10786));
 sg13g2_buf_2 place10790 (.A(net10789),
    .X(net10790));
 sg13g2_o21ai_1 _16267_ (.B1(net10393),
    .Y(_09752_),
    .A1(net10405),
    .A2(_09106_));
 sg13g2_buf_2 place10789 (.A(net10787),
    .X(net10789));
 sg13g2_buf_2 place10787 (.A(net10786),
    .X(net10787));
 sg13g2_a22oi_1 _16270_ (.Y(_09755_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[60] ),
    .B2(net10647),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[28] ),
    .A1(net10644));
 sg13g2_inv_1 _16271_ (.Y(_09756_),
    .A(_09755_));
 sg13g2_a221oi_1 _16272_ (.B2(_09117_),
    .C1(_09756_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh ),
    .Y(_09757_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[60] ));
 sg13g2_nor2_1 _16273_ (.A(net10284),
    .B(_09757_),
    .Y(_09758_));
 sg13g2_a221oi_1 _16274_ (.B2(_09752_),
    .C1(_09758_),
    .B1(net9698),
    .A1(net10698),
    .Y(_09759_),
    .A2(net10545));
 sg13g2_o21ai_1 _16275_ (.B1(_09759_),
    .Y(_02164_),
    .A1(_09376_),
    .A2(_09749_));
 sg13g2_buf_16 clkbuf_leaf_59_clk (.X(clknet_leaf_59_clk),
    .A(clknet_8_1_0_clk));
 sg13g2_buf_2 place10776 (.A(net10775),
    .X(net10776));
 sg13g2_buf_2 place10777 (.A(net10775),
    .X(net10777));
 sg13g2_xnor2_1 _16279_ (.Y(_09763_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[29] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[29] ));
 sg13g2_a21o_1 _16280_ (.A2(_09679_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[25] ),
    .B1(net10493),
    .X(_09764_));
 sg13g2_o21ai_1 _16281_ (.B1(_09764_),
    .Y(_09765_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[25] ),
    .A2(_09679_));
 sg13g2_o21ai_1 _16282_ (.B1(_09729_),
    .Y(_09766_),
    .A1(_09727_),
    .A2(_09765_));
 sg13g2_a21oi_1 _16283_ (.A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[27] ),
    .A2(_09766_),
    .Y(_09767_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[27] ));
 sg13g2_nor2_1 _16284_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[27] ),
    .B(_09766_),
    .Y(_09768_));
 sg13g2_nand2_1 _16285_ (.Y(_09769_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[28] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[28] ));
 sg13g2_o21ai_1 _16286_ (.B1(_09769_),
    .Y(_09770_),
    .A1(_09767_),
    .A2(_09768_));
 sg13g2_nand3_1 _16287_ (.B(_09693_),
    .C(_09726_),
    .A(_09668_),
    .Y(_09771_));
 sg13g2_nor4_2 _16288_ (.A(_09564_),
    .B(_09581_),
    .C(_09670_),
    .Y(_09772_),
    .D(_09771_));
 sg13g2_or2_1 _16289_ (.X(_09773_),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[28] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[28] ));
 sg13g2_o21ai_1 _16290_ (.B1(_09773_),
    .Y(_09774_),
    .A1(_09770_),
    .A2(_09772_));
 sg13g2_xnor2_1 _16291_ (.Y(_09775_),
    .A(_09763_),
    .B(_09774_));
 sg13g2_buf_2 place10773 (.A(net10772),
    .X(net10773));
 sg13g2_buf_2 place10797 (.A(net10796),
    .X(net10797));
 sg13g2_o21ai_1 _16294_ (.B1(_09453_),
    .Y(_09778_),
    .A1(net10404),
    .A2(_09147_));
 sg13g2_buf_2 place11009 (.A(net11008),
    .X(net11009));
 sg13g2_buf_2 place10897 (.A(net10894),
    .X(net10897));
 sg13g2_buf_2 place10884 (.A(_00007_),
    .X(net10884));
 sg13g2_a22oi_1 _16298_ (.Y(_09782_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[61] ),
    .B2(net10648),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[29] ),
    .A1(net10643));
 sg13g2_inv_1 _16299_ (.Y(_09783_),
    .A(_09782_));
 sg13g2_a221oi_1 _16300_ (.B2(_09117_),
    .C1(_09783_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh ),
    .Y(_09784_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[61] ));
 sg13g2_nor2_1 _16301_ (.A(net10284),
    .B(_09784_),
    .Y(_09785_));
 sg13g2_a221oi_1 _16302_ (.B2(_09778_),
    .C1(_09785_),
    .B1(net9698),
    .A1(net10698),
    .Y(_09786_),
    .A2(net10543));
 sg13g2_o21ai_1 _16303_ (.B1(_09786_),
    .Y(_02165_),
    .A1(_09376_),
    .A2(_09775_));
 sg13g2_or2_1 _16304_ (.X(_09787_),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[29] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[29] ));
 sg13g2_and2_1 _16305_ (.A(_09773_),
    .B(_09787_),
    .X(_09788_));
 sg13g2_o21ai_1 _16306_ (.B1(_09788_),
    .Y(_09789_),
    .A1(_09770_),
    .A2(_09772_));
 sg13g2_nand2_1 _16307_ (.Y(_09790_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[29] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[29] ));
 sg13g2_nand2_1 _16308_ (.Y(_09791_),
    .A(_09789_),
    .B(_09790_));
 sg13g2_buf_2 place10902 (.A(net10901),
    .X(net10902));
 sg13g2_buf_2 place10866 (.A(net10861),
    .X(net10866));
 sg13g2_xor2_1 _16311_ (.B(net10674),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[30] ),
    .X(_09794_));
 sg13g2_xnor2_1 _16312_ (.Y(_09795_),
    .A(_09791_),
    .B(_09794_));
 sg13g2_buf_2 place10758 (.A(net10755),
    .X(net10758));
 sg13g2_buf_2 place10784 (.A(_00001_),
    .X(net10784));
 sg13g2_o21ai_1 _16315_ (.B1(_09453_),
    .Y(_09798_),
    .A1(net10404),
    .A2(_09178_));
 sg13g2_buf_2 place10883 (.A(_00007_),
    .X(net10883));
 sg13g2_buf_2 place10885 (.A(net10884),
    .X(net10885));
 sg13g2_a22oi_1 _16318_ (.Y(_09801_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[62] ),
    .B2(net10648),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[30] ),
    .A1(net10643));
 sg13g2_inv_1 _16319_ (.Y(_09802_),
    .A(_09801_));
 sg13g2_a221oi_1 _16320_ (.B2(_09117_),
    .C1(_09802_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh ),
    .Y(_09803_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[62] ));
 sg13g2_nor2_1 _16321_ (.A(net10284),
    .B(_09803_),
    .Y(_09804_));
 sg13g2_a221oi_1 _16322_ (.B2(_09798_),
    .C1(_09804_),
    .B1(net9698),
    .A1(net10698),
    .Y(_09805_),
    .A2(net10537));
 sg13g2_o21ai_1 _16323_ (.B1(_09805_),
    .Y(_02167_),
    .A1(_09376_),
    .A2(_09795_));
 sg13g2_buf_2 place10870 (.A(net10869),
    .X(net10870));
 sg13g2_nand2_1 _16325_ (.Y(_09807_),
    .A(net10648),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[63] ));
 sg13g2_a22oi_1 _16326_ (.Y(_09808_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.count_instr[31] ),
    .B2(net10643),
    .A2(\u_ac_controller_soc_inst.u_picorv32.count_instr[63] ),
    .A1(net10640));
 sg13g2_nand3_1 _16327_ (.B(_09807_),
    .C(_09808_),
    .A(_08320_),
    .Y(_09809_));
 sg13g2_o21ai_1 _16328_ (.B1(_09809_),
    .Y(_09810_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[31] ),
    .A2(_08320_));
 sg13g2_nand2_1 _16329_ (.Y(_09811_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[30] ),
    .B(net10674));
 sg13g2_buf_2 place10892 (.A(net10884),
    .X(net10892));
 sg13g2_buf_2 place10898 (.A(net10897),
    .X(net10898));
 sg13g2_xor2_1 _16332_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[31] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[31] ),
    .X(_09814_));
 sg13g2_nor2_1 _16333_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[30] ),
    .B(net10674),
    .Y(_09815_));
 sg13g2_nand2_1 _16334_ (.Y(_09816_),
    .A(_09814_),
    .B(_09815_));
 sg13g2_o21ai_1 _16335_ (.B1(_09816_),
    .Y(_09817_),
    .A1(_09811_),
    .A2(_09814_));
 sg13g2_a21o_2 _16336_ (.A2(_09208_),
    .A1(net10399),
    .B1(_09490_),
    .X(_09818_));
 sg13g2_inv_16 _16337_ (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[4] ),
    .Y(_09819_));
 sg13g2_o21ai_1 _16338_ (.B1(net10284),
    .Y(_09820_),
    .A1(_09819_),
    .A2(_08586_));
 sg13g2_a221oi_1 _16339_ (.B2(net9698),
    .C1(_09820_),
    .B1(_09818_),
    .A1(net10713),
    .Y(_09821_),
    .A2(_09817_));
 sg13g2_or2_1 _16340_ (.X(_09822_),
    .B(_09815_),
    .A(_09814_));
 sg13g2_a21oi_1 _16341_ (.A1(_09789_),
    .A2(_09790_),
    .Y(_09823_),
    .B1(_09822_));
 sg13g2_and4_1 _16342_ (.A(_09789_),
    .B(_09790_),
    .C(_09811_),
    .D(_09814_),
    .X(_09824_));
 sg13g2_o21ai_1 _16343_ (.B1(net10713),
    .Y(_09825_),
    .A1(_09823_),
    .A2(_09824_));
 sg13g2_a22oi_1 _16344_ (.Y(_02168_),
    .B1(_09821_),
    .B2(_09825_),
    .A2(_09810_),
    .A1(net10287));
 sg13g2_buf_16 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_8_54_0_clk));
 sg13g2_buf_2 place10887 (.A(net10886),
    .X(net10887));
 sg13g2_buf_2 place10782 (.A(_00002_),
    .X(net10782));
 sg13g2_buf_2 place10871 (.A(net10869),
    .X(net10871));
 sg13g2_buf_2 place10868 (.A(net10867),
    .X(net10868));
 sg13g2_buf_2 place11001 (.A(net11000),
    .X(net11001));
 sg13g2_buf_2 place11010 (.A(net11009),
    .X(net11010));
 sg13g2_buf_2 place10785 (.A(net10784),
    .X(net10785));
 sg13g2_buf_2 place10775 (.A(_00002_),
    .X(net10775));
 sg13g2_buf_2 place10960 (.A(net10958),
    .X(net10960));
 sg13g2_buf_2 place10735 (.A(_00103_),
    .X(net10735));
 sg13g2_buf_2 place10847 (.A(net10846),
    .X(net10847));
 sg13g2_buf_2 place10770 (.A(_00003_),
    .X(net10770));
 sg13g2_buf_2 place10907 (.A(net10906),
    .X(net10907));
 sg13g2_buf_2 place10865 (.A(net10861),
    .X(net10865));
 sg13g2_buf_2 place10961 (.A(net10960),
    .X(net10961));
 sg13g2_buf_2 place10963 (.A(net10962),
    .X(net10963));
 sg13g2_buf_2 place10772 (.A(net10771),
    .X(net10772));
 sg13g2_buf_2 place10771 (.A(_00003_),
    .X(net10771));
 sg13g2_buf_2 place10765 (.A(net10764),
    .X(net10765));
 sg13g2_buf_2 place10792 (.A(net10786),
    .X(net10792));
 sg13g2_buf_2 place10905 (.A(net10904),
    .X(net10905));
 sg13g2_buf_2 place10795 (.A(net10793),
    .X(net10795));
 sg13g2_buf_2 place10959 (.A(net10958),
    .X(net10959));
 sg13g2_buf_2 place10967 (.A(net10965),
    .X(net10967));
 sg13g2_buf_2 place10857 (.A(net10845),
    .X(net10857));
 sg13g2_buf_2 place10862 (.A(net10861),
    .X(net10862));
 sg13g2_buf_2 place10766 (.A(net10765),
    .X(net10766));
 sg13g2_buf_2 place10767 (.A(net10765),
    .X(net10767));
 sg13g2_buf_2 place10783 (.A(net10782),
    .X(net10783));
 sg13g2_buf_2 place10794 (.A(net10793),
    .X(net10794));
 sg13g2_buf_2 place10860 (.A(net10859),
    .X(net10860));
 sg13g2_buf_2 place10760 (.A(net10759),
    .X(net10760));
 sg13g2_buf_2 place10796 (.A(net10795),
    .X(net10796));
 sg13g2_buf_2 place10803 (.A(net10799),
    .X(net10803));
 sg13g2_nor2b_2 _16380_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_branch ),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.latched_store ),
    .Y(_09828_));
 sg13g2_buf_2 place10750 (.A(net10748),
    .X(net10750));
 sg13g2_buf_2 place10709 (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[3] ),
    .X(net10709));
 sg13g2_buf_2 place10698 (.A(net10697),
    .X(net10698));
 sg13g2_buf_2 place10695 (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[6] ),
    .X(net10695));
 sg13g2_buf_2 place10696 (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[6] ),
    .X(net10696));
 sg13g2_buf_2 place10846 (.A(net10845),
    .X(net10846));
 sg13g2_mux2_1 _16387_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[0] ),
    .S(\u_ac_controller_soc_inst.u_picorv32.latched_stalu ),
    .X(_09835_));
 sg13g2_nand2_2 _16388_ (.Y(_09836_),
    .A(net10384),
    .B(_09835_));
 sg13g2_buf_2 place10693 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[11] ),
    .X(net10693));
 sg13g2_buf_2 place10692 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[12] ),
    .X(net10692));
 sg13g2_buf_2 place10691 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[13] ),
    .X(net10691));
 sg13g2_buf_2 place10903 (.A(net10902),
    .X(net10903));
 sg13g2_buf_2 place10690 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[15] ),
    .X(net10690));
 sg13g2_nand2b_2 _16394_ (.Y(_09842_),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_rd[3] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.latched_rd[4] ));
 sg13g2_nor2_2 _16395_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[2] ),
    .B(_09842_),
    .Y(_09843_));
 sg13g2_buf_2 place10904 (.A(net10893),
    .X(net10904));
 sg13g2_inv_1 _16397_ (.Y(_09845_),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[1] ));
 sg13g2_buf_2 place10734 (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[0] ),
    .X(net10734));
 sg13g2_inv_8 _16399_ (.Y(_09847_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[1] ));
 sg13g2_nor2_2 _16400_ (.A(net11019),
    .B(_09847_),
    .Y(_09848_));
 sg13g2_o21ai_1 _16401_ (.B1(_09848_),
    .Y(_09849_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.latched_store ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.latched_branch ));
 sg13g2_nor3_2 _16402_ (.A(_09845_),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_rd[0] ),
    .C(_09849_),
    .Y(_09850_));
 sg13g2_buf_2 place10689 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[16] ),
    .X(net10689));
 sg13g2_nand2_2 _16404_ (.Y(_09852_),
    .A(_09843_),
    .B(_09850_));
 sg13g2_buf_2 place10688 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[17] ),
    .X(net10688));
 sg13g2_buf_2 place10741 (.A(_00103_),
    .X(net10741));
 sg13g2_buf_2 place10753 (.A(net10752),
    .X(net10753));
 sg13g2_nand2_1 _16408_ (.Y(_09856_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][0] ),
    .B(net10135));
 sg13g2_o21ai_1 _16409_ (.B1(_09856_),
    .Y(_00690_),
    .A1(net10276),
    .A2(net10135));
 sg13g2_nand2b_2 _16410_ (.Y(_09857_),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_store ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.latched_branch ));
 sg13g2_buf_2 place10726 (.A(net10725),
    .X(net10726));
 sg13g2_buf_2 place10755 (.A(net10752),
    .X(net10755));
 sg13g2_mux2_1 _16413_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[10] ),
    .S(net10630),
    .X(_09860_));
 sg13g2_inv_2 _16414_ (.Y(_09861_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[7] ));
 sg13g2_nand4_1 _16415_ (.B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[2] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.reg_pc[4] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[3] ),
    .Y(_09862_),
    .D(\u_ac_controller_soc_inst.u_picorv32.reg_pc[5] ));
 sg13g2_buf_2 place10694 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[10] ),
    .X(net10694));
 sg13g2_nand2_1 _16417_ (.Y(_09864_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[8] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[9] ));
 sg13g2_nor4_2 _16418_ (.A(_09285_),
    .B(_09861_),
    .C(_09862_),
    .Y(_09865_),
    .D(_09864_));
 sg13g2_xnor2_1 _16419_ (.Y(_09866_),
    .A(net10498),
    .B(_09865_));
 sg13g2_nand2_1 _16420_ (.Y(_09867_),
    .A(_09857_),
    .B(_09866_));
 sg13g2_o21ai_1 _16421_ (.B1(_09867_),
    .Y(_09868_),
    .A1(_09857_),
    .A2(_09860_));
 sg13g2_buf_2 place10699 (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[4] ),
    .X(net10699));
 sg13g2_buf_2 place10802 (.A(net10801),
    .X(net10802));
 sg13g2_nand2_1 _16424_ (.Y(_09871_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][10] ),
    .B(net10138));
 sg13g2_o21ai_1 _16425_ (.B1(_09871_),
    .Y(_00691_),
    .A1(net10138),
    .A2(net10131));
 sg13g2_mux2_1 _16426_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[11] ),
    .S(net10630),
    .X(_09872_));
 sg13g2_buf_2 place10683 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[21] ),
    .X(net10683));
 sg13g2_and2_1 _16428_ (.A(net10498),
    .B(_09865_),
    .X(_09874_));
 sg13g2_xnor2_1 _16429_ (.Y(_09875_),
    .A(net10497),
    .B(_09874_));
 sg13g2_nor2_1 _16430_ (.A(_09828_),
    .B(_09875_),
    .Y(_09876_));
 sg13g2_a21oi_2 _16431_ (.B1(_09876_),
    .Y(_09877_),
    .A2(_09872_),
    .A1(net10384));
 sg13g2_buf_2 place10859 (.A(net10858),
    .X(net10859));
 sg13g2_buf_2 place10682 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[22] ),
    .X(net10682));
 sg13g2_nand2_1 _16434_ (.Y(_09880_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][11] ),
    .B(net10141));
 sg13g2_o21ai_1 _16435_ (.B1(_09880_),
    .Y(_00692_),
    .A1(net10141),
    .A2(net9985));
 sg13g2_mux2_1 _16436_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[12] ),
    .S(net10630),
    .X(_09881_));
 sg13g2_nand2_1 _16437_ (.Y(_09882_),
    .A(net10497),
    .B(_09874_));
 sg13g2_xor2_1 _16438_ (.B(_09882_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[12] ),
    .X(_09883_));
 sg13g2_nor2_1 _16439_ (.A(net10385),
    .B(_09883_),
    .Y(_09884_));
 sg13g2_a21oi_2 _16440_ (.B1(_09884_),
    .Y(_09885_),
    .A2(_09881_),
    .A1(net10385));
 sg13g2_buf_2 place10681 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[24] ),
    .X(net10681));
 sg13g2_buf_2 place10687 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[18] ),
    .X(net10687));
 sg13g2_nand2_1 _16443_ (.Y(_09888_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][12] ),
    .B(net10136));
 sg13g2_o21ai_1 _16444_ (.B1(_09888_),
    .Y(_00693_),
    .A1(net10136),
    .A2(net9801));
 sg13g2_mux2_1 _16445_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[13] ),
    .S(\u_ac_controller_soc_inst.u_picorv32.latched_stalu ),
    .X(_09889_));
 sg13g2_and4_2 _16446_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[10] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[11] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.reg_pc[12] ),
    .D(_09865_),
    .X(_09890_));
 sg13g2_buf_2 place10779 (.A(net10778),
    .X(net10779));
 sg13g2_xnor2_1 _16448_ (.Y(_09892_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[13] ),
    .B(_09890_));
 sg13g2_nor2_1 _16449_ (.A(net10384),
    .B(_09892_),
    .Y(_09893_));
 sg13g2_a21oi_2 _16450_ (.B1(_09893_),
    .Y(_09894_),
    .A2(_09889_),
    .A1(net10384));
 sg13g2_buf_2 place10686 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[19] ),
    .X(net10686));
 sg13g2_buf_2 place10679 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[26] ),
    .X(net10679));
 sg13g2_nand2_1 _16453_ (.Y(_09897_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][13] ),
    .B(net10135));
 sg13g2_o21ai_1 _16454_ (.B1(_09897_),
    .Y(_00694_),
    .A1(net10135),
    .A2(net9981));
 sg13g2_mux2_1 _16455_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[14] ),
    .S(\u_ac_controller_soc_inst.u_picorv32.latched_stalu ),
    .X(_09898_));
 sg13g2_nand2_1 _16456_ (.Y(_09899_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[13] ),
    .B(_09890_));
 sg13g2_xor2_1 _16457_ (.B(_09899_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[14] ),
    .X(_09900_));
 sg13g2_nor2_1 _16458_ (.A(net10388),
    .B(_09900_),
    .Y(_09901_));
 sg13g2_a21oi_2 _16459_ (.B1(_09901_),
    .Y(_09902_),
    .A2(_09898_),
    .A1(net10388));
 sg13g2_buf_2 place10678 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[27] ),
    .X(net10678));
 sg13g2_buf_2 place10778 (.A(_00002_),
    .X(net10778));
 sg13g2_nand2_1 _16462_ (.Y(_09905_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][14] ),
    .B(_09852_));
 sg13g2_o21ai_1 _16463_ (.B1(_09905_),
    .Y(_00695_),
    .A1(_09852_),
    .A2(net9796));
 sg13g2_mux2_1 _16464_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[15] ),
    .S(net10627),
    .X(_09906_));
 sg13g2_and3_2 _16465_ (.X(_09907_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[13] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[14] ),
    .C(_09890_));
 sg13g2_buf_2 place10677 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[28] ),
    .X(net10677));
 sg13g2_xnor2_1 _16467_ (.Y(_09909_),
    .A(net10496),
    .B(_09907_));
 sg13g2_nor2_1 _16468_ (.A(net10388),
    .B(_09909_),
    .Y(_09910_));
 sg13g2_a21oi_2 _16469_ (.B1(_09910_),
    .Y(_09911_),
    .A2(_09906_),
    .A1(net10388));
 sg13g2_buf_2 place10781 (.A(net10778),
    .X(net10781));
 sg13g2_buf_2 place10676 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[29] ),
    .X(net10676));
 sg13g2_nand2_1 _16472_ (.Y(_09914_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][15] ),
    .B(net10138));
 sg13g2_o21ai_1 _16473_ (.B1(_09914_),
    .Y(_00696_),
    .A1(net10138),
    .A2(net9792));
 sg13g2_mux2_1 _16474_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[16] ),
    .S(net10627),
    .X(_09915_));
 sg13g2_nand2_1 _16475_ (.Y(_09916_),
    .A(net10496),
    .B(_09907_));
 sg13g2_xor2_1 _16476_ (.B(_09916_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[16] ),
    .X(_09917_));
 sg13g2_nor2_1 _16477_ (.A(net10388),
    .B(_09917_),
    .Y(_09918_));
 sg13g2_a21oi_2 _16478_ (.B1(_09918_),
    .Y(_09919_),
    .A2(_09915_),
    .A1(net10388));
 sg13g2_buf_2 place10680 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[25] ),
    .X(net10680));
 sg13g2_buf_2 place10675 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[2] ),
    .X(net10675));
 sg13g2_nand2_1 _16481_ (.Y(_09922_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][16] ),
    .B(net10138));
 sg13g2_o21ai_1 _16482_ (.B1(_09922_),
    .Y(_00697_),
    .A1(net10138),
    .A2(net9745));
 sg13g2_mux2_1 _16483_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[17] ),
    .S(net10627),
    .X(_09923_));
 sg13g2_buf_2 place10742 (.A(net10741),
    .X(net10742));
 sg13g2_nand3_1 _16485_ (.B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[16] ),
    .C(_09907_),
    .A(net10496),
    .Y(_09925_));
 sg13g2_xor2_1 _16486_ (.B(_09925_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[17] ),
    .X(_09926_));
 sg13g2_nor2_1 _16487_ (.A(net10388),
    .B(_09926_),
    .Y(_09927_));
 sg13g2_a21oi_2 _16488_ (.B1(_09927_),
    .Y(_09928_),
    .A2(_09923_),
    .A1(net10388));
 sg13g2_buf_2 place10685 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[20] ),
    .X(net10685));
 sg13g2_buf_2 place10780 (.A(net10779),
    .X(net10780));
 sg13g2_buf_2 place10774 (.A(net10771),
    .X(net10774));
 sg13g2_nand2_1 _16492_ (.Y(_09932_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][17] ),
    .B(net10137));
 sg13g2_o21ai_1 _16493_ (.B1(_09932_),
    .Y(_00698_),
    .A1(net10137),
    .A2(net9742));
 sg13g2_mux2_1 _16494_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[18] ),
    .S(net10627),
    .X(_09933_));
 sg13g2_and4_2 _16495_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[15] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[16] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.reg_pc[17] ),
    .D(_09907_),
    .X(_09934_));
 sg13g2_buf_2 place10684 (.A(net10683),
    .X(net10684));
 sg13g2_xnor2_1 _16497_ (.Y(_09936_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[18] ),
    .B(_09934_));
 sg13g2_nor2_1 _16498_ (.A(net10387),
    .B(_09936_),
    .Y(_09937_));
 sg13g2_a21oi_2 _16499_ (.B1(_09937_),
    .Y(_09938_),
    .A2(_09933_),
    .A1(net10387));
 sg13g2_buf_2 place11011 (.A(net11010),
    .X(net11011));
 sg13g2_buf_2 place10894 (.A(net10893),
    .X(net10894));
 sg13g2_nand2_1 _16502_ (.Y(_09941_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][18] ),
    .B(net10140));
 sg13g2_o21ai_1 _16503_ (.B1(_09941_),
    .Y(_00699_),
    .A1(net10140),
    .A2(net9735));
 sg13g2_buf_2 place11005 (.A(net11004),
    .X(net11005));
 sg13g2_mux2_1 _16505_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[19] ),
    .S(net10627),
    .X(_09943_));
 sg13g2_nand2_1 _16506_ (.Y(_09944_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[18] ),
    .B(_09934_));
 sg13g2_xor2_1 _16507_ (.B(_09944_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[19] ),
    .X(_09945_));
 sg13g2_nor2_1 _16508_ (.A(net10390),
    .B(_09945_),
    .Y(_09946_));
 sg13g2_a21oi_2 _16509_ (.B1(_09946_),
    .Y(_09947_),
    .A2(_09943_),
    .A1(net10390));
 sg13g2_buf_2 place10671 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[5] ),
    .X(net10671));
 sg13g2_buf_2 place10759 (.A(net10758),
    .X(net10759));
 sg13g2_nand2_1 _16512_ (.Y(_09950_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][19] ),
    .B(net10143));
 sg13g2_o21ai_1 _16513_ (.B1(_09950_),
    .Y(_00700_),
    .A1(net10143),
    .A2(net9724));
 sg13g2_buf_2 place11002 (.A(net10990),
    .X(net11002));
 sg13g2_mux2_1 _16515_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[1] ),
    .S(net10631),
    .X(_09952_));
 sg13g2_and2_1 _16516_ (.A(net10385),
    .B(_09952_),
    .X(_09953_));
 sg13g2_a21oi_2 _16517_ (.B1(_09953_),
    .Y(_09954_),
    .A2(_09857_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[1] ));
 sg13g2_buf_2 place10670 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[6] ),
    .X(net10670));
 sg13g2_buf_2 place10858 (.A(net10857),
    .X(net10858));
 sg13g2_nand2_1 _16520_ (.Y(_09957_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][1] ),
    .B(net10134));
 sg13g2_o21ai_1 _16521_ (.B1(_09957_),
    .Y(_00701_),
    .A1(net10137),
    .A2(net10228));
 sg13g2_buf_2 place10674 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[30] ),
    .X(net10674));
 sg13g2_mux2_1 _16523_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[20] ),
    .S(net10628),
    .X(_09959_));
 sg13g2_nand3_1 _16524_ (.B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[19] ),
    .C(_09934_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[18] ),
    .Y(_09960_));
 sg13g2_xor2_1 _16525_ (.B(_09960_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[20] ),
    .X(_09961_));
 sg13g2_nor2_1 _16526_ (.A(net10389),
    .B(_09961_),
    .Y(_09962_));
 sg13g2_a21oi_2 _16527_ (.B1(_09962_),
    .Y(_09963_),
    .A2(_09959_),
    .A1(net10387));
 sg13g2_buf_2 place10743 (.A(net10742),
    .X(net10743));
 sg13g2_buf_16 clkbuf_leaf_140_clk (.X(clknet_leaf_140_clk),
    .A(clknet_8_28_0_clk));
 sg13g2_nand2_1 _16530_ (.Y(_09966_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][20] ),
    .B(net10139));
 sg13g2_o21ai_1 _16531_ (.B1(_09966_),
    .Y(_00702_),
    .A1(net10139),
    .A2(net9719));
 sg13g2_mux2_1 _16532_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[21] ),
    .S(net10628),
    .X(_09967_));
 sg13g2_and4_2 _16533_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[18] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[19] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.reg_pc[20] ),
    .D(_09934_),
    .X(_09968_));
 sg13g2_buf_2 place10673 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[3] ),
    .X(net10673));
 sg13g2_xnor2_1 _16535_ (.Y(_09970_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[21] ),
    .B(_09968_));
 sg13g2_nor2_1 _16536_ (.A(net10389),
    .B(_09970_),
    .Y(_09971_));
 sg13g2_a21oi_2 _16537_ (.B1(_09971_),
    .Y(_09972_),
    .A2(_09967_),
    .A1(net10389));
 sg13g2_buf_2 place11008 (.A(net11007),
    .X(net11008));
 sg13g2_buf_2 place10746 (.A(net10745),
    .X(net10746));
 sg13g2_nand2_1 _16540_ (.Y(_09975_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][21] ),
    .B(net10139));
 sg13g2_o21ai_1 _16541_ (.B1(_09975_),
    .Y(_00703_),
    .A1(net10139),
    .A2(net9714));
 sg13g2_mux2_1 _16542_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[22] ),
    .S(net10629),
    .X(_09976_));
 sg13g2_nand2_1 _16543_ (.Y(_09977_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[21] ),
    .B(_09968_));
 sg13g2_xor2_1 _16544_ (.B(_09977_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[22] ),
    .X(_09978_));
 sg13g2_nor2_1 _16545_ (.A(net10389),
    .B(_09978_),
    .Y(_09979_));
 sg13g2_a21oi_2 _16546_ (.B1(_09979_),
    .Y(_09980_),
    .A2(_09976_),
    .A1(net10389));
 sg13g2_buf_2 place11007 (.A(net11006),
    .X(net11007));
 sg13g2_buf_2 place11006 (.A(net11005),
    .X(net11006));
 sg13g2_nand2_1 _16549_ (.Y(_09983_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][22] ),
    .B(net10140));
 sg13g2_o21ai_1 _16550_ (.B1(_09983_),
    .Y(_00704_),
    .A1(net10140),
    .A2(net9696));
 sg13g2_mux2_1 _16551_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[23] ),
    .S(net10629),
    .X(_09984_));
 sg13g2_nand3_1 _16552_ (.B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[22] ),
    .C(_09968_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[21] ),
    .Y(_09985_));
 sg13g2_xor2_1 _16553_ (.B(_09985_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[23] ),
    .X(_09986_));
 sg13g2_nor2_1 _16554_ (.A(net10390),
    .B(_09986_),
    .Y(_09987_));
 sg13g2_a21oi_2 _16555_ (.B1(_09987_),
    .Y(_09988_),
    .A2(_09984_),
    .A1(net10390));
 sg13g2_buf_2 place10697 (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[4] ),
    .X(net10697));
 sg13g2_buf_2 place10886 (.A(net10885),
    .X(net10886));
 sg13g2_nand2_1 _16558_ (.Y(_09991_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][23] ),
    .B(net10140));
 sg13g2_o21ai_1 _16559_ (.B1(_09991_),
    .Y(_00705_),
    .A1(net10140),
    .A2(net9690));
 sg13g2_mux2_1 _16560_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[24] ),
    .S(net10629),
    .X(_09992_));
 sg13g2_inv_2 _16561_ (.Y(_09993_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[24] ));
 sg13g2_nand4_1 _16562_ (.B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[22] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.reg_pc[23] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[21] ),
    .Y(_09994_),
    .D(_09968_));
 sg13g2_xnor2_1 _16563_ (.Y(_09995_),
    .A(_09993_),
    .B(_09994_));
 sg13g2_nor2_1 _16564_ (.A(net10391),
    .B(_09995_),
    .Y(_09996_));
 sg13g2_a21oi_2 _16565_ (.B1(_09996_),
    .Y(_09997_),
    .A2(_09992_),
    .A1(net10391));
 sg13g2_buf_2 place11004 (.A(net11003),
    .X(net11004));
 sg13g2_buf_2 place10757 (.A(net10756),
    .X(net10757));
 sg13g2_nand2_1 _16568_ (.Y(_10000_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][24] ),
    .B(net10140));
 sg13g2_o21ai_1 _16569_ (.B1(_10000_),
    .Y(_00706_),
    .A1(net10140),
    .A2(net9685));
 sg13g2_mux2_1 _16570_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[25] ),
    .S(net10629),
    .X(_10001_));
 sg13g2_nor2_2 _16571_ (.A(_09993_),
    .B(_09994_),
    .Y(_10002_));
 sg13g2_xnor2_1 _16572_ (.Y(_10003_),
    .A(net10493),
    .B(_10002_));
 sg13g2_nand2_1 _16573_ (.Y(_10004_),
    .A(net10381),
    .B(_10003_));
 sg13g2_o21ai_1 _16574_ (.B1(_10004_),
    .Y(_10005_),
    .A1(net10381),
    .A2(_10001_));
 sg13g2_buf_2 place10733 (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[1] ),
    .X(net10733));
 sg13g2_buf_2 place10715 (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[1] ),
    .X(net10715));
 sg13g2_nand2_1 _16577_ (.Y(_10008_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][25] ),
    .B(net10142));
 sg13g2_o21ai_1 _16578_ (.B1(_10008_),
    .Y(_00707_),
    .A1(net10142),
    .A2(net9679));
 sg13g2_nand2_1 _16579_ (.Y(_10009_),
    .A(net10493),
    .B(_10002_));
 sg13g2_xnor2_1 _16580_ (.Y(_10010_),
    .A(net10492),
    .B(_10009_));
 sg13g2_nor2b_1 _16581_ (.A(net10629),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_out[26] ),
    .Y(_10011_));
 sg13g2_a21oi_2 _16582_ (.B1(_10011_),
    .Y(_10012_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[26] ),
    .A1(net10629));
 sg13g2_nor2_1 _16583_ (.A(net10381),
    .B(_10012_),
    .Y(_10013_));
 sg13g2_a21oi_2 _16584_ (.B1(_10013_),
    .Y(_10014_),
    .A2(_10010_),
    .A1(net10381));
 sg13g2_buf_2 place10800 (.A(net10799),
    .X(net10800));
 sg13g2_buf_2 place10668 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[9] ),
    .X(net10668));
 sg13g2_buf_2 place10672 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[4] ),
    .X(net10672));
 sg13g2_nand2_1 _16588_ (.Y(_10018_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][26] ),
    .B(net10143));
 sg13g2_o21ai_1 _16589_ (.B1(_10018_),
    .Y(_00708_),
    .A1(net10143),
    .A2(net9675));
 sg13g2_mux2_1 _16590_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[27] ),
    .S(net10629),
    .X(_10019_));
 sg13g2_nand3_1 _16591_ (.B(net10492),
    .C(_10002_),
    .A(net10493),
    .Y(_10020_));
 sg13g2_xor2_1 _16592_ (.B(_10020_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[27] ),
    .X(_10021_));
 sg13g2_nor2_1 _16593_ (.A(net10391),
    .B(_10021_),
    .Y(_10022_));
 sg13g2_a21oi_2 _16594_ (.B1(_10022_),
    .Y(_10023_),
    .A2(_10019_),
    .A1(net10391));
 sg13g2_buf_2 place10716 (.A(net10715),
    .X(net10716));
 sg13g2_buf_2 place10745 (.A(net10744),
    .X(net10745));
 sg13g2_nand2_1 _16597_ (.Y(_10026_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][27] ),
    .B(net10143));
 sg13g2_o21ai_1 _16598_ (.B1(_10026_),
    .Y(_00709_),
    .A1(net10143),
    .A2(net9651));
 sg13g2_buf_2 place10718 (.A(net10717),
    .X(net10718));
 sg13g2_mux2_1 _16600_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[28] ),
    .S(net10628),
    .X(_10028_));
 sg13g2_inv_2 _16601_ (.Y(_10029_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[28] ));
 sg13g2_nand4_1 _16602_ (.B(net10492),
    .C(\u_ac_controller_soc_inst.u_picorv32.reg_pc[27] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[25] ),
    .Y(_10030_),
    .D(_10002_));
 sg13g2_xnor2_1 _16603_ (.Y(_10031_),
    .A(_10029_),
    .B(_10030_));
 sg13g2_nor2_1 _16604_ (.A(net10391),
    .B(_10031_),
    .Y(_10032_));
 sg13g2_a21oi_2 _16605_ (.B1(_10032_),
    .Y(_10033_),
    .A2(_10028_),
    .A1(net10391));
 sg13g2_buf_2 place10700 (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[4] ),
    .X(net10700));
 sg13g2_buf_2 place10701 (.A(net10700),
    .X(net10701));
 sg13g2_nand2_1 _16608_ (.Y(_10036_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][28] ),
    .B(net10143));
 sg13g2_o21ai_1 _16609_ (.B1(_10036_),
    .Y(_00710_),
    .A1(net10143),
    .A2(net9646));
 sg13g2_mux2_1 _16610_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[29] ),
    .S(net10628),
    .X(_10037_));
 sg13g2_nor2_2 _16611_ (.A(_10029_),
    .B(_10030_),
    .Y(_10038_));
 sg13g2_xnor2_1 _16612_ (.Y(_10039_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[29] ),
    .B(_10038_));
 sg13g2_nor2_1 _16613_ (.A(net10391),
    .B(_10039_),
    .Y(_10040_));
 sg13g2_a21oi_2 _16614_ (.B1(_10040_),
    .Y(_10041_),
    .A2(_10037_),
    .A1(net10391));
 sg13g2_buf_2 place10669 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[8] ),
    .X(net10669));
 sg13g2_buf_2 place10722 (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[1] ),
    .X(net10722));
 sg13g2_nand2_1 _16617_ (.Y(_10044_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][29] ),
    .B(net10142));
 sg13g2_o21ai_1 _16618_ (.B1(_10044_),
    .Y(_00711_),
    .A1(net10142),
    .A2(net9643));
 sg13g2_mux2_1 _16619_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[2] ),
    .S(net10631),
    .X(_10045_));
 sg13g2_and2_1 _16620_ (.A(net10385),
    .B(_10045_),
    .X(_10046_));
 sg13g2_a21oi_2 _16621_ (.B1(_10046_),
    .Y(_10047_),
    .A2(_09857_),
    .A1(_00130_));
 sg13g2_buf_2 place10725 (.A(net10723),
    .X(net10725));
 sg13g2_buf_2 place10721 (.A(net10716),
    .X(net10721));
 sg13g2_nand2_1 _16624_ (.Y(_10050_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][2] ),
    .B(net10137));
 sg13g2_o21ai_1 _16625_ (.B1(_10050_),
    .Y(_00712_),
    .A1(net10137),
    .A2(net10224));
 sg13g2_nand2_1 _16626_ (.Y(_10051_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[29] ),
    .B(_10038_));
 sg13g2_xnor2_1 _16627_ (.Y(_10052_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[30] ),
    .B(_10051_));
 sg13g2_nor2b_1 _16628_ (.A(net10628),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_out[30] ),
    .Y(_10053_));
 sg13g2_a21oi_2 _16629_ (.B1(_10053_),
    .Y(_10054_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[30] ),
    .A1(net10629));
 sg13g2_nor2_1 _16630_ (.A(net10381),
    .B(_10054_),
    .Y(_10055_));
 sg13g2_a21oi_2 _16631_ (.B1(_10055_),
    .Y(_10056_),
    .A2(_10052_),
    .A1(net10381));
 sg13g2_buf_2 place10667 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20] ),
    .X(net10667));
 sg13g2_buf_2 place10724 (.A(net10723),
    .X(net10724));
 sg13g2_nand2_1 _16634_ (.Y(_10059_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][30] ),
    .B(net10141));
 sg13g2_o21ai_1 _16635_ (.B1(_10059_),
    .Y(_00713_),
    .A1(net10141),
    .A2(net9638));
 sg13g2_nand3_1 _16636_ (.B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[30] ),
    .C(_10038_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[29] ),
    .Y(_10060_));
 sg13g2_xnor2_1 _16637_ (.Y(_10061_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[31] ),
    .B(_10060_));
 sg13g2_nor2b_1 _16638_ (.A(net10628),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_out[31] ),
    .Y(_10062_));
 sg13g2_a21oi_2 _16639_ (.B1(_10062_),
    .Y(_10063_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[31] ),
    .A1(net10628));
 sg13g2_nor2_1 _16640_ (.A(net10381),
    .B(_10063_),
    .Y(_10064_));
 sg13g2_a21oi_2 _16641_ (.B1(_10064_),
    .Y(_10065_),
    .A2(_10061_),
    .A1(net10381));
 sg13g2_buf_16 clkbuf_leaf_144_clk (.X(clknet_leaf_144_clk),
    .A(clknet_8_97_0_clk));
 sg13g2_buf_16 clkbuf_leaf_143_clk (.X(clknet_leaf_143_clk),
    .A(clknet_8_98_0_clk));
 sg13g2_nand2_1 _16644_ (.Y(_10068_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][31] ),
    .B(_09852_));
 sg13g2_o21ai_1 _16645_ (.B1(_10068_),
    .Y(_00714_),
    .A1(_09852_),
    .A2(net9636));
 sg13g2_mux2_1 _16646_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[3] ),
    .S(net10631),
    .X(_10069_));
 sg13g2_xnor2_1 _16647_ (.Y(_10070_),
    .A(net10490),
    .B(net10491));
 sg13g2_nor2_1 _16648_ (.A(net10386),
    .B(_10070_),
    .Y(_10071_));
 sg13g2_a21oi_2 _16649_ (.B1(_10071_),
    .Y(_10072_),
    .A2(_10069_),
    .A1(net10386));
 sg13g2_buf_2 place10702 (.A(net10701),
    .X(net10702));
 sg13g2_buf_2 place10706 (.A(net10703),
    .X(net10706));
 sg13g2_nand2_1 _16652_ (.Y(_10075_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][3] ),
    .B(net10138));
 sg13g2_o21ai_1 _16653_ (.B1(_10075_),
    .Y(_00715_),
    .A1(net10138),
    .A2(net10220));
 sg13g2_mux2_1 _16654_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[4] ),
    .S(net10631),
    .X(_10076_));
 sg13g2_nand2_1 _16655_ (.Y(_10077_),
    .A(net10490),
    .B(net10491));
 sg13g2_xor2_1 _16656_ (.B(_10077_),
    .A(net10489),
    .X(_10078_));
 sg13g2_nor2_1 _16657_ (.A(net10386),
    .B(_10078_),
    .Y(_10079_));
 sg13g2_a21oi_2 _16658_ (.B1(_10079_),
    .Y(_10080_),
    .A2(_10076_),
    .A1(net10386));
 sg13g2_buf_2 place10703 (.A(net10701),
    .X(net10703));
 sg13g2_buf_2 place10663 (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[8] ),
    .X(net10663));
 sg13g2_nand2_1 _16661_ (.Y(_10083_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][4] ),
    .B(net10139));
 sg13g2_o21ai_1 _16662_ (.B1(_10083_),
    .Y(_00716_),
    .A1(net10139),
    .A2(net10182));
 sg13g2_mux2_1 _16663_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[5] ),
    .S(net10631),
    .X(_10084_));
 sg13g2_nand3_1 _16664_ (.B(net10491),
    .C(net10489),
    .A(net10490),
    .Y(_10085_));
 sg13g2_xor2_1 _16665_ (.B(_10085_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[5] ),
    .X(_10086_));
 sg13g2_nor2_1 _16666_ (.A(net10386),
    .B(_10086_),
    .Y(_10087_));
 sg13g2_a21oi_2 _16667_ (.B1(_10087_),
    .Y(_10088_),
    .A2(_10084_),
    .A1(net10386));
 sg13g2_buf_2 place10705 (.A(net10704),
    .X(net10705));
 sg13g2_buf_2 place10704 (.A(net10703),
    .X(net10704));
 sg13g2_nand2_1 _16670_ (.Y(_10091_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][5] ),
    .B(net10137));
 sg13g2_o21ai_1 _16671_ (.B1(_10091_),
    .Y(_00717_),
    .A1(net10137),
    .A2(net10178));
 sg13g2_mux2_1 _16672_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[6] ),
    .S(net10631),
    .X(_10092_));
 sg13g2_xnor2_1 _16673_ (.Y(_10093_),
    .A(_09285_),
    .B(_09862_));
 sg13g2_nor2_1 _16674_ (.A(net10385),
    .B(_10093_),
    .Y(_10094_));
 sg13g2_a21oi_2 _16675_ (.B1(_10094_),
    .Y(_10095_),
    .A2(_10092_),
    .A1(net10385));
 sg13g2_buf_2 place10707 (.A(net10706),
    .X(net10707));
 sg13g2_buf_2 place10655 (.A(net10653),
    .X(net10655));
 sg13g2_nand2_1 _16678_ (.Y(_10098_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][6] ),
    .B(net10136));
 sg13g2_o21ai_1 _16679_ (.B1(_10098_),
    .Y(_00718_),
    .A1(net10136),
    .A2(net10172));
 sg13g2_nor2_1 _16680_ (.A(_09285_),
    .B(_09862_),
    .Y(_10099_));
 sg13g2_xnor2_1 _16681_ (.Y(_10100_),
    .A(_09861_),
    .B(_10099_));
 sg13g2_mux2_1 _16682_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[7] ),
    .S(net10631),
    .X(_10101_));
 sg13g2_and2_1 _16683_ (.A(net10385),
    .B(_10101_),
    .X(_10102_));
 sg13g2_a21oi_2 _16684_ (.B1(_10102_),
    .Y(_10103_),
    .A2(_10100_),
    .A1(_09857_));
 sg13g2_buf_2 place10662 (.A(net10661),
    .X(net10662));
 sg13g2_buf_2 place10666 (.A(net10664),
    .X(net10666));
 sg13g2_nand2_1 _16687_ (.Y(_10106_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][7] ),
    .B(net10136));
 sg13g2_o21ai_1 _16688_ (.B1(_10106_),
    .Y(_00719_),
    .A1(net10136),
    .A2(net10167));
 sg13g2_mux2_1 _16689_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[8] ),
    .S(net10630),
    .X(_10107_));
 sg13g2_nor3_1 _16690_ (.A(_09285_),
    .B(_09861_),
    .C(_09862_),
    .Y(_10108_));
 sg13g2_xnor2_1 _16691_ (.Y(_10109_),
    .A(net10488),
    .B(_10108_));
 sg13g2_nor2_1 _16692_ (.A(net10384),
    .B(_10109_),
    .Y(_10110_));
 sg13g2_a21oi_2 _16693_ (.B1(_10110_),
    .Y(_10111_),
    .A2(_10107_),
    .A1(net10384));
 sg13g2_buf_2 place10654 (.A(net10653),
    .X(net10654));
 sg13g2_buf_2 place10653 (.A(net10652),
    .X(net10653));
 sg13g2_nand2_1 _16696_ (.Y(_10114_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][8] ),
    .B(net10135));
 sg13g2_o21ai_1 _16697_ (.B1(_10114_),
    .Y(_00720_),
    .A1(net10135),
    .A2(net10128));
 sg13g2_mux2_1 _16698_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_out[9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[9] ),
    .S(net10630),
    .X(_10115_));
 sg13g2_nand2_1 _16699_ (.Y(_10116_),
    .A(net10488),
    .B(_10108_));
 sg13g2_xor2_1 _16700_ (.B(_10116_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[9] ),
    .X(_10117_));
 sg13g2_nor2_1 _16701_ (.A(_09828_),
    .B(_10117_),
    .Y(_10118_));
 sg13g2_a21oi_2 _16702_ (.B1(_10118_),
    .Y(_10119_),
    .A2(_10115_),
    .A1(net10386));
 sg13g2_buf_2 place10650 (.A(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycleh ),
    .X(net10650));
 sg13g2_buf_2 place10644 (.A(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstr ),
    .X(net10644));
 sg13g2_nand2_1 _16705_ (.Y(_10122_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][9] ),
    .B(net10136));
 sg13g2_o21ai_1 _16706_ (.B1(_10122_),
    .Y(_00721_),
    .A1(net10136),
    .A2(net9975));
 sg13g2_inv_1 _16707_ (.Y(_10123_),
    .A(_09849_));
 sg13g2_and3_2 _16708_ (.X(_10124_),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[1] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_rd[0] ),
    .C(_10123_));
 sg13g2_buf_2 place10639 (.A(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh ),
    .X(net10639));
 sg13g2_nand2_2 _16710_ (.Y(_10126_),
    .A(_09843_),
    .B(_10124_));
 sg13g2_buf_2 place10637 (.A(net10636),
    .X(net10637));
 sg13g2_buf_2 place10627 (.A(\u_ac_controller_soc_inst.u_picorv32.latched_stalu ),
    .X(net10627));
 sg13g2_buf_2 place10710 (.A(net10709),
    .X(net10710));
 sg13g2_nand2_1 _16714_ (.Y(_10130_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][0] ),
    .B(net9965));
 sg13g2_o21ai_1 _16715_ (.B1(_10130_),
    .Y(_00722_),
    .A1(net10279),
    .A2(net9965));
 sg13g2_nand2_1 _16716_ (.Y(_10131_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][10] ),
    .B(net9968));
 sg13g2_o21ai_1 _16717_ (.B1(_10131_),
    .Y(_00723_),
    .A1(net10131),
    .A2(net9968));
 sg13g2_nand2_1 _16718_ (.Y(_10132_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][11] ),
    .B(net9972));
 sg13g2_o21ai_1 _16719_ (.B1(_10132_),
    .Y(_00724_),
    .A1(net9985),
    .A2(net9972));
 sg13g2_nand2_1 _16720_ (.Y(_10133_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][12] ),
    .B(net9966));
 sg13g2_o21ai_1 _16721_ (.B1(_10133_),
    .Y(_00725_),
    .A1(net9801),
    .A2(net9966));
 sg13g2_nand2_1 _16722_ (.Y(_10134_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][13] ),
    .B(net9965));
 sg13g2_o21ai_1 _16723_ (.B1(_10134_),
    .Y(_00726_),
    .A1(net9981),
    .A2(net9965));
 sg13g2_nand2_1 _16724_ (.Y(_10135_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][14] ),
    .B(net9969));
 sg13g2_o21ai_1 _16725_ (.B1(_10135_),
    .Y(_00727_),
    .A1(net9795),
    .A2(net9969));
 sg13g2_nand2_1 _16726_ (.Y(_10136_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][15] ),
    .B(net9968));
 sg13g2_o21ai_1 _16727_ (.B1(_10136_),
    .Y(_00728_),
    .A1(net9793),
    .A2(net9968));
 sg13g2_nand2_1 _16728_ (.Y(_10137_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][16] ),
    .B(net9968));
 sg13g2_o21ai_1 _16729_ (.B1(_10137_),
    .Y(_00729_),
    .A1(net9745),
    .A2(net9968));
 sg13g2_buf_2 place10661 (.A(\u_ac_controller_soc_inst.u_picorv32.decoder_trigger ),
    .X(net10661));
 sg13g2_nand2_1 _16731_ (.Y(_10139_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][17] ),
    .B(net9967));
 sg13g2_o21ai_1 _16732_ (.B1(_10139_),
    .Y(_00730_),
    .A1(net9742),
    .A2(net9967));
 sg13g2_nand2_1 _16733_ (.Y(_10140_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][18] ),
    .B(net9970));
 sg13g2_o21ai_1 _16734_ (.B1(_10140_),
    .Y(_00731_),
    .A1(net9738),
    .A2(net9970));
 sg13g2_buf_2 place10626 (.A(\u_ac_controller_soc_inst.cbus_addr[11] ),
    .X(net10626));
 sg13g2_nand2_1 _16736_ (.Y(_10142_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][19] ),
    .B(net9973));
 sg13g2_o21ai_1 _16737_ (.B1(_10142_),
    .Y(_00732_),
    .A1(net9724),
    .A2(net9973));
 sg13g2_nand2_1 _16738_ (.Y(_10143_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][1] ),
    .B(net9965));
 sg13g2_o21ai_1 _16739_ (.B1(_10143_),
    .Y(_00733_),
    .A1(net10227),
    .A2(net9965));
 sg13g2_nand2_1 _16740_ (.Y(_10144_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][20] ),
    .B(net9971));
 sg13g2_o21ai_1 _16741_ (.B1(_10144_),
    .Y(_00734_),
    .A1(net9718),
    .A2(net9971));
 sg13g2_nand2_1 _16742_ (.Y(_10145_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][21] ),
    .B(net9971));
 sg13g2_o21ai_1 _16743_ (.B1(_10145_),
    .Y(_00735_),
    .A1(net9714),
    .A2(net9971));
 sg13g2_nand2_1 _16744_ (.Y(_10146_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][22] ),
    .B(net9970));
 sg13g2_o21ai_1 _16745_ (.B1(_10146_),
    .Y(_00736_),
    .A1(net9696),
    .A2(net9970));
 sg13g2_nand2_1 _16746_ (.Y(_10147_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][23] ),
    .B(net9970));
 sg13g2_o21ai_1 _16747_ (.B1(_10147_),
    .Y(_00737_),
    .A1(net9691),
    .A2(net9971));
 sg13g2_nand2_1 _16748_ (.Y(_10148_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][24] ),
    .B(net9970));
 sg13g2_o21ai_1 _16749_ (.B1(_10148_),
    .Y(_00738_),
    .A1(net9685),
    .A2(net9970));
 sg13g2_nand2_1 _16750_ (.Y(_10149_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][25] ),
    .B(net9972));
 sg13g2_o21ai_1 _16751_ (.B1(_10149_),
    .Y(_00739_),
    .A1(net9679),
    .A2(net9972));
 sg13g2_buf_2 place10649 (.A(net10647),
    .X(net10649));
 sg13g2_nand2_1 _16753_ (.Y(_10151_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][26] ),
    .B(net9973));
 sg13g2_o21ai_1 _16754_ (.B1(_10151_),
    .Y(_00740_),
    .A1(net9675),
    .A2(net9973));
 sg13g2_nand2_1 _16755_ (.Y(_10152_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][27] ),
    .B(net9973));
 sg13g2_o21ai_1 _16756_ (.B1(_10152_),
    .Y(_00741_),
    .A1(_10023_),
    .A2(net9973));
 sg13g2_buf_2 place10625 (.A(\u_ac_controller_soc_inst.cbus_addr[13] ),
    .X(net10625));
 sg13g2_nand2_1 _16758_ (.Y(_10154_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][28] ),
    .B(net9973));
 sg13g2_o21ai_1 _16759_ (.B1(_10154_),
    .Y(_00742_),
    .A1(net9646),
    .A2(net9973));
 sg13g2_nand2_1 _16760_ (.Y(_10155_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][29] ),
    .B(net9972));
 sg13g2_o21ai_1 _16761_ (.B1(_10155_),
    .Y(_00743_),
    .A1(_10041_),
    .A2(net9972));
 sg13g2_nand2_1 _16762_ (.Y(_10156_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][2] ),
    .B(net9967));
 sg13g2_o21ai_1 _16763_ (.B1(_10156_),
    .Y(_00744_),
    .A1(net10222),
    .A2(net9967));
 sg13g2_nand2_1 _16764_ (.Y(_10157_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][30] ),
    .B(net9969));
 sg13g2_o21ai_1 _16765_ (.B1(_10157_),
    .Y(_00745_),
    .A1(net9638),
    .A2(net9969));
 sg13g2_nand2_1 _16766_ (.Y(_10158_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][31] ),
    .B(net9969));
 sg13g2_o21ai_1 _16767_ (.B1(_10158_),
    .Y(_00746_),
    .A1(net9636),
    .A2(net9969));
 sg13g2_nand2_1 _16768_ (.Y(_10159_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][3] ),
    .B(net9968));
 sg13g2_o21ai_1 _16769_ (.B1(_10159_),
    .Y(_00747_),
    .A1(net10221),
    .A2(net9968));
 sg13g2_nand2_1 _16770_ (.Y(_10160_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][4] ),
    .B(net9971));
 sg13g2_o21ai_1 _16771_ (.B1(_10160_),
    .Y(_00748_),
    .A1(net10181),
    .A2(net9971));
 sg13g2_nand2_1 _16772_ (.Y(_10161_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][5] ),
    .B(net9967));
 sg13g2_o21ai_1 _16773_ (.B1(_10161_),
    .Y(_00749_),
    .A1(net10174),
    .A2(net9967));
 sg13g2_nand2_1 _16774_ (.Y(_10162_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][6] ),
    .B(net9966));
 sg13g2_o21ai_1 _16775_ (.B1(_10162_),
    .Y(_00750_),
    .A1(net10171),
    .A2(net9966));
 sg13g2_nand2_1 _16776_ (.Y(_10163_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][7] ),
    .B(net9966));
 sg13g2_o21ai_1 _16777_ (.B1(_10163_),
    .Y(_00751_),
    .A1(net10167),
    .A2(net9966));
 sg13g2_nand2_1 _16778_ (.Y(_10164_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][8] ),
    .B(_10126_));
 sg13g2_o21ai_1 _16779_ (.B1(_10164_),
    .Y(_00752_),
    .A1(net10128),
    .A2(_10126_));
 sg13g2_nand2_1 _16780_ (.Y(_10165_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][9] ),
    .B(net9966));
 sg13g2_o21ai_1 _16781_ (.B1(_10165_),
    .Y(_00753_),
    .A1(net9975),
    .A2(net9966));
 sg13g2_buf_2 place10660 (.A(\u_ac_controller_soc_inst.u_picorv32.decoder_trigger ),
    .X(net10660));
 sg13g2_nor2_2 _16783_ (.A(_00084_),
    .B(_09842_),
    .Y(_10167_));
 sg13g2_nor3_2 _16784_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[4] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_rd[3] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.latched_rd[2] ),
    .Y(_10168_));
 sg13g2_nor4_2 _16785_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[1] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_rd[0] ),
    .C(_09849_),
    .Y(_10169_),
    .D(_10168_));
 sg13g2_buf_2 place10657 (.A(net10652),
    .X(net10657));
 sg13g2_nand2_2 _16787_ (.Y(_10171_),
    .A(_10167_),
    .B(_10169_));
 sg13g2_buf_2 place10624 (.A(\u_ac_controller_soc_inst.cbus_addr[20] ),
    .X(net10624));
 sg13g2_buf_2 place10647 (.A(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycleh ),
    .X(net10647));
 sg13g2_buf_2 place10623 (.A(\u_ac_controller_soc_inst.cbus_addr[21] ),
    .X(net10623));
 sg13g2_nand2_1 _16791_ (.Y(_10175_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][0] ),
    .B(net10122));
 sg13g2_o21ai_1 _16792_ (.B1(_10175_),
    .Y(_00754_),
    .A1(net10277),
    .A2(net10122));
 sg13g2_nand2_1 _16793_ (.Y(_10176_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][10] ),
    .B(net10123));
 sg13g2_o21ai_1 _16794_ (.B1(_10176_),
    .Y(_00755_),
    .A1(net10131),
    .A2(net10123));
 sg13g2_nand2_1 _16795_ (.Y(_10177_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][11] ),
    .B(net10119));
 sg13g2_o21ai_1 _16796_ (.B1(_10177_),
    .Y(_00756_),
    .A1(net9985),
    .A2(net10119));
 sg13g2_nand2_1 _16797_ (.Y(_10178_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][12] ),
    .B(net10125));
 sg13g2_o21ai_1 _16798_ (.B1(_10178_),
    .Y(_00757_),
    .A1(net9800),
    .A2(net10125));
 sg13g2_nand2_1 _16799_ (.Y(_10179_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][13] ),
    .B(net10122));
 sg13g2_o21ai_1 _16800_ (.B1(_10179_),
    .Y(_00758_),
    .A1(net9979),
    .A2(net10122));
 sg13g2_nand2_1 _16801_ (.Y(_10180_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][14] ),
    .B(net10119));
 sg13g2_o21ai_1 _16802_ (.B1(_10180_),
    .Y(_00759_),
    .A1(net9798),
    .A2(net10118));
 sg13g2_nand2_1 _16803_ (.Y(_10181_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][15] ),
    .B(net10123));
 sg13g2_o21ai_1 _16804_ (.B1(_10181_),
    .Y(_00760_),
    .A1(net9791),
    .A2(net10123));
 sg13g2_nand2_1 _16805_ (.Y(_10182_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][16] ),
    .B(net10123));
 sg13g2_o21ai_1 _16806_ (.B1(_10182_),
    .Y(_00761_),
    .A1(net9745),
    .A2(net10123));
 sg13g2_buf_2 place10622 (.A(\u_ac_controller_soc_inst.cbus_addr[23] ),
    .X(net10622));
 sg13g2_nand2_1 _16808_ (.Y(_10184_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][17] ),
    .B(net10124));
 sg13g2_o21ai_1 _16809_ (.B1(_10184_),
    .Y(_00762_),
    .A1(net9742),
    .A2(net10124));
 sg13g2_nand2_1 _16810_ (.Y(_10185_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][18] ),
    .B(net10118));
 sg13g2_o21ai_1 _16811_ (.B1(_10185_),
    .Y(_00763_),
    .A1(net9738),
    .A2(net10118));
 sg13g2_buf_2 place10633 (.A(\u_ac_controller_soc_inst.u_picorv32.instr_sub ),
    .X(net10633));
 sg13g2_nand2_1 _16813_ (.Y(_10187_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][19] ),
    .B(net10121));
 sg13g2_o21ai_1 _16814_ (.B1(_10187_),
    .Y(_00764_),
    .A1(net9724),
    .A2(net10121));
 sg13g2_nand2_1 _16815_ (.Y(_10188_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][1] ),
    .B(net10124));
 sg13g2_o21ai_1 _16816_ (.B1(_10188_),
    .Y(_00765_),
    .A1(net10227),
    .A2(net10124));
 sg13g2_nand2_1 _16817_ (.Y(_10189_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][20] ),
    .B(net10117));
 sg13g2_o21ai_1 _16818_ (.B1(_10189_),
    .Y(_00766_),
    .A1(net9719),
    .A2(net10117));
 sg13g2_nand2_1 _16819_ (.Y(_10190_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][21] ),
    .B(_10171_));
 sg13g2_o21ai_1 _16820_ (.B1(_10190_),
    .Y(_00767_),
    .A1(net9713),
    .A2(_10171_));
 sg13g2_nand2_1 _16821_ (.Y(_10191_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][22] ),
    .B(net10117));
 sg13g2_o21ai_1 _16822_ (.B1(_10191_),
    .Y(_00768_),
    .A1(net9695),
    .A2(net10117));
 sg13g2_nand2_1 _16823_ (.Y(_10192_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][23] ),
    .B(net10117));
 sg13g2_o21ai_1 _16824_ (.B1(_10192_),
    .Y(_00769_),
    .A1(net9692),
    .A2(net10117));
 sg13g2_nand2_1 _16825_ (.Y(_10193_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][24] ),
    .B(net10117));
 sg13g2_o21ai_1 _16826_ (.B1(_10193_),
    .Y(_00770_),
    .A1(net9687),
    .A2(net10117));
 sg13g2_nand2_1 _16827_ (.Y(_10194_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][25] ),
    .B(net10120));
 sg13g2_o21ai_1 _16828_ (.B1(_10194_),
    .Y(_00771_),
    .A1(net9679),
    .A2(net10120));
 sg13g2_buf_2 place10628 (.A(net10627),
    .X(net10628));
 sg13g2_nand2_1 _16830_ (.Y(_10196_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][26] ),
    .B(net10121));
 sg13g2_o21ai_1 _16831_ (.B1(_10196_),
    .Y(_00772_),
    .A1(net9674),
    .A2(net10121));
 sg13g2_nand2_1 _16832_ (.Y(_10197_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][27] ),
    .B(net10121));
 sg13g2_o21ai_1 _16833_ (.B1(_10197_),
    .Y(_00773_),
    .A1(_10023_),
    .A2(net10121));
 sg13g2_buf_2 place10618 (.A(\u_ac_controller_soc_inst.cbus_addr[3] ),
    .X(net10618));
 sg13g2_nand2_1 _16835_ (.Y(_10199_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][28] ),
    .B(net10121));
 sg13g2_o21ai_1 _16836_ (.B1(_10199_),
    .Y(_00774_),
    .A1(net9647),
    .A2(net10121));
 sg13g2_nand2_1 _16837_ (.Y(_10200_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][29] ),
    .B(net10120));
 sg13g2_o21ai_1 _16838_ (.B1(_10200_),
    .Y(_00775_),
    .A1(_10041_),
    .A2(net10120));
 sg13g2_nand2_1 _16839_ (.Y(_10201_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][2] ),
    .B(net10124));
 sg13g2_o21ai_1 _16840_ (.B1(_10201_),
    .Y(_00776_),
    .A1(net10224),
    .A2(net10124));
 sg13g2_nand2_1 _16841_ (.Y(_10202_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][30] ),
    .B(net10119));
 sg13g2_o21ai_1 _16842_ (.B1(_10202_),
    .Y(_00777_),
    .A1(net9638),
    .A2(net10119));
 sg13g2_nand2_1 _16843_ (.Y(_10203_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][31] ),
    .B(net10119));
 sg13g2_o21ai_1 _16844_ (.B1(_10203_),
    .Y(_00778_),
    .A1(net9635),
    .A2(net10119));
 sg13g2_nand2_1 _16845_ (.Y(_10204_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][3] ),
    .B(net10123));
 sg13g2_o21ai_1 _16846_ (.B1(_10204_),
    .Y(_00779_),
    .A1(net10220),
    .A2(net10123));
 sg13g2_nand2_1 _16847_ (.Y(_10205_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][4] ),
    .B(_10171_));
 sg13g2_o21ai_1 _16848_ (.B1(_10205_),
    .Y(_00780_),
    .A1(net10182),
    .A2(_10171_));
 sg13g2_nand2_1 _16849_ (.Y(_10206_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][5] ),
    .B(net10124));
 sg13g2_o21ai_1 _16850_ (.B1(_10206_),
    .Y(_00781_),
    .A1(_10088_),
    .A2(net10124));
 sg13g2_nand2_1 _16851_ (.Y(_10207_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][6] ),
    .B(net10125));
 sg13g2_o21ai_1 _16852_ (.B1(_10207_),
    .Y(_00782_),
    .A1(net10171),
    .A2(net10125));
 sg13g2_nand2_1 _16853_ (.Y(_10208_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][7] ),
    .B(net10125));
 sg13g2_o21ai_1 _16854_ (.B1(_10208_),
    .Y(_00783_),
    .A1(net10167),
    .A2(net10125));
 sg13g2_nand2_1 _16855_ (.Y(_10209_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][8] ),
    .B(net10118));
 sg13g2_o21ai_1 _16856_ (.B1(_10209_),
    .Y(_00784_),
    .A1(_10111_),
    .A2(net10118));
 sg13g2_nand2_1 _16857_ (.Y(_10210_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][9] ),
    .B(net10125));
 sg13g2_o21ai_1 _16858_ (.B1(_10210_),
    .Y(_00785_),
    .A1(net9975),
    .A2(net10125));
 sg13g2_and3_2 _16859_ (.X(_10211_),
    .A(_09845_),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_rd[0] ),
    .C(_10123_));
 sg13g2_buf_2 place10629 (.A(net10628),
    .X(net10629));
 sg13g2_nand2_2 _16861_ (.Y(_10213_),
    .A(_10167_),
    .B(_10211_));
 sg13g2_buf_2 place10615 (.A(\u_ac_controller_soc_inst.cbus_addr[5] ),
    .X(net10615));
 sg13g2_buf_2 place10614 (.A(\u_ac_controller_soc_inst.cbus_addr[6] ),
    .X(net10614));
 sg13g2_buf_2 place10616 (.A(\u_ac_controller_soc_inst.cbus_addr[5] ),
    .X(net10616));
 sg13g2_nand2_1 _16865_ (.Y(_10217_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][0] ),
    .B(_10213_));
 sg13g2_o21ai_1 _16866_ (.B1(_10217_),
    .Y(_00786_),
    .A1(net10277),
    .A2(net9955));
 sg13g2_nand2_1 _16867_ (.Y(_10218_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][10] ),
    .B(net9957));
 sg13g2_o21ai_1 _16868_ (.B1(_10218_),
    .Y(_00787_),
    .A1(net10131),
    .A2(net9957));
 sg13g2_nand2_1 _16869_ (.Y(_10219_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][11] ),
    .B(net9964));
 sg13g2_o21ai_1 _16870_ (.B1(_10219_),
    .Y(_00788_),
    .A1(net9985),
    .A2(net9962));
 sg13g2_nand2_1 _16871_ (.Y(_10220_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][12] ),
    .B(net9955));
 sg13g2_o21ai_1 _16872_ (.B1(_10220_),
    .Y(_00789_),
    .A1(net9800),
    .A2(net9956));
 sg13g2_nand2_1 _16873_ (.Y(_10221_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][13] ),
    .B(net9955));
 sg13g2_o21ai_1 _16874_ (.B1(_10221_),
    .Y(_00790_),
    .A1(net9979),
    .A2(net9955));
 sg13g2_nand2_1 _16875_ (.Y(_10222_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][14] ),
    .B(net9961));
 sg13g2_o21ai_1 _16876_ (.B1(_10222_),
    .Y(_00791_),
    .A1(net9798),
    .A2(net9961));
 sg13g2_nand2_1 _16877_ (.Y(_10223_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][15] ),
    .B(net9957));
 sg13g2_o21ai_1 _16878_ (.B1(_10223_),
    .Y(_00792_),
    .A1(net9791),
    .A2(net9957));
 sg13g2_nand2_1 _16879_ (.Y(_10224_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][16] ),
    .B(net9958));
 sg13g2_o21ai_1 _16880_ (.B1(_10224_),
    .Y(_00793_),
    .A1(net9744),
    .A2(net9958));
 sg13g2_buf_2 place10612 (.A(\u_ac_controller_soc_inst.cbus_addr[8] ),
    .X(net10612));
 sg13g2_nand2_1 _16882_ (.Y(_10226_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][17] ),
    .B(net9958));
 sg13g2_o21ai_1 _16883_ (.B1(_10226_),
    .Y(_00794_),
    .A1(net9742),
    .A2(net9958));
 sg13g2_nand2_1 _16884_ (.Y(_10227_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][18] ),
    .B(net9961));
 sg13g2_o21ai_1 _16885_ (.B1(_10227_),
    .Y(_00795_),
    .A1(net9738),
    .A2(net9959));
 sg13g2_buf_2 place10611 (.A(\u_ac_controller_soc_inst.cbus_addr[9] ),
    .X(net10611));
 sg13g2_nand2_1 _16887_ (.Y(_10229_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][19] ),
    .B(net9963));
 sg13g2_o21ai_1 _16888_ (.B1(_10229_),
    .Y(_00796_),
    .A1(net9724),
    .A2(net9963));
 sg13g2_nand2_1 _16889_ (.Y(_10230_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][1] ),
    .B(net9955));
 sg13g2_o21ai_1 _16890_ (.B1(_10230_),
    .Y(_00797_),
    .A1(net10227),
    .A2(net9955));
 sg13g2_nand2_1 _16891_ (.Y(_10231_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][20] ),
    .B(net9960));
 sg13g2_o21ai_1 _16892_ (.B1(_10231_),
    .Y(_00798_),
    .A1(net9719),
    .A2(net9960));
 sg13g2_nand2_1 _16893_ (.Y(_10232_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][21] ),
    .B(net9959));
 sg13g2_o21ai_1 _16894_ (.B1(_10232_),
    .Y(_00799_),
    .A1(net9714),
    .A2(net9959));
 sg13g2_nand2_1 _16895_ (.Y(_10233_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][22] ),
    .B(net9960));
 sg13g2_o21ai_1 _16896_ (.B1(_10233_),
    .Y(_00800_),
    .A1(net9695),
    .A2(net9960));
 sg13g2_nand2_1 _16897_ (.Y(_10234_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][23] ),
    .B(net9960));
 sg13g2_o21ai_1 _16898_ (.B1(_10234_),
    .Y(_00801_),
    .A1(net9692),
    .A2(net9960));
 sg13g2_nand2_1 _16899_ (.Y(_10235_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][24] ),
    .B(net9960));
 sg13g2_o21ai_1 _16900_ (.B1(_10235_),
    .Y(_00802_),
    .A1(net9687),
    .A2(net9960));
 sg13g2_nand2_1 _16901_ (.Y(_10236_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][25] ),
    .B(net9964));
 sg13g2_o21ai_1 _16902_ (.B1(_10236_),
    .Y(_00803_),
    .A1(net9679),
    .A2(net9964));
 sg13g2_buf_2 place10610 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_do_rdata ),
    .X(net10610));
 sg13g2_nand2_1 _16904_ (.Y(_10238_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][26] ),
    .B(net9963));
 sg13g2_o21ai_1 _16905_ (.B1(_10238_),
    .Y(_00804_),
    .A1(net9674),
    .A2(net9963));
 sg13g2_nand2_1 _16906_ (.Y(_10239_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][27] ),
    .B(net9963));
 sg13g2_o21ai_1 _16907_ (.B1(_10239_),
    .Y(_00805_),
    .A1(_10023_),
    .A2(net9963));
 sg13g2_buf_2 place10648 (.A(net10647),
    .X(net10648));
 sg13g2_nand2_1 _16909_ (.Y(_10241_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][28] ),
    .B(net9963));
 sg13g2_o21ai_1 _16910_ (.B1(_10241_),
    .Y(_00806_),
    .A1(net9647),
    .A2(net9963));
 sg13g2_nand2_1 _16911_ (.Y(_10242_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][29] ),
    .B(net9964));
 sg13g2_o21ai_1 _16912_ (.B1(_10242_),
    .Y(_00807_),
    .A1(_10041_),
    .A2(net9964));
 sg13g2_nand2_1 _16913_ (.Y(_10243_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][2] ),
    .B(net9958));
 sg13g2_o21ai_1 _16914_ (.B1(_10243_),
    .Y(_00808_),
    .A1(net10224),
    .A2(net9958));
 sg13g2_nand2_1 _16915_ (.Y(_10244_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][30] ),
    .B(net9962));
 sg13g2_o21ai_1 _16916_ (.B1(_10244_),
    .Y(_00809_),
    .A1(net9638),
    .A2(net9962));
 sg13g2_nand2_1 _16917_ (.Y(_10245_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][31] ),
    .B(net9962));
 sg13g2_o21ai_1 _16918_ (.B1(_10245_),
    .Y(_00810_),
    .A1(net9635),
    .A2(net9961));
 sg13g2_nand2_1 _16919_ (.Y(_10246_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][3] ),
    .B(net9957));
 sg13g2_o21ai_1 _16920_ (.B1(_10246_),
    .Y(_00811_),
    .A1(net10220),
    .A2(net9957));
 sg13g2_nand2_1 _16921_ (.Y(_10247_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][4] ),
    .B(net9959));
 sg13g2_o21ai_1 _16922_ (.B1(_10247_),
    .Y(_00812_),
    .A1(net10182),
    .A2(net9959));
 sg13g2_nand2_1 _16923_ (.Y(_10248_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][5] ),
    .B(net9958));
 sg13g2_o21ai_1 _16924_ (.B1(_10248_),
    .Y(_00813_),
    .A1(_10088_),
    .A2(net9958));
 sg13g2_nand2_1 _16925_ (.Y(_10249_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][6] ),
    .B(net9956));
 sg13g2_o21ai_1 _16926_ (.B1(_10249_),
    .Y(_00814_),
    .A1(net10171),
    .A2(net9956));
 sg13g2_nand2_1 _16927_ (.Y(_10250_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][7] ),
    .B(net9956));
 sg13g2_o21ai_1 _16928_ (.B1(_10250_),
    .Y(_00815_),
    .A1(net10167),
    .A2(net9956));
 sg13g2_nand2_1 _16929_ (.Y(_10251_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][8] ),
    .B(net9961));
 sg13g2_o21ai_1 _16930_ (.B1(_10251_),
    .Y(_00816_),
    .A1(net10127),
    .A2(net9961));
 sg13g2_nand2_1 _16931_ (.Y(_10252_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][9] ),
    .B(net9956));
 sg13g2_o21ai_1 _16932_ (.B1(_10252_),
    .Y(_00817_),
    .A1(net9975),
    .A2(net9956));
 sg13g2_nand2_2 _16933_ (.Y(_10253_),
    .A(_09850_),
    .B(_10167_));
 sg13g2_buf_2 place10609 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_do_wdata ),
    .X(net10609));
 sg13g2_buf_2 place10608 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[12] ),
    .X(net10608));
 sg13g2_buf_16 clkbuf_leaf_145_clk (.X(clknet_leaf_145_clk),
    .A(clknet_8_96_0_clk));
 sg13g2_nand2_1 _16937_ (.Y(_10257_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][0] ),
    .B(_10253_));
 sg13g2_o21ai_1 _16938_ (.B1(_10257_),
    .Y(_00818_),
    .A1(net10277),
    .A2(net10107));
 sg13g2_nand2_1 _16939_ (.Y(_10258_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][10] ),
    .B(net10108));
 sg13g2_o21ai_1 _16940_ (.B1(_10258_),
    .Y(_00819_),
    .A1(net10131),
    .A2(net10108));
 sg13g2_nand2_1 _16941_ (.Y(_10259_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][11] ),
    .B(net10112));
 sg13g2_o21ai_1 _16942_ (.B1(_10259_),
    .Y(_00820_),
    .A1(_09877_),
    .A2(net10112));
 sg13g2_nand2_1 _16943_ (.Y(_10260_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][12] ),
    .B(net10110));
 sg13g2_o21ai_1 _16944_ (.B1(_10260_),
    .Y(_00821_),
    .A1(net9800),
    .A2(net10110));
 sg13g2_nand2_1 _16945_ (.Y(_10261_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][13] ),
    .B(net10107));
 sg13g2_o21ai_1 _16946_ (.B1(_10261_),
    .Y(_00822_),
    .A1(net9979),
    .A2(net10107));
 sg13g2_nand2_1 _16947_ (.Y(_10262_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][14] ),
    .B(net10111));
 sg13g2_o21ai_1 _16948_ (.B1(_10262_),
    .Y(_00823_),
    .A1(net9798),
    .A2(net10111));
 sg13g2_nand2_1 _16949_ (.Y(_10263_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][15] ),
    .B(net10108));
 sg13g2_o21ai_1 _16950_ (.B1(_10263_),
    .Y(_00824_),
    .A1(net9791),
    .A2(net10108));
 sg13g2_nand2_1 _16951_ (.Y(_10264_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][16] ),
    .B(net10108));
 sg13g2_o21ai_1 _16952_ (.B1(_10264_),
    .Y(_00825_),
    .A1(net9745),
    .A2(net10108));
 sg13g2_buf_2 place10652 (.A(\u_ac_controller_soc_inst.u_picorv32.instr_jal ),
    .X(net10652));
 sg13g2_nand2_1 _16954_ (.Y(_10266_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][17] ),
    .B(net10109));
 sg13g2_o21ai_1 _16955_ (.B1(_10266_),
    .Y(_00826_),
    .A1(net9742),
    .A2(net10109));
 sg13g2_nand2_1 _16956_ (.Y(_10267_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][18] ),
    .B(net10115));
 sg13g2_o21ai_1 _16957_ (.B1(_10267_),
    .Y(_00827_),
    .A1(net9738),
    .A2(net10115));
 sg13g2_buf_2 place10607 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[13] ),
    .X(net10607));
 sg13g2_nand2_1 _16959_ (.Y(_10269_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][19] ),
    .B(net10114));
 sg13g2_o21ai_1 _16960_ (.B1(_10269_),
    .Y(_00828_),
    .A1(net9724),
    .A2(net10114));
 sg13g2_nand2_1 _16961_ (.Y(_10270_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][1] ),
    .B(net10107));
 sg13g2_o21ai_1 _16962_ (.B1(_10270_),
    .Y(_00829_),
    .A1(net10227),
    .A2(net10107));
 sg13g2_nand2_1 _16963_ (.Y(_10271_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][20] ),
    .B(net10116));
 sg13g2_o21ai_1 _16964_ (.B1(_10271_),
    .Y(_00830_),
    .A1(net9719),
    .A2(net10116));
 sg13g2_nand2_1 _16965_ (.Y(_10272_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][21] ),
    .B(net10115));
 sg13g2_o21ai_1 _16966_ (.B1(_10272_),
    .Y(_00831_),
    .A1(net9713),
    .A2(net10115));
 sg13g2_nand2_1 _16967_ (.Y(_10273_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][22] ),
    .B(net10116));
 sg13g2_o21ai_1 _16968_ (.B1(_10273_),
    .Y(_00832_),
    .A1(net9695),
    .A2(net10116));
 sg13g2_nand2_1 _16969_ (.Y(_10274_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][23] ),
    .B(net10116));
 sg13g2_o21ai_1 _16970_ (.B1(_10274_),
    .Y(_00833_),
    .A1(net9692),
    .A2(net10116));
 sg13g2_nand2_1 _16971_ (.Y(_10275_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][24] ),
    .B(net10116));
 sg13g2_o21ai_1 _16972_ (.B1(_10275_),
    .Y(_00834_),
    .A1(net9687),
    .A2(net10116));
 sg13g2_nand2_1 _16973_ (.Y(_10276_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][25] ),
    .B(net10113));
 sg13g2_o21ai_1 _16974_ (.B1(_10276_),
    .Y(_00835_),
    .A1(net9679),
    .A2(net10113));
 sg13g2_buf_2 place10621 (.A(net10620),
    .X(net10621));
 sg13g2_nand2_1 _16976_ (.Y(_10278_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][26] ),
    .B(net10114));
 sg13g2_o21ai_1 _16977_ (.B1(_10278_),
    .Y(_00836_),
    .A1(net9674),
    .A2(net10114));
 sg13g2_nand2_1 _16978_ (.Y(_10279_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][27] ),
    .B(net10114));
 sg13g2_o21ai_1 _16979_ (.B1(_10279_),
    .Y(_00837_),
    .A1(net9651),
    .A2(net10114));
 sg13g2_buf_16 clkbuf_leaf_150_clk (.X(clknet_leaf_150_clk),
    .A(clknet_8_28_0_clk));
 sg13g2_nand2_1 _16981_ (.Y(_10281_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][28] ),
    .B(net10114));
 sg13g2_o21ai_1 _16982_ (.B1(_10281_),
    .Y(_00838_),
    .A1(net9647),
    .A2(net10114));
 sg13g2_nand2_1 _16983_ (.Y(_10282_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][29] ),
    .B(net10112));
 sg13g2_o21ai_1 _16984_ (.B1(_10282_),
    .Y(_00839_),
    .A1(net9643),
    .A2(net10112));
 sg13g2_nand2_1 _16985_ (.Y(_10283_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][2] ),
    .B(net10109));
 sg13g2_o21ai_1 _16986_ (.B1(_10283_),
    .Y(_00840_),
    .A1(net10224),
    .A2(net10109));
 sg13g2_nand2_1 _16987_ (.Y(_10284_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][30] ),
    .B(net10112));
 sg13g2_o21ai_1 _16988_ (.B1(_10284_),
    .Y(_00841_),
    .A1(net9640),
    .A2(net10113));
 sg13g2_nand2_1 _16989_ (.Y(_10285_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][31] ),
    .B(net10111));
 sg13g2_o21ai_1 _16990_ (.B1(_10285_),
    .Y(_00842_),
    .A1(net9636),
    .A2(net10111));
 sg13g2_nand2_1 _16991_ (.Y(_10286_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][3] ),
    .B(net10108));
 sg13g2_o21ai_1 _16992_ (.B1(_10286_),
    .Y(_00843_),
    .A1(net10220),
    .A2(net10108));
 sg13g2_nand2_1 _16993_ (.Y(_10287_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][4] ),
    .B(net10115));
 sg13g2_o21ai_1 _16994_ (.B1(_10287_),
    .Y(_00844_),
    .A1(net10182),
    .A2(net10115));
 sg13g2_nand2_1 _16995_ (.Y(_10288_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][5] ),
    .B(net10109));
 sg13g2_o21ai_1 _16996_ (.B1(_10288_),
    .Y(_00845_),
    .A1(_10088_),
    .A2(net10109));
 sg13g2_nand2_1 _16997_ (.Y(_10289_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][6] ),
    .B(net10110));
 sg13g2_o21ai_1 _16998_ (.B1(_10289_),
    .Y(_00846_),
    .A1(net10171),
    .A2(net10110));
 sg13g2_nand2_1 _16999_ (.Y(_10290_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][7] ),
    .B(net10110));
 sg13g2_o21ai_1 _17000_ (.B1(_10290_),
    .Y(_00847_),
    .A1(net10167),
    .A2(net10110));
 sg13g2_nand2_1 _17001_ (.Y(_10291_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][8] ),
    .B(net10111));
 sg13g2_o21ai_1 _17002_ (.B1(_10291_),
    .Y(_00848_),
    .A1(net10127),
    .A2(net10111));
 sg13g2_nand2_1 _17003_ (.Y(_10292_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][9] ),
    .B(net10110));
 sg13g2_o21ai_1 _17004_ (.B1(_10292_),
    .Y(_00849_),
    .A1(net9974),
    .A2(net10110));
 sg13g2_nand2_1 _17005_ (.Y(_10293_),
    .A(_10124_),
    .B(_10167_));
 sg13g2_buf_16 clkbuf_leaf_147_clk (.X(clknet_leaf_147_clk),
    .A(clknet_8_96_0_clk));
 sg13g2_buf_2 place10606 (.A(_00086_),
    .X(net10606));
 sg13g2_buf_2 place10619 (.A(\u_ac_controller_soc_inst.cbus_addr[3] ),
    .X(net10619));
 sg13g2_nand2_1 _17009_ (.Y(_10297_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][0] ),
    .B(net9945));
 sg13g2_o21ai_1 _17010_ (.B1(_10297_),
    .Y(_00850_),
    .A1(net10278),
    .A2(net9945));
 sg13g2_nand2_1 _17011_ (.Y(_10298_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][10] ),
    .B(net9948));
 sg13g2_o21ai_1 _17012_ (.B1(_10298_),
    .Y(_00851_),
    .A1(net10131),
    .A2(net9948));
 sg13g2_nand2_1 _17013_ (.Y(_10299_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][11] ),
    .B(net9951));
 sg13g2_o21ai_1 _17014_ (.B1(_10299_),
    .Y(_00852_),
    .A1(net9985),
    .A2(net9951));
 sg13g2_nand2_1 _17015_ (.Y(_10300_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][12] ),
    .B(net9946));
 sg13g2_o21ai_1 _17016_ (.B1(_10300_),
    .Y(_00853_),
    .A1(net9800),
    .A2(net9946));
 sg13g2_nand2_1 _17017_ (.Y(_10301_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][13] ),
    .B(net9945));
 sg13g2_o21ai_1 _17018_ (.B1(_10301_),
    .Y(_00854_),
    .A1(net9978),
    .A2(net9945));
 sg13g2_nand2_1 _17019_ (.Y(_10302_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][14] ),
    .B(net9949));
 sg13g2_o21ai_1 _17020_ (.B1(_10302_),
    .Y(_00855_),
    .A1(net9798),
    .A2(net9949));
 sg13g2_nand2_1 _17021_ (.Y(_10303_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][15] ),
    .B(net9948));
 sg13g2_o21ai_1 _17022_ (.B1(_10303_),
    .Y(_00856_),
    .A1(net9791),
    .A2(net9948));
 sg13g2_nand2_1 _17023_ (.Y(_10304_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][16] ),
    .B(net9948));
 sg13g2_o21ai_1 _17024_ (.B1(_10304_),
    .Y(_00857_),
    .A1(net9744),
    .A2(net9948));
 sg13g2_buf_16 clkbuf_leaf_149_clk (.X(clknet_leaf_149_clk),
    .A(clknet_8_29_0_clk));
 sg13g2_nand2_1 _17026_ (.Y(_10306_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][17] ),
    .B(net9947));
 sg13g2_o21ai_1 _17027_ (.B1(_10306_),
    .Y(_00858_),
    .A1(net9742),
    .A2(net9947));
 sg13g2_nand2_1 _17028_ (.Y(_10307_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][18] ),
    .B(net9949));
 sg13g2_o21ai_1 _17029_ (.B1(_10307_),
    .Y(_00859_),
    .A1(net9738),
    .A2(net9949));
 sg13g2_buf_16 clkbuf_leaf_148_clk (.X(clknet_leaf_148_clk),
    .A(clknet_8_96_0_clk));
 sg13g2_nand2_1 _17031_ (.Y(_10309_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][19] ),
    .B(net9952));
 sg13g2_o21ai_1 _17032_ (.B1(_10309_),
    .Y(_00860_),
    .A1(net9723),
    .A2(net9952));
 sg13g2_nand2_1 _17033_ (.Y(_10310_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][1] ),
    .B(net9945));
 sg13g2_o21ai_1 _17034_ (.B1(_10310_),
    .Y(_00861_),
    .A1(net10227),
    .A2(net9945));
 sg13g2_nand2_1 _17035_ (.Y(_10311_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][20] ),
    .B(net9954));
 sg13g2_o21ai_1 _17036_ (.B1(_10311_),
    .Y(_00862_),
    .A1(net9719),
    .A2(net9954));
 sg13g2_nand2_1 _17037_ (.Y(_10312_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][21] ),
    .B(net9953));
 sg13g2_o21ai_1 _17038_ (.B1(_10312_),
    .Y(_00863_),
    .A1(net9712),
    .A2(net9953));
 sg13g2_nand2_1 _17039_ (.Y(_10313_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][22] ),
    .B(net9954));
 sg13g2_o21ai_1 _17040_ (.B1(_10313_),
    .Y(_00864_),
    .A1(net9695),
    .A2(net9954));
 sg13g2_nand2_1 _17041_ (.Y(_10314_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][23] ),
    .B(net9954));
 sg13g2_o21ai_1 _17042_ (.B1(_10314_),
    .Y(_00865_),
    .A1(net9692),
    .A2(net9954));
 sg13g2_nand2_1 _17043_ (.Y(_10315_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][24] ),
    .B(net9954));
 sg13g2_o21ai_1 _17044_ (.B1(_10315_),
    .Y(_00866_),
    .A1(net9687),
    .A2(net9954));
 sg13g2_nand2_1 _17045_ (.Y(_10316_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][25] ),
    .B(net9951));
 sg13g2_o21ai_1 _17046_ (.B1(_10316_),
    .Y(_00867_),
    .A1(net9680),
    .A2(net9951));
 sg13g2_buf_2 place10656 (.A(net10655),
    .X(net10656));
 sg13g2_nand2_1 _17048_ (.Y(_10318_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][26] ),
    .B(net9952));
 sg13g2_o21ai_1 _17049_ (.B1(_10318_),
    .Y(_00868_),
    .A1(net9675),
    .A2(net9952));
 sg13g2_nand2_1 _17050_ (.Y(_10319_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][27] ),
    .B(net9952));
 sg13g2_o21ai_1 _17051_ (.B1(_10319_),
    .Y(_00869_),
    .A1(_10023_),
    .A2(net9952));
 sg13g2_buf_2 place10643 (.A(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstr ),
    .X(net10643));
 sg13g2_nand2_1 _17053_ (.Y(_10321_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][28] ),
    .B(net9952));
 sg13g2_o21ai_1 _17054_ (.B1(_10321_),
    .Y(_00870_),
    .A1(net9647),
    .A2(net9952));
 sg13g2_nand2_1 _17055_ (.Y(_10322_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][29] ),
    .B(net9951));
 sg13g2_o21ai_1 _17056_ (.B1(_10322_),
    .Y(_00871_),
    .A1(_10041_),
    .A2(net9951));
 sg13g2_nand2_1 _17057_ (.Y(_10323_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][2] ),
    .B(net9947));
 sg13g2_o21ai_1 _17058_ (.B1(_10323_),
    .Y(_00872_),
    .A1(net10224),
    .A2(net9947));
 sg13g2_nand2_1 _17059_ (.Y(_10324_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][30] ),
    .B(net9950));
 sg13g2_o21ai_1 _17060_ (.B1(_10324_),
    .Y(_00873_),
    .A1(net9640),
    .A2(net9950));
 sg13g2_nand2_1 _17061_ (.Y(_10325_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][31] ),
    .B(net9950));
 sg13g2_o21ai_1 _17062_ (.B1(_10325_),
    .Y(_00874_),
    .A1(net9635),
    .A2(net9950));
 sg13g2_nand2_1 _17063_ (.Y(_10326_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][3] ),
    .B(net9948));
 sg13g2_o21ai_1 _17064_ (.B1(_10326_),
    .Y(_00875_),
    .A1(net10220),
    .A2(net9948));
 sg13g2_nand2_1 _17065_ (.Y(_10327_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][4] ),
    .B(net9953));
 sg13g2_o21ai_1 _17066_ (.B1(_10327_),
    .Y(_00876_),
    .A1(net10182),
    .A2(net9953));
 sg13g2_nand2_1 _17067_ (.Y(_10328_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][5] ),
    .B(net9947));
 sg13g2_o21ai_1 _17068_ (.B1(_10328_),
    .Y(_00877_),
    .A1(_10088_),
    .A2(net9947));
 sg13g2_nand2_1 _17069_ (.Y(_10329_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][6] ),
    .B(net9946));
 sg13g2_o21ai_1 _17070_ (.B1(_10329_),
    .Y(_00878_),
    .A1(net10170),
    .A2(net9946));
 sg13g2_nand2_1 _17071_ (.Y(_10330_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][7] ),
    .B(net9946));
 sg13g2_o21ai_1 _17072_ (.B1(_10330_),
    .Y(_00879_),
    .A1(net10167),
    .A2(net9946));
 sg13g2_nand2_1 _17073_ (.Y(_10331_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][8] ),
    .B(net9949));
 sg13g2_o21ai_1 _17074_ (.B1(_10331_),
    .Y(_00880_),
    .A1(_10111_),
    .A2(net9949));
 sg13g2_nand2_1 _17075_ (.Y(_10332_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][9] ),
    .B(net9946));
 sg13g2_o21ai_1 _17076_ (.B1(_10332_),
    .Y(_00881_),
    .A1(net9974),
    .A2(net9946));
 sg13g2_nand2b_2 _17077_ (.Y(_10333_),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_rd[4] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.latched_rd[3] ));
 sg13g2_nor2_2 _17078_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[2] ),
    .B(_10333_),
    .Y(_10334_));
 sg13g2_nand2_2 _17079_ (.Y(_10335_),
    .A(_10169_),
    .B(_10334_));
 sg13g2_buf_2 place10651 (.A(net10650),
    .X(net10651));
 sg13g2_buf_2 place10640 (.A(net10639),
    .X(net10640));
 sg13g2_buf_2 place10642 (.A(net10641),
    .X(net10642));
 sg13g2_nand2_1 _17083_ (.Y(_10339_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][0] ),
    .B(_10335_));
 sg13g2_o21ai_1 _17084_ (.B1(_10339_),
    .Y(_00882_),
    .A1(net10277),
    .A2(_10335_));
 sg13g2_nand2_1 _17085_ (.Y(_10340_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][10] ),
    .B(net10106));
 sg13g2_o21ai_1 _17086_ (.B1(_10340_),
    .Y(_00883_),
    .A1(net10133),
    .A2(net10106));
 sg13g2_nand2_1 _17087_ (.Y(_10341_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][11] ),
    .B(net10099));
 sg13g2_o21ai_1 _17088_ (.B1(_10341_),
    .Y(_00884_),
    .A1(net9982),
    .A2(net10099));
 sg13g2_nand2_1 _17089_ (.Y(_10342_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][12] ),
    .B(net10104));
 sg13g2_o21ai_1 _17090_ (.B1(_10342_),
    .Y(_00885_),
    .A1(net9802),
    .A2(net10104));
 sg13g2_nand2_1 _17091_ (.Y(_10343_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][13] ),
    .B(_10335_));
 sg13g2_o21ai_1 _17092_ (.B1(_10343_),
    .Y(_00886_),
    .A1(net9980),
    .A2(_10335_));
 sg13g2_nand2_1 _17093_ (.Y(_10344_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][14] ),
    .B(net10097));
 sg13g2_o21ai_1 _17094_ (.B1(_10344_),
    .Y(_00887_),
    .A1(net9797),
    .A2(net10097));
 sg13g2_nand2_1 _17095_ (.Y(_10345_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][15] ),
    .B(net10106));
 sg13g2_o21ai_1 _17096_ (.B1(_10345_),
    .Y(_00888_),
    .A1(net9793),
    .A2(net10106));
 sg13g2_nand2_1 _17097_ (.Y(_10346_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][16] ),
    .B(net10105));
 sg13g2_o21ai_1 _17098_ (.B1(_10346_),
    .Y(_00889_),
    .A1(net9744),
    .A2(net10105));
 sg13g2_buf_2 place10603 (.A(_00129_),
    .X(net10603));
 sg13g2_nand2_1 _17100_ (.Y(_10348_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][17] ),
    .B(net10103));
 sg13g2_o21ai_1 _17101_ (.B1(_10348_),
    .Y(_00890_),
    .A1(net9741),
    .A2(net10103));
 sg13g2_nand2_1 _17102_ (.Y(_10349_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][18] ),
    .B(net10098));
 sg13g2_o21ai_1 _17103_ (.B1(_10349_),
    .Y(_00891_),
    .A1(net9735),
    .A2(net10098));
 sg13g2_buf_2 place10636 (.A(net10634),
    .X(net10636));
 sg13g2_nand2_1 _17105_ (.Y(_10351_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][19] ),
    .B(net10102));
 sg13g2_o21ai_1 _17106_ (.B1(_10351_),
    .Y(_00892_),
    .A1(net9722),
    .A2(net10102));
 sg13g2_nand2_1 _17107_ (.Y(_10352_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][1] ),
    .B(net10103));
 sg13g2_o21ai_1 _17108_ (.B1(_10352_),
    .Y(_00893_),
    .A1(net10229),
    .A2(net10103));
 sg13g2_nand2_1 _17109_ (.Y(_10353_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][20] ),
    .B(net10098));
 sg13g2_o21ai_1 _17110_ (.B1(_10353_),
    .Y(_00894_),
    .A1(net9716),
    .A2(net10098));
 sg13g2_nand2_1 _17111_ (.Y(_10354_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][21] ),
    .B(net10098));
 sg13g2_o21ai_1 _17112_ (.B1(_10354_),
    .Y(_00895_),
    .A1(net9715),
    .A2(net10098));
 sg13g2_nand2_1 _17113_ (.Y(_10355_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][22] ),
    .B(net10099));
 sg13g2_o21ai_1 _17114_ (.B1(_10355_),
    .Y(_00896_),
    .A1(net9694),
    .A2(net10099));
 sg13g2_nand2_1 _17115_ (.Y(_10356_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][23] ),
    .B(net10099));
 sg13g2_o21ai_1 _17116_ (.B1(_10356_),
    .Y(_00897_),
    .A1(net9689),
    .A2(net10099));
 sg13g2_nand2_1 _17117_ (.Y(_10357_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][24] ),
    .B(net10099));
 sg13g2_o21ai_1 _17118_ (.B1(_10357_),
    .Y(_00898_),
    .A1(net9688),
    .A2(net10099));
 sg13g2_nand2_1 _17119_ (.Y(_10358_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][25] ),
    .B(net10100));
 sg13g2_o21ai_1 _17120_ (.B1(_10358_),
    .Y(_00899_),
    .A1(net9680),
    .A2(net10100));
 sg13g2_buf_2 place10632 (.A(\u_ac_controller_soc_inst.u_picorv32.is_slli_srli_srai ),
    .X(net10632));
 sg13g2_nand2_1 _17122_ (.Y(_10360_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][26] ),
    .B(net10101));
 sg13g2_o21ai_1 _17123_ (.B1(_10360_),
    .Y(_00900_),
    .A1(net9676),
    .A2(net10101));
 sg13g2_nand2_1 _17124_ (.Y(_10361_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][27] ),
    .B(net10100));
 sg13g2_o21ai_1 _17125_ (.B1(_10361_),
    .Y(_00901_),
    .A1(net9651),
    .A2(net10100));
 sg13g2_buf_2 place10658 (.A(net10657),
    .X(net10658));
 sg13g2_nand2_1 _17127_ (.Y(_10363_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][28] ),
    .B(net10102));
 sg13g2_o21ai_1 _17128_ (.B1(_10363_),
    .Y(_00902_),
    .A1(net9646),
    .A2(net10102));
 sg13g2_nand2_1 _17129_ (.Y(_10364_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][29] ),
    .B(net10100));
 sg13g2_o21ai_1 _17130_ (.B1(_10364_),
    .Y(_00903_),
    .A1(net9641),
    .A2(net10100));
 sg13g2_nand2_1 _17131_ (.Y(_10365_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][2] ),
    .B(net10103));
 sg13g2_o21ai_1 _17132_ (.B1(_10365_),
    .Y(_00904_),
    .A1(net10223),
    .A2(net10103));
 sg13g2_nand2_1 _17133_ (.Y(_10366_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][30] ),
    .B(net10101));
 sg13g2_o21ai_1 _17134_ (.B1(_10366_),
    .Y(_00905_),
    .A1(net9639),
    .A2(net10101));
 sg13g2_nand2_1 _17135_ (.Y(_10367_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][31] ),
    .B(net10102));
 sg13g2_o21ai_1 _17136_ (.B1(_10367_),
    .Y(_00906_),
    .A1(net9633),
    .A2(net10102));
 sg13g2_nand2_1 _17137_ (.Y(_10368_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][3] ),
    .B(net10105));
 sg13g2_o21ai_1 _17138_ (.B1(_10368_),
    .Y(_00907_),
    .A1(net10219),
    .A2(net10105));
 sg13g2_nand2_1 _17139_ (.Y(_10369_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][4] ),
    .B(net10105));
 sg13g2_o21ai_1 _17140_ (.B1(_10369_),
    .Y(_00908_),
    .A1(net10180),
    .A2(net10105));
 sg13g2_nand2_1 _17141_ (.Y(_10370_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][5] ),
    .B(net10106));
 sg13g2_o21ai_1 _17142_ (.B1(_10370_),
    .Y(_00909_),
    .A1(net10175),
    .A2(net10106));
 sg13g2_nand2_1 _17143_ (.Y(_10371_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][6] ),
    .B(net10104));
 sg13g2_o21ai_1 _17144_ (.B1(_10371_),
    .Y(_00910_),
    .A1(net10171),
    .A2(net10104));
 sg13g2_nand2_1 _17145_ (.Y(_10372_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][7] ),
    .B(net10104));
 sg13g2_o21ai_1 _17146_ (.B1(_10372_),
    .Y(_00911_),
    .A1(net10169),
    .A2(net10104));
 sg13g2_nand2_1 _17147_ (.Y(_10373_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][8] ),
    .B(net10097));
 sg13g2_o21ai_1 _17148_ (.B1(_10373_),
    .Y(_00912_),
    .A1(net10128),
    .A2(net10097));
 sg13g2_nand2_1 _17149_ (.Y(_10374_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][9] ),
    .B(net10104));
 sg13g2_o21ai_1 _17150_ (.B1(_10374_),
    .Y(_00913_),
    .A1(net9976),
    .A2(net10104));
 sg13g2_nand2_2 _17151_ (.Y(_10375_),
    .A(_10211_),
    .B(_10334_));
 sg13g2_buf_2 place10631 (.A(\u_ac_controller_soc_inst.u_picorv32.latched_stalu ),
    .X(net10631));
 sg13g2_buf_2 place10605 (.A(\u_ac_controller_soc_inst.cbus_wdata[0] ),
    .X(net10605));
 sg13g2_buf_2 place10596 (.A(net10595),
    .X(net10596));
 sg13g2_nand2_1 _17155_ (.Y(_10379_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][0] ),
    .B(_10375_));
 sg13g2_o21ai_1 _17156_ (.B1(_10379_),
    .Y(_00914_),
    .A1(net10278),
    .A2(_10375_));
 sg13g2_nand2_1 _17157_ (.Y(_10380_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][10] ),
    .B(net9938));
 sg13g2_o21ai_1 _17158_ (.B1(_10380_),
    .Y(_00915_),
    .A1(net10133),
    .A2(net9938));
 sg13g2_nand2_1 _17159_ (.Y(_10381_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][11] ),
    .B(net9942));
 sg13g2_o21ai_1 _17160_ (.B1(_10381_),
    .Y(_00916_),
    .A1(net9982),
    .A2(net9941));
 sg13g2_nand2_1 _17161_ (.Y(_10382_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][12] ),
    .B(net9939));
 sg13g2_o21ai_1 _17162_ (.B1(_10382_),
    .Y(_00917_),
    .A1(net9802),
    .A2(net9939));
 sg13g2_nand2_1 _17163_ (.Y(_10383_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][13] ),
    .B(net9936));
 sg13g2_o21ai_1 _17164_ (.B1(_10383_),
    .Y(_00918_),
    .A1(net9980),
    .A2(net9936));
 sg13g2_nand2_1 _17165_ (.Y(_10384_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][14] ),
    .B(_10375_));
 sg13g2_o21ai_1 _17166_ (.B1(_10384_),
    .Y(_00919_),
    .A1(net9797),
    .A2(_10375_));
 sg13g2_nand2_1 _17167_ (.Y(_10385_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][15] ),
    .B(net9938));
 sg13g2_o21ai_1 _17168_ (.B1(_10385_),
    .Y(_00920_),
    .A1(net9793),
    .A2(net9938));
 sg13g2_nand2_1 _17169_ (.Y(_10386_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][16] ),
    .B(net9937));
 sg13g2_o21ai_1 _17170_ (.B1(_10386_),
    .Y(_00921_),
    .A1(net9746),
    .A2(net9937));
 sg13g2_buf_2 place10595 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[0] ),
    .X(net10595));
 sg13g2_nand2_1 _17172_ (.Y(_10388_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][17] ),
    .B(net9936));
 sg13g2_o21ai_1 _17173_ (.B1(_10388_),
    .Y(_00922_),
    .A1(net9741),
    .A2(net9936));
 sg13g2_nand2_1 _17174_ (.Y(_10389_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][18] ),
    .B(net9940));
 sg13g2_o21ai_1 _17175_ (.B1(_10389_),
    .Y(_00923_),
    .A1(net9735),
    .A2(net9940));
 sg13g2_buf_2 place10613 (.A(\u_ac_controller_soc_inst.cbus_addr[7] ),
    .X(net10613));
 sg13g2_nand2_1 _17177_ (.Y(_10391_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][19] ),
    .B(net9944));
 sg13g2_o21ai_1 _17178_ (.B1(_10391_),
    .Y(_00924_),
    .A1(net9722),
    .A2(net9944));
 sg13g2_nand2_1 _17179_ (.Y(_10392_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][1] ),
    .B(net9936));
 sg13g2_o21ai_1 _17180_ (.B1(_10392_),
    .Y(_00925_),
    .A1(net10229),
    .A2(net9936));
 sg13g2_nand2_1 _17181_ (.Y(_10393_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][20] ),
    .B(net9940));
 sg13g2_o21ai_1 _17182_ (.B1(_10393_),
    .Y(_00926_),
    .A1(net9716),
    .A2(net9940));
 sg13g2_nand2_1 _17183_ (.Y(_10394_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][21] ),
    .B(net9940));
 sg13g2_o21ai_1 _17184_ (.B1(_10394_),
    .Y(_00927_),
    .A1(net9712),
    .A2(net9940));
 sg13g2_nand2_1 _17185_ (.Y(_10395_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][22] ),
    .B(net9941));
 sg13g2_o21ai_1 _17186_ (.B1(_10395_),
    .Y(_00928_),
    .A1(net9694),
    .A2(net9941));
 sg13g2_nand2_1 _17187_ (.Y(_10396_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][23] ),
    .B(net9941));
 sg13g2_o21ai_1 _17188_ (.B1(_10396_),
    .Y(_00929_),
    .A1(_09988_),
    .A2(net9941));
 sg13g2_nand2_1 _17189_ (.Y(_10397_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][24] ),
    .B(net9941));
 sg13g2_o21ai_1 _17190_ (.B1(_10397_),
    .Y(_00930_),
    .A1(net9688),
    .A2(net9941));
 sg13g2_nand2_1 _17191_ (.Y(_10398_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][25] ),
    .B(net9943));
 sg13g2_o21ai_1 _17192_ (.B1(_10398_),
    .Y(_00931_),
    .A1(_10005_),
    .A2(net9943));
 sg13g2_buf_2 place10593 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[10] ),
    .X(net10593));
 sg13g2_nand2_1 _17194_ (.Y(_10400_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][26] ),
    .B(net9942));
 sg13g2_o21ai_1 _17195_ (.B1(_10400_),
    .Y(_00932_),
    .A1(net9676),
    .A2(net9942));
 sg13g2_nand2_1 _17196_ (.Y(_10401_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][27] ),
    .B(net9943));
 sg13g2_o21ai_1 _17197_ (.B1(_10401_),
    .Y(_00933_),
    .A1(net9651),
    .A2(net9943));
 sg13g2_buf_2 place10594 (.A(net10593),
    .X(net10594));
 sg13g2_nand2_1 _17199_ (.Y(_10403_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][28] ),
    .B(net9944));
 sg13g2_o21ai_1 _17200_ (.B1(_10403_),
    .Y(_00934_),
    .A1(net9646),
    .A2(net9944));
 sg13g2_nand2_1 _17201_ (.Y(_10404_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][29] ),
    .B(net9943));
 sg13g2_o21ai_1 _17202_ (.B1(_10404_),
    .Y(_00935_),
    .A1(net9641),
    .A2(net9943));
 sg13g2_nand2_1 _17203_ (.Y(_10405_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][2] ),
    .B(net9938));
 sg13g2_o21ai_1 _17204_ (.B1(_10405_),
    .Y(_00936_),
    .A1(net10225),
    .A2(net9938));
 sg13g2_nand2_1 _17205_ (.Y(_10406_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][30] ),
    .B(net9944));
 sg13g2_o21ai_1 _17206_ (.B1(_10406_),
    .Y(_00937_),
    .A1(net9639),
    .A2(net9944));
 sg13g2_nand2_1 _17207_ (.Y(_10407_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][31] ),
    .B(net9944));
 sg13g2_o21ai_1 _17208_ (.B1(_10407_),
    .Y(_00938_),
    .A1(net9633),
    .A2(net9944));
 sg13g2_nand2_1 _17209_ (.Y(_10408_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][3] ),
    .B(net9937));
 sg13g2_o21ai_1 _17210_ (.B1(_10408_),
    .Y(_00939_),
    .A1(net10219),
    .A2(net9937));
 sg13g2_nand2_1 _17211_ (.Y(_10409_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][4] ),
    .B(net9937));
 sg13g2_o21ai_1 _17212_ (.B1(_10409_),
    .Y(_00940_),
    .A1(net10180),
    .A2(net9937));
 sg13g2_nand2_1 _17213_ (.Y(_10410_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][5] ),
    .B(net9938));
 sg13g2_o21ai_1 _17214_ (.B1(_10410_),
    .Y(_00941_),
    .A1(net10175),
    .A2(net9938));
 sg13g2_nand2_1 _17215_ (.Y(_10411_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][6] ),
    .B(net9939));
 sg13g2_o21ai_1 _17216_ (.B1(_10411_),
    .Y(_00942_),
    .A1(net10171),
    .A2(net9939));
 sg13g2_nand2_1 _17217_ (.Y(_10412_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][7] ),
    .B(net9939));
 sg13g2_o21ai_1 _17218_ (.B1(_10412_),
    .Y(_00943_),
    .A1(net10168),
    .A2(net9939));
 sg13g2_nand2_1 _17219_ (.Y(_10413_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][8] ),
    .B(net9940));
 sg13g2_o21ai_1 _17220_ (.B1(_10413_),
    .Y(_00944_),
    .A1(net10128),
    .A2(net9940));
 sg13g2_nand2_1 _17221_ (.Y(_10414_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][9] ),
    .B(net9939));
 sg13g2_o21ai_1 _17222_ (.B1(_10414_),
    .Y(_00945_),
    .A1(net9976),
    .A2(net9939));
 sg13g2_nand2_2 _17223_ (.Y(_10415_),
    .A(_09850_),
    .B(_10334_));
 sg13g2_buf_16 clkbuf_leaf_152_clk (.X(clknet_leaf_152_clk),
    .A(clknet_8_29_0_clk));
 sg13g2_buf_16 clkbuf_leaf_151_clk (.X(clknet_leaf_151_clk),
    .A(clknet_8_30_0_clk));
 sg13g2_buf_2 place10592 (.A(net10591),
    .X(net10592));
 sg13g2_nand2_1 _17227_ (.Y(_10419_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][0] ),
    .B(_10415_));
 sg13g2_o21ai_1 _17228_ (.B1(_10419_),
    .Y(_00946_),
    .A1(net10278),
    .A2(_10415_));
 sg13g2_nand2_1 _17229_ (.Y(_10420_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][10] ),
    .B(net10090));
 sg13g2_o21ai_1 _17230_ (.B1(_10420_),
    .Y(_00947_),
    .A1(net10133),
    .A2(net10090));
 sg13g2_nand2_1 _17231_ (.Y(_10421_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][11] ),
    .B(net10094));
 sg13g2_o21ai_1 _17232_ (.B1(_10421_),
    .Y(_00948_),
    .A1(net9982),
    .A2(net10094));
 sg13g2_nand2_1 _17233_ (.Y(_10422_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][12] ),
    .B(net10089));
 sg13g2_o21ai_1 _17234_ (.B1(_10422_),
    .Y(_00949_),
    .A1(net9802),
    .A2(net10089));
 sg13g2_nand2_1 _17235_ (.Y(_10423_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][13] ),
    .B(net10088));
 sg13g2_o21ai_1 _17236_ (.B1(_10423_),
    .Y(_00950_),
    .A1(net9981),
    .A2(net10088));
 sg13g2_nand2_1 _17237_ (.Y(_10424_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][14] ),
    .B(net10092));
 sg13g2_o21ai_1 _17238_ (.B1(_10424_),
    .Y(_00951_),
    .A1(net9797),
    .A2(net10092));
 sg13g2_nand2_1 _17239_ (.Y(_10425_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][15] ),
    .B(net10091));
 sg13g2_o21ai_1 _17240_ (.B1(_10425_),
    .Y(_00952_),
    .A1(net9793),
    .A2(net10091));
 sg13g2_nand2_1 _17241_ (.Y(_10426_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][16] ),
    .B(net10090));
 sg13g2_o21ai_1 _17242_ (.B1(_10426_),
    .Y(_00953_),
    .A1(net9744),
    .A2(net10090));
 sg13g2_buf_2 place10591 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[11] ),
    .X(net10591));
 sg13g2_nand2_1 _17244_ (.Y(_10428_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][17] ),
    .B(net10088));
 sg13g2_o21ai_1 _17245_ (.B1(_10428_),
    .Y(_00954_),
    .A1(net9741),
    .A2(net10088));
 sg13g2_nand2_1 _17246_ (.Y(_10429_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][18] ),
    .B(net10093));
 sg13g2_o21ai_1 _17247_ (.B1(_10429_),
    .Y(_00955_),
    .A1(net9735),
    .A2(net10093));
 sg13g2_buf_2 place10641 (.A(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh ),
    .X(net10641));
 sg13g2_nand2_1 _17249_ (.Y(_10431_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][19] ),
    .B(net10096));
 sg13g2_o21ai_1 _17250_ (.B1(_10431_),
    .Y(_00956_),
    .A1(net9722),
    .A2(net10096));
 sg13g2_nand2_1 _17251_ (.Y(_10432_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][1] ),
    .B(net10088));
 sg13g2_o21ai_1 _17252_ (.B1(_10432_),
    .Y(_00957_),
    .A1(net10228),
    .A2(net10088));
 sg13g2_nand2_1 _17253_ (.Y(_10433_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][20] ),
    .B(net10093));
 sg13g2_o21ai_1 _17254_ (.B1(_10433_),
    .Y(_00958_),
    .A1(net9716),
    .A2(net10093));
 sg13g2_nand2_1 _17255_ (.Y(_10434_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][21] ),
    .B(net10093));
 sg13g2_o21ai_1 _17256_ (.B1(_10434_),
    .Y(_00959_),
    .A1(net9712),
    .A2(net10093));
 sg13g2_nand2_1 _17257_ (.Y(_10435_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][22] ),
    .B(net10094));
 sg13g2_o21ai_1 _17258_ (.B1(_10435_),
    .Y(_00960_),
    .A1(net9694),
    .A2(net10094));
 sg13g2_nand2_1 _17259_ (.Y(_10436_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][23] ),
    .B(net10094));
 sg13g2_o21ai_1 _17260_ (.B1(_10436_),
    .Y(_00961_),
    .A1(_09988_),
    .A2(net10092));
 sg13g2_nand2_1 _17261_ (.Y(_10437_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][24] ),
    .B(net10094));
 sg13g2_o21ai_1 _17262_ (.B1(_10437_),
    .Y(_00962_),
    .A1(net9688),
    .A2(net10094));
 sg13g2_nand2_1 _17263_ (.Y(_10438_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][25] ),
    .B(net10095));
 sg13g2_o21ai_1 _17264_ (.B1(_10438_),
    .Y(_00963_),
    .A1(net9680),
    .A2(net10095));
 sg13g2_buf_2 place10589 (.A(net10588),
    .X(net10589));
 sg13g2_nand2_1 _17266_ (.Y(_10440_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][26] ),
    .B(net10095));
 sg13g2_o21ai_1 _17267_ (.B1(_10440_),
    .Y(_00964_),
    .A1(net9676),
    .A2(net10092));
 sg13g2_nand2_1 _17268_ (.Y(_10441_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][27] ),
    .B(net10095));
 sg13g2_o21ai_1 _17269_ (.B1(_10441_),
    .Y(_00965_),
    .A1(net9650),
    .A2(net10095));
 sg13g2_buf_2 place10588 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[12] ),
    .X(net10588));
 sg13g2_nand2_1 _17271_ (.Y(_10443_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][28] ),
    .B(net10096));
 sg13g2_o21ai_1 _17272_ (.B1(_10443_),
    .Y(_00966_),
    .A1(net9646),
    .A2(net10096));
 sg13g2_nand2_1 _17273_ (.Y(_10444_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][29] ),
    .B(net10095));
 sg13g2_o21ai_1 _17274_ (.B1(_10444_),
    .Y(_00967_),
    .A1(net9641),
    .A2(net10095));
 sg13g2_nand2_1 _17275_ (.Y(_10445_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][2] ),
    .B(net10091));
 sg13g2_o21ai_1 _17276_ (.B1(_10445_),
    .Y(_00968_),
    .A1(net10225),
    .A2(net10091));
 sg13g2_nand2_1 _17277_ (.Y(_10446_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][30] ),
    .B(net10096));
 sg13g2_o21ai_1 _17278_ (.B1(_10446_),
    .Y(_00969_),
    .A1(net9639),
    .A2(net10096));
 sg13g2_nand2_1 _17279_ (.Y(_10447_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][31] ),
    .B(net10096));
 sg13g2_o21ai_1 _17280_ (.B1(_10447_),
    .Y(_00970_),
    .A1(net9633),
    .A2(net10096));
 sg13g2_nand2_1 _17281_ (.Y(_10448_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][3] ),
    .B(net10091));
 sg13g2_o21ai_1 _17282_ (.B1(_10448_),
    .Y(_00971_),
    .A1(net10219),
    .A2(net10091));
 sg13g2_nand2_1 _17283_ (.Y(_10449_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][4] ),
    .B(net10090));
 sg13g2_o21ai_1 _17284_ (.B1(_10449_),
    .Y(_00972_),
    .A1(net10180),
    .A2(net10090));
 sg13g2_nand2_1 _17285_ (.Y(_10450_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][5] ),
    .B(net10091));
 sg13g2_o21ai_1 _17286_ (.B1(_10450_),
    .Y(_00973_),
    .A1(net10175),
    .A2(net10091));
 sg13g2_nand2_1 _17287_ (.Y(_10451_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][6] ),
    .B(net10089));
 sg13g2_o21ai_1 _17288_ (.B1(_10451_),
    .Y(_00974_),
    .A1(net10171),
    .A2(net10089));
 sg13g2_nand2_1 _17289_ (.Y(_10452_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][7] ),
    .B(net10089));
 sg13g2_o21ai_1 _17290_ (.B1(_10452_),
    .Y(_00975_),
    .A1(net10168),
    .A2(net10089));
 sg13g2_nand2_1 _17291_ (.Y(_10453_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][8] ),
    .B(net10093));
 sg13g2_o21ai_1 _17292_ (.B1(_10453_),
    .Y(_00976_),
    .A1(net10128),
    .A2(net10093));
 sg13g2_nand2_1 _17293_ (.Y(_10454_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][9] ),
    .B(net10089));
 sg13g2_o21ai_1 _17294_ (.B1(_10454_),
    .Y(_00977_),
    .A1(net9976),
    .A2(net10089));
 sg13g2_nand2_2 _17295_ (.Y(_10455_),
    .A(_10124_),
    .B(_10334_));
 sg13g2_buf_16 clkbuf_leaf_153_clk (.X(clknet_leaf_153_clk),
    .A(clknet_8_29_0_clk));
 sg13g2_buf_2 place10601 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[2] ),
    .X(net10601));
 sg13g2_buf_2 place10586 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[13] ),
    .X(net10586));
 sg13g2_nand2_1 _17299_ (.Y(_10459_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][0] ),
    .B(_10455_));
 sg13g2_o21ai_1 _17300_ (.B1(_10459_),
    .Y(_00978_),
    .A1(net10280),
    .A2(_10455_));
 sg13g2_nand2_1 _17301_ (.Y(_10460_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][10] ),
    .B(net9927));
 sg13g2_o21ai_1 _17302_ (.B1(_10460_),
    .Y(_00979_),
    .A1(net10133),
    .A2(net9927));
 sg13g2_nand2_1 _17303_ (.Y(_10461_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][11] ),
    .B(net9934));
 sg13g2_o21ai_1 _17304_ (.B1(_10461_),
    .Y(_00980_),
    .A1(_09877_),
    .A2(net9932));
 sg13g2_nand2_1 _17305_ (.Y(_10462_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][12] ),
    .B(net9929));
 sg13g2_o21ai_1 _17306_ (.B1(_10462_),
    .Y(_00981_),
    .A1(net9802),
    .A2(net9929));
 sg13g2_nand2_1 _17307_ (.Y(_10463_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][13] ),
    .B(net9926));
 sg13g2_o21ai_1 _17308_ (.B1(_10463_),
    .Y(_00982_),
    .A1(net9981),
    .A2(net9926));
 sg13g2_nand2_1 _17309_ (.Y(_10464_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][14] ),
    .B(net9932));
 sg13g2_o21ai_1 _17310_ (.B1(_10464_),
    .Y(_00983_),
    .A1(net9797),
    .A2(net9931));
 sg13g2_nand2_1 _17311_ (.Y(_10465_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][15] ),
    .B(net9928));
 sg13g2_o21ai_1 _17312_ (.B1(_10465_),
    .Y(_00984_),
    .A1(net9794),
    .A2(net9928));
 sg13g2_nand2_1 _17313_ (.Y(_10466_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][16] ),
    .B(_10455_));
 sg13g2_o21ai_1 _17314_ (.B1(_10466_),
    .Y(_00985_),
    .A1(net9744),
    .A2(_10455_));
 sg13g2_buf_16 clkbuf_leaf_154_clk (.X(clknet_leaf_154_clk),
    .A(clknet_8_31_0_clk));
 sg13g2_nand2_1 _17316_ (.Y(_10468_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][17] ),
    .B(net9926));
 sg13g2_o21ai_1 _17317_ (.B1(_10468_),
    .Y(_00986_),
    .A1(net9741),
    .A2(net9926));
 sg13g2_nand2_1 _17318_ (.Y(_10469_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][18] ),
    .B(net9931));
 sg13g2_o21ai_1 _17319_ (.B1(_10469_),
    .Y(_00987_),
    .A1(_09938_),
    .A2(net9931));
 sg13g2_buf_2 place10602 (.A(net10601),
    .X(net10602));
 sg13g2_nand2_1 _17321_ (.Y(_10471_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][19] ),
    .B(net9935));
 sg13g2_o21ai_1 _17322_ (.B1(_10471_),
    .Y(_00988_),
    .A1(net9722),
    .A2(net9935));
 sg13g2_nand2_1 _17323_ (.Y(_10472_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][1] ),
    .B(net9926));
 sg13g2_o21ai_1 _17324_ (.B1(_10472_),
    .Y(_00989_),
    .A1(net10229),
    .A2(net9926));
 sg13g2_nand2_1 _17325_ (.Y(_10473_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][20] ),
    .B(net9930));
 sg13g2_o21ai_1 _17326_ (.B1(_10473_),
    .Y(_00990_),
    .A1(net9716),
    .A2(net9930));
 sg13g2_nand2_1 _17327_ (.Y(_10474_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][21] ),
    .B(net9930));
 sg13g2_o21ai_1 _17328_ (.B1(_10474_),
    .Y(_00991_),
    .A1(net9712),
    .A2(net9930));
 sg13g2_nand2_1 _17329_ (.Y(_10475_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][22] ),
    .B(net9932));
 sg13g2_o21ai_1 _17330_ (.B1(_10475_),
    .Y(_00992_),
    .A1(net9694),
    .A2(net9932));
 sg13g2_nand2_1 _17331_ (.Y(_10476_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][23] ),
    .B(net9932));
 sg13g2_o21ai_1 _17332_ (.B1(_10476_),
    .Y(_00993_),
    .A1(_09988_),
    .A2(net9932));
 sg13g2_nand2_1 _17333_ (.Y(_10477_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][24] ),
    .B(net9932));
 sg13g2_o21ai_1 _17334_ (.B1(_10477_),
    .Y(_00994_),
    .A1(net9688),
    .A2(net9932));
 sg13g2_nand2_1 _17335_ (.Y(_10478_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][25] ),
    .B(net9934));
 sg13g2_o21ai_1 _17336_ (.B1(_10478_),
    .Y(_00995_),
    .A1(net9680),
    .A2(net9934));
 sg13g2_buf_2 place10585 (.A(net10584),
    .X(net10585));
 sg13g2_nand2_1 _17338_ (.Y(_10480_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][26] ),
    .B(net9934));
 sg13g2_o21ai_1 _17339_ (.B1(_10480_),
    .Y(_00996_),
    .A1(net9676),
    .A2(net9933));
 sg13g2_nand2_1 _17340_ (.Y(_10481_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][27] ),
    .B(net9934));
 sg13g2_o21ai_1 _17341_ (.B1(_10481_),
    .Y(_00997_),
    .A1(net9651),
    .A2(net9934));
 sg13g2_buf_16 clkbuf_leaf_161_clk (.X(clknet_leaf_161_clk),
    .A(clknet_8_74_0_clk));
 sg13g2_nand2_1 _17343_ (.Y(_10483_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][28] ),
    .B(net9935));
 sg13g2_o21ai_1 _17344_ (.B1(_10483_),
    .Y(_00998_),
    .A1(net9646),
    .A2(net9935));
 sg13g2_nand2_1 _17345_ (.Y(_10484_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][29] ),
    .B(net9934));
 sg13g2_o21ai_1 _17346_ (.B1(_10484_),
    .Y(_00999_),
    .A1(net9641),
    .A2(net9934));
 sg13g2_nand2_1 _17347_ (.Y(_10485_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][2] ),
    .B(net9928));
 sg13g2_o21ai_1 _17348_ (.B1(_10485_),
    .Y(_01000_),
    .A1(net10225),
    .A2(net9928));
 sg13g2_nand2_1 _17349_ (.Y(_10486_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][30] ),
    .B(net9935));
 sg13g2_o21ai_1 _17350_ (.B1(_10486_),
    .Y(_01001_),
    .A1(net9639),
    .A2(net9935));
 sg13g2_nand2_1 _17351_ (.Y(_10487_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][31] ),
    .B(net9935));
 sg13g2_o21ai_1 _17352_ (.B1(_10487_),
    .Y(_01002_),
    .A1(net9633),
    .A2(net9935));
 sg13g2_nand2_1 _17353_ (.Y(_10488_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][3] ),
    .B(net9927));
 sg13g2_o21ai_1 _17354_ (.B1(_10488_),
    .Y(_01003_),
    .A1(net10220),
    .A2(net9928));
 sg13g2_nand2_1 _17355_ (.Y(_10489_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][4] ),
    .B(net9927));
 sg13g2_o21ai_1 _17356_ (.B1(_10489_),
    .Y(_01004_),
    .A1(net10180),
    .A2(net9927));
 sg13g2_nand2_1 _17357_ (.Y(_10490_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][5] ),
    .B(net9928));
 sg13g2_o21ai_1 _17358_ (.B1(_10490_),
    .Y(_01005_),
    .A1(net10176),
    .A2(net9928));
 sg13g2_nand2_1 _17359_ (.Y(_10491_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][6] ),
    .B(net9929));
 sg13g2_o21ai_1 _17360_ (.B1(_10491_),
    .Y(_01006_),
    .A1(net10171),
    .A2(net9929));
 sg13g2_nand2_1 _17361_ (.Y(_10492_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][7] ),
    .B(net9929));
 sg13g2_o21ai_1 _17362_ (.B1(_10492_),
    .Y(_01007_),
    .A1(net10168),
    .A2(net9929));
 sg13g2_nand2_1 _17363_ (.Y(_10493_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][8] ),
    .B(net9931));
 sg13g2_o21ai_1 _17364_ (.B1(_10493_),
    .Y(_01008_),
    .A1(net10128),
    .A2(net9931));
 sg13g2_nand2_1 _17365_ (.Y(_10494_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][9] ),
    .B(net9929));
 sg13g2_o21ai_1 _17366_ (.B1(_10494_),
    .Y(_01009_),
    .A1(net9977),
    .A2(net9929));
 sg13g2_buf_16 clkbuf_leaf_160_clk (.X(clknet_leaf_160_clk),
    .A(clknet_8_74_0_clk));
 sg13g2_nand2_2 _17368_ (.Y(_10496_),
    .A(_10168_),
    .B(_10211_));
 sg13g2_buf_16 clkbuf_leaf_157_clk (.X(clknet_leaf_157_clk),
    .A(clknet_8_25_0_clk));
 sg13g2_buf_16 clkbuf_leaf_156_clk (.X(clknet_leaf_156_clk),
    .A(clknet_8_24_0_clk));
 sg13g2_buf_16 clkbuf_leaf_155_clk (.X(clknet_leaf_155_clk),
    .A(clknet_8_29_0_clk));
 sg13g2_nand2_1 _17372_ (.Y(_10500_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][0] ),
    .B(_10496_));
 sg13g2_o21ai_1 _17373_ (.B1(_10500_),
    .Y(_01010_),
    .A1(net10278),
    .A2(net9922));
 sg13g2_buf_2 place10590 (.A(net10588),
    .X(net10590));
 sg13g2_nand2_1 _17375_ (.Y(_10502_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][10] ),
    .B(net9921));
 sg13g2_o21ai_1 _17376_ (.B1(_10502_),
    .Y(_01011_),
    .A1(net10132),
    .A2(net9921));
 sg13g2_buf_2 place10583 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[15] ),
    .X(net10583));
 sg13g2_nand2_1 _17378_ (.Y(_10504_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][11] ),
    .B(net9917));
 sg13g2_o21ai_1 _17379_ (.B1(_10504_),
    .Y(_01012_),
    .A1(net9983),
    .A2(net9917));
 sg13g2_buf_16 clkbuf_leaf_158_clk (.X(clknet_leaf_158_clk),
    .A(clknet_8_25_0_clk));
 sg13g2_nand2_1 _17381_ (.Y(_10506_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][12] ),
    .B(net9925));
 sg13g2_o21ai_1 _17382_ (.B1(_10506_),
    .Y(_01013_),
    .A1(net9801),
    .A2(net9925));
 sg13g2_buf_2 place10587 (.A(net10586),
    .X(net10587));
 sg13g2_nand2_1 _17384_ (.Y(_10508_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][13] ),
    .B(net9922));
 sg13g2_o21ai_1 _17385_ (.B1(_10508_),
    .Y(_01014_),
    .A1(net9980),
    .A2(net9922));
 sg13g2_buf_2 place10604 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[1] ),
    .X(net10604));
 sg13g2_nand2_1 _17387_ (.Y(_10510_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][14] ),
    .B(net9916));
 sg13g2_o21ai_1 _17388_ (.B1(_10510_),
    .Y(_01015_),
    .A1(net9796),
    .A2(net9916));
 sg13g2_buf_2 place10630 (.A(\u_ac_controller_soc_inst.u_picorv32.latched_stalu ),
    .X(net10630));
 sg13g2_nand2_1 _17390_ (.Y(_10512_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][15] ),
    .B(net9923));
 sg13g2_o21ai_1 _17391_ (.B1(_10512_),
    .Y(_01016_),
    .A1(net9792),
    .A2(net9923));
 sg13g2_buf_2 place10580 (.A(net10579),
    .X(net10580));
 sg13g2_nand2_1 _17393_ (.Y(_10514_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][16] ),
    .B(net9924));
 sg13g2_o21ai_1 _17394_ (.B1(_10514_),
    .Y(_01017_),
    .A1(net9745),
    .A2(net9923));
 sg13g2_buf_2 place10579 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[16] ),
    .X(net10579));
 sg13g2_buf_2 place10645 (.A(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstr ),
    .X(net10645));
 sg13g2_nand2_1 _17397_ (.Y(_10517_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][17] ),
    .B(net9923));
 sg13g2_o21ai_1 _17398_ (.B1(_10517_),
    .Y(_01018_),
    .A1(net9739),
    .A2(net9923));
 sg13g2_buf_2 place10617 (.A(\u_ac_controller_soc_inst.cbus_addr[4] ),
    .X(net10617));
 sg13g2_nand2_1 _17400_ (.Y(_10519_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][18] ),
    .B(_10496_));
 sg13g2_o21ai_1 _17401_ (.B1(_10519_),
    .Y(_01019_),
    .A1(net9737),
    .A2(_10496_));
 sg13g2_buf_2 place10620 (.A(\u_ac_controller_soc_inst.cbus_addr[2] ),
    .X(net10620));
 sg13g2_buf_2 place10584 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[14] ),
    .X(net10584));
 sg13g2_nand2_1 _17404_ (.Y(_10522_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][19] ),
    .B(net9918));
 sg13g2_o21ai_1 _17405_ (.B1(_10522_),
    .Y(_01020_),
    .A1(net9721),
    .A2(net9918));
 sg13g2_buf_2 place10638 (.A(net10633),
    .X(net10638));
 sg13g2_nand2_1 _17407_ (.Y(_10524_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][1] ),
    .B(net9922));
 sg13g2_o21ai_1 _17408_ (.B1(_10524_),
    .Y(_01021_),
    .A1(net10229),
    .A2(net9922));
 sg13g2_buf_2 place10635 (.A(net10634),
    .X(net10635));
 sg13g2_nand2_1 _17410_ (.Y(_10526_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][20] ),
    .B(net9921));
 sg13g2_o21ai_1 _17411_ (.B1(_10526_),
    .Y(_01022_),
    .A1(net9720),
    .A2(net9921));
 sg13g2_buf_2 place10581 (.A(net10580),
    .X(net10581));
 sg13g2_nand2_1 _17413_ (.Y(_10528_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][21] ),
    .B(net9921));
 sg13g2_o21ai_1 _17414_ (.B1(_10528_),
    .Y(_01023_),
    .A1(net9715),
    .A2(net9921));
 sg13g2_buf_2 place10600 (.A(\u_ac_controller_soc_inst.cbus_wstrb[2] ),
    .X(net10600));
 sg13g2_nand2_1 _17416_ (.Y(_10530_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][22] ),
    .B(net9919));
 sg13g2_o21ai_1 _17417_ (.B1(_10530_),
    .Y(_01024_),
    .A1(_09980_),
    .A2(net9919));
 sg13g2_buf_16 clkbuf_leaf_163_clk (.X(clknet_leaf_163_clk),
    .A(clknet_8_97_0_clk));
 sg13g2_nand2_1 _17419_ (.Y(_10532_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][23] ),
    .B(net9917));
 sg13g2_o21ai_1 _17420_ (.B1(_10532_),
    .Y(_01025_),
    .A1(net9689),
    .A2(net9917));
 sg13g2_buf_16 clkbuf_leaf_162_clk (.X(clknet_leaf_162_clk),
    .A(clknet_8_96_0_clk));
 sg13g2_nand2_1 _17422_ (.Y(_10534_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][24] ),
    .B(net9919));
 sg13g2_o21ai_1 _17423_ (.B1(_10534_),
    .Y(_01026_),
    .A1(_09997_),
    .A2(net9919));
 sg13g2_buf_2 place10573 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[19] ),
    .X(net10573));
 sg13g2_nand2_1 _17425_ (.Y(_10536_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][25] ),
    .B(net9920));
 sg13g2_o21ai_1 _17426_ (.B1(_10536_),
    .Y(_01027_),
    .A1(net9681),
    .A2(net9920));
 sg13g2_buf_2 place10574 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[19] ),
    .X(net10574));
 sg13g2_buf_2 place10582 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[15] ),
    .X(net10582));
 sg13g2_nand2_1 _17429_ (.Y(_10539_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][26] ),
    .B(net9918));
 sg13g2_o21ai_1 _17430_ (.B1(_10539_),
    .Y(_01028_),
    .A1(net9674),
    .A2(net9918));
 sg13g2_buf_2 place10598 (.A(net10596),
    .X(net10598));
 sg13g2_nand2_1 _17432_ (.Y(_10541_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][27] ),
    .B(net9920));
 sg13g2_o21ai_1 _17433_ (.B1(_10541_),
    .Y(_01029_),
    .A1(net9652),
    .A2(net9920));
 sg13g2_buf_2 place10570 (.A(net10569),
    .X(net10570));
 sg13g2_buf_2 place10567 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[20] ),
    .X(net10567));
 sg13g2_nand2_1 _17436_ (.Y(_10544_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][28] ),
    .B(net9918));
 sg13g2_o21ai_1 _17437_ (.B1(_10544_),
    .Y(_01030_),
    .A1(_10033_),
    .A2(net9918));
 sg13g2_buf_2 place10568 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[1] ),
    .X(net10568));
 sg13g2_nand2_1 _17439_ (.Y(_10546_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][29] ),
    .B(net9920));
 sg13g2_o21ai_1 _17440_ (.B1(_10546_),
    .Y(_01031_),
    .A1(net9641),
    .A2(net9920));
 sg13g2_buf_2 place10569 (.A(net10568),
    .X(net10569));
 sg13g2_nand2_1 _17442_ (.Y(_10548_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][2] ),
    .B(net9923));
 sg13g2_o21ai_1 _17443_ (.B1(_10548_),
    .Y(_01032_),
    .A1(_10047_),
    .A2(net9923));
 sg13g2_buf_2 place10563 (.A(net10562),
    .X(net10563));
 sg13g2_nand2_1 _17445_ (.Y(_10550_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][30] ),
    .B(net9917));
 sg13g2_o21ai_1 _17446_ (.B1(_10550_),
    .Y(_01033_),
    .A1(_10056_),
    .A2(net9917));
 sg13g2_buf_2 place10566 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[20] ),
    .X(net10566));
 sg13g2_nand2_1 _17448_ (.Y(_10552_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][31] ),
    .B(net9918));
 sg13g2_o21ai_1 _17449_ (.B1(_10552_),
    .Y(_01034_),
    .A1(net9632),
    .A2(net9918));
 sg13g2_buf_2 place10564 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[21] ),
    .X(net10564));
 sg13g2_nand2_1 _17451_ (.Y(_10554_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][3] ),
    .B(net9924));
 sg13g2_o21ai_1 _17452_ (.B1(_10554_),
    .Y(_01035_),
    .A1(net10221),
    .A2(net9924));
 sg13g2_buf_2 place10560 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[22] ),
    .X(net10560));
 sg13g2_nand2_1 _17454_ (.Y(_10556_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][4] ),
    .B(net9921));
 sg13g2_o21ai_1 _17455_ (.B1(_10556_),
    .Y(_01036_),
    .A1(net10180),
    .A2(net9921));
 sg13g2_buf_2 place10561 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[22] ),
    .X(net10561));
 sg13g2_nand2_1 _17457_ (.Y(_10558_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][5] ),
    .B(net9924));
 sg13g2_o21ai_1 _17458_ (.B1(_10558_),
    .Y(_01037_),
    .A1(net10177),
    .A2(net9924));
 sg13g2_buf_16 clkbuf_leaf_164_clk (.X(clknet_leaf_164_clk),
    .A(clknet_8_97_0_clk));
 sg13g2_nand2_1 _17460_ (.Y(_10560_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][6] ),
    .B(net9925));
 sg13g2_o21ai_1 _17461_ (.B1(_10560_),
    .Y(_01038_),
    .A1(net10172),
    .A2(net9925));
 sg13g2_buf_2 place10559 (.A(net10558),
    .X(net10559));
 sg13g2_nand2_1 _17463_ (.Y(_10562_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][7] ),
    .B(net9925));
 sg13g2_o21ai_1 _17464_ (.B1(_10562_),
    .Y(_01039_),
    .A1(net10169),
    .A2(net9925));
 sg13g2_buf_2 place10558 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[23] ),
    .X(net10558));
 sg13g2_nand2_1 _17466_ (.Y(_10564_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][8] ),
    .B(net9916));
 sg13g2_o21ai_1 _17467_ (.B1(_10564_),
    .Y(_01040_),
    .A1(net10129),
    .A2(net9916));
 sg13g2_buf_16 clkbuf_leaf_170_clk (.X(clknet_leaf_170_clk),
    .A(clknet_8_79_0_clk));
 sg13g2_nand2_1 _17469_ (.Y(_10566_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][9] ),
    .B(net9925));
 sg13g2_o21ai_1 _17470_ (.B1(_10566_),
    .Y(_01041_),
    .A1(net9977),
    .A2(net9925));
 sg13g2_nor2_2 _17471_ (.A(_00084_),
    .B(_10333_),
    .Y(_10567_));
 sg13g2_nand2_2 _17472_ (.Y(_10568_),
    .A(_10169_),
    .B(_10567_));
 sg13g2_buf_16 clkbuf_leaf_166_clk (.X(clknet_leaf_166_clk),
    .A(clknet_8_75_0_clk));
 sg13g2_buf_2 place10554 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[24] ),
    .X(net10554));
 sg13g2_buf_2 place10556 (.A(net10555),
    .X(net10556));
 sg13g2_nand2_1 _17476_ (.Y(_10572_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][0] ),
    .B(_10568_));
 sg13g2_o21ai_1 _17477_ (.B1(_10572_),
    .Y(_01042_),
    .A1(net10280),
    .A2(_10568_));
 sg13g2_nand2_1 _17478_ (.Y(_10573_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][10] ),
    .B(net10086));
 sg13g2_o21ai_1 _17479_ (.B1(_10573_),
    .Y(_01043_),
    .A1(net10132),
    .A2(net10086));
 sg13g2_nand2_1 _17480_ (.Y(_10574_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][11] ),
    .B(net10083));
 sg13g2_o21ai_1 _17481_ (.B1(_10574_),
    .Y(_01044_),
    .A1(net9983),
    .A2(net10083));
 sg13g2_nand2_1 _17482_ (.Y(_10575_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][12] ),
    .B(net10084));
 sg13g2_o21ai_1 _17483_ (.B1(_10575_),
    .Y(_01045_),
    .A1(_09885_),
    .A2(net10084));
 sg13g2_nand2_1 _17484_ (.Y(_10576_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][13] ),
    .B(net10084));
 sg13g2_o21ai_1 _17485_ (.B1(_10576_),
    .Y(_01046_),
    .A1(net9980),
    .A2(net10084));
 sg13g2_nand2_1 _17486_ (.Y(_10577_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][14] ),
    .B(net10079));
 sg13g2_o21ai_1 _17487_ (.B1(_10577_),
    .Y(_01047_),
    .A1(net9797),
    .A2(net10079));
 sg13g2_nand2_1 _17488_ (.Y(_10578_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][15] ),
    .B(net10087));
 sg13g2_o21ai_1 _17489_ (.B1(_10578_),
    .Y(_01048_),
    .A1(net9793),
    .A2(net10087));
 sg13g2_nand2_1 _17490_ (.Y(_10579_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][16] ),
    .B(_10568_));
 sg13g2_o21ai_1 _17491_ (.B1(_10579_),
    .Y(_01049_),
    .A1(net9746),
    .A2(_10568_));
 sg13g2_buf_16 clkbuf_leaf_172_clk (.X(clknet_leaf_172_clk),
    .A(clknet_8_90_0_clk));
 sg13g2_nand2_1 _17493_ (.Y(_10581_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][17] ),
    .B(net10084));
 sg13g2_o21ai_1 _17494_ (.B1(_10581_),
    .Y(_01050_),
    .A1(net9741),
    .A2(net10085));
 sg13g2_nand2_1 _17495_ (.Y(_10582_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][18] ),
    .B(net10081));
 sg13g2_o21ai_1 _17496_ (.B1(_10582_),
    .Y(_01051_),
    .A1(net9735),
    .A2(net10081));
 sg13g2_buf_2 place10553 (.A(net10552),
    .X(net10553));
 sg13g2_nand2_1 _17498_ (.Y(_10584_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][19] ),
    .B(net10080));
 sg13g2_o21ai_1 _17499_ (.B1(_10584_),
    .Y(_01052_),
    .A1(_09947_),
    .A2(net10080));
 sg13g2_nand2_1 _17500_ (.Y(_10585_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][1] ),
    .B(net10084));
 sg13g2_o21ai_1 _17501_ (.B1(_10585_),
    .Y(_01053_),
    .A1(net10226),
    .A2(net10084));
 sg13g2_nand2_1 _17502_ (.Y(_10586_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][20] ),
    .B(net10081));
 sg13g2_o21ai_1 _17503_ (.B1(_10586_),
    .Y(_01054_),
    .A1(net9716),
    .A2(net10081));
 sg13g2_nand2_1 _17504_ (.Y(_10587_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][21] ),
    .B(net10082));
 sg13g2_o21ai_1 _17505_ (.B1(_10587_),
    .Y(_01055_),
    .A1(_09972_),
    .A2(net10081));
 sg13g2_nand2_1 _17506_ (.Y(_10588_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][22] ),
    .B(net10082));
 sg13g2_o21ai_1 _17507_ (.B1(_10588_),
    .Y(_01056_),
    .A1(net9696),
    .A2(net10082));
 sg13g2_nand2_1 _17508_ (.Y(_10589_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][23] ),
    .B(net10082));
 sg13g2_o21ai_1 _17509_ (.B1(_10589_),
    .Y(_01057_),
    .A1(net9690),
    .A2(net10082));
 sg13g2_nand2_1 _17510_ (.Y(_10590_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][24] ),
    .B(net10081));
 sg13g2_o21ai_1 _17511_ (.B1(_10590_),
    .Y(_01058_),
    .A1(net9684),
    .A2(net10082));
 sg13g2_nand2_1 _17512_ (.Y(_10591_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][25] ),
    .B(net10083));
 sg13g2_o21ai_1 _17513_ (.B1(_10591_),
    .Y(_01059_),
    .A1(net9681),
    .A2(net10083));
 sg13g2_buf_2 place10557 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[23] ),
    .X(net10557));
 sg13g2_nand2_1 _17515_ (.Y(_10593_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][26] ),
    .B(net10080));
 sg13g2_o21ai_1 _17516_ (.B1(_10593_),
    .Y(_01060_),
    .A1(net9674),
    .A2(net10080));
 sg13g2_nand2_1 _17517_ (.Y(_10594_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][27] ),
    .B(net10083));
 sg13g2_o21ai_1 _17518_ (.B1(_10594_),
    .Y(_01061_),
    .A1(net9652),
    .A2(net10083));
 sg13g2_buf_2 place10552 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[25] ),
    .X(net10552));
 sg13g2_nand2_1 _17520_ (.Y(_10596_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][28] ),
    .B(net10080));
 sg13g2_o21ai_1 _17521_ (.B1(_10596_),
    .Y(_01062_),
    .A1(_10033_),
    .A2(net10080));
 sg13g2_nand2_1 _17522_ (.Y(_10597_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][29] ),
    .B(net10083));
 sg13g2_o21ai_1 _17523_ (.B1(_10597_),
    .Y(_01063_),
    .A1(net9641),
    .A2(net10083));
 sg13g2_nand2_1 _17524_ (.Y(_10598_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][2] ),
    .B(net10087));
 sg13g2_o21ai_1 _17525_ (.B1(_10598_),
    .Y(_01064_),
    .A1(net10225),
    .A2(net10087));
 sg13g2_nand2_1 _17526_ (.Y(_10599_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][30] ),
    .B(net10079));
 sg13g2_o21ai_1 _17527_ (.B1(_10599_),
    .Y(_01065_),
    .A1(net9637),
    .A2(net10079));
 sg13g2_nand2_1 _17528_ (.Y(_10600_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][31] ),
    .B(net10080));
 sg13g2_o21ai_1 _17529_ (.B1(_10600_),
    .Y(_01066_),
    .A1(net9632),
    .A2(net10080));
 sg13g2_nand2_1 _17530_ (.Y(_10601_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][3] ),
    .B(net10086));
 sg13g2_o21ai_1 _17531_ (.B1(_10601_),
    .Y(_01067_),
    .A1(net10219),
    .A2(_10568_));
 sg13g2_nand2_1 _17532_ (.Y(_10602_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][4] ),
    .B(net10086));
 sg13g2_o21ai_1 _17533_ (.B1(_10602_),
    .Y(_01068_),
    .A1(net10179),
    .A2(net10086));
 sg13g2_nand2_1 _17534_ (.Y(_10603_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][5] ),
    .B(net10087));
 sg13g2_o21ai_1 _17535_ (.B1(_10603_),
    .Y(_01069_),
    .A1(net10176),
    .A2(net10087));
 sg13g2_nand2_1 _17536_ (.Y(_10604_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][6] ),
    .B(net10085));
 sg13g2_o21ai_1 _17537_ (.B1(_10604_),
    .Y(_01070_),
    .A1(net10173),
    .A2(net10085));
 sg13g2_nand2_1 _17538_ (.Y(_10605_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][7] ),
    .B(net10085));
 sg13g2_o21ai_1 _17539_ (.B1(_10605_),
    .Y(_01071_),
    .A1(net10168),
    .A2(net10085));
 sg13g2_nand2_1 _17540_ (.Y(_10606_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][8] ),
    .B(net10079));
 sg13g2_o21ai_1 _17541_ (.B1(_10606_),
    .Y(_01072_),
    .A1(net10129),
    .A2(net10079));
 sg13g2_nand2_1 _17542_ (.Y(_10607_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][9] ),
    .B(net10085));
 sg13g2_o21ai_1 _17543_ (.B1(_10607_),
    .Y(_01073_),
    .A1(net9977),
    .A2(net10085));
 sg13g2_nand2_2 _17544_ (.Y(_10608_),
    .A(_10211_),
    .B(_10567_));
 sg13g2_buf_2 place10548 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[26] ),
    .X(net10548));
 sg13g2_buf_2 place10555 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[24] ),
    .X(net10555));
 sg13g2_buf_2 place10549 (.A(net10548),
    .X(net10549));
 sg13g2_nand2_1 _17548_ (.Y(_10612_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][0] ),
    .B(_10608_));
 sg13g2_o21ai_1 _17549_ (.B1(_10612_),
    .Y(_01074_),
    .A1(net10280),
    .A2(net9907));
 sg13g2_nand2_1 _17550_ (.Y(_10613_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][10] ),
    .B(net9908));
 sg13g2_o21ai_1 _17551_ (.B1(_10613_),
    .Y(_01075_),
    .A1(net10132),
    .A2(net9908));
 sg13g2_nand2_1 _17552_ (.Y(_10614_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][11] ),
    .B(net9913));
 sg13g2_o21ai_1 _17553_ (.B1(_10614_),
    .Y(_01076_),
    .A1(net9983),
    .A2(net9913));
 sg13g2_nand2_1 _17554_ (.Y(_10615_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][12] ),
    .B(net9909));
 sg13g2_o21ai_1 _17555_ (.B1(_10615_),
    .Y(_01077_),
    .A1(net9799),
    .A2(net9909));
 sg13g2_nand2_1 _17556_ (.Y(_10616_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][13] ),
    .B(net9909));
 sg13g2_o21ai_1 _17557_ (.B1(_10616_),
    .Y(_01078_),
    .A1(net9980),
    .A2(net9909));
 sg13g2_nand2_1 _17558_ (.Y(_10617_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][14] ),
    .B(net9914));
 sg13g2_o21ai_1 _17559_ (.B1(_10617_),
    .Y(_01079_),
    .A1(net9797),
    .A2(net9914));
 sg13g2_nand2_1 _17560_ (.Y(_10618_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][15] ),
    .B(net9908));
 sg13g2_o21ai_1 _17561_ (.B1(_10618_),
    .Y(_01080_),
    .A1(net9794),
    .A2(net9908));
 sg13g2_nand2_1 _17562_ (.Y(_10619_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][16] ),
    .B(net9907));
 sg13g2_o21ai_1 _17563_ (.B1(_10619_),
    .Y(_01081_),
    .A1(net9746),
    .A2(net9907));
 sg13g2_buf_2 place10551 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[25] ),
    .X(net10551));
 sg13g2_nand2_1 _17565_ (.Y(_10621_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][17] ),
    .B(net9909));
 sg13g2_o21ai_1 _17566_ (.B1(_10621_),
    .Y(_01082_),
    .A1(net9741),
    .A2(net9910));
 sg13g2_nand2_1 _17567_ (.Y(_10622_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][18] ),
    .B(net9911));
 sg13g2_o21ai_1 _17568_ (.B1(_10622_),
    .Y(_01083_),
    .A1(net9735),
    .A2(net9911));
 sg13g2_buf_2 place10546 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[27] ),
    .X(net10546));
 sg13g2_nand2_1 _17570_ (.Y(_10624_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][19] ),
    .B(net9915));
 sg13g2_o21ai_1 _17571_ (.B1(_10624_),
    .Y(_01084_),
    .A1(_09947_),
    .A2(net9915));
 sg13g2_nand2_1 _17572_ (.Y(_10625_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][1] ),
    .B(net9909));
 sg13g2_o21ai_1 _17573_ (.B1(_10625_),
    .Y(_01085_),
    .A1(_09954_),
    .A2(net9909));
 sg13g2_nand2_1 _17574_ (.Y(_10626_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][20] ),
    .B(net9911));
 sg13g2_o21ai_1 _17575_ (.B1(_10626_),
    .Y(_01086_),
    .A1(_09963_),
    .A2(net9911));
 sg13g2_nand2_1 _17576_ (.Y(_10627_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][21] ),
    .B(net9911));
 sg13g2_o21ai_1 _17577_ (.B1(_10627_),
    .Y(_01087_),
    .A1(_09972_),
    .A2(net9911));
 sg13g2_nand2_1 _17578_ (.Y(_10628_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][22] ),
    .B(net9912));
 sg13g2_o21ai_1 _17579_ (.B1(_10628_),
    .Y(_01088_),
    .A1(net9696),
    .A2(net9912));
 sg13g2_nand2_1 _17580_ (.Y(_10629_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][23] ),
    .B(net9912));
 sg13g2_o21ai_1 _17581_ (.B1(_10629_),
    .Y(_01089_),
    .A1(net9690),
    .A2(net9912));
 sg13g2_nand2_1 _17582_ (.Y(_10630_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][24] ),
    .B(net9912));
 sg13g2_o21ai_1 _17583_ (.B1(_10630_),
    .Y(_01090_),
    .A1(net9684),
    .A2(net9912));
 sg13g2_nand2_1 _17584_ (.Y(_10631_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][25] ),
    .B(net9913));
 sg13g2_o21ai_1 _17585_ (.B1(_10631_),
    .Y(_01091_),
    .A1(net9681),
    .A2(net9913));
 sg13g2_buf_16 clkbuf_leaf_173_clk (.X(clknet_leaf_173_clk),
    .A(clknet_8_88_0_clk));
 sg13g2_nand2_1 _17587_ (.Y(_10633_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][26] ),
    .B(net9915));
 sg13g2_o21ai_1 _17588_ (.B1(_10633_),
    .Y(_01092_),
    .A1(_10014_),
    .A2(net9915));
 sg13g2_nand2_1 _17589_ (.Y(_10634_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][27] ),
    .B(net9913));
 sg13g2_o21ai_1 _17590_ (.B1(_10634_),
    .Y(_01093_),
    .A1(net9652),
    .A2(net9913));
 sg13g2_buf_2 place10547 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[27] ),
    .X(net10547));
 sg13g2_nand2_1 _17592_ (.Y(_10636_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][28] ),
    .B(net9915));
 sg13g2_o21ai_1 _17593_ (.B1(_10636_),
    .Y(_01094_),
    .A1(_10033_),
    .A2(net9915));
 sg13g2_nand2_1 _17594_ (.Y(_10637_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][29] ),
    .B(net9913));
 sg13g2_o21ai_1 _17595_ (.B1(_10637_),
    .Y(_01095_),
    .A1(net9642),
    .A2(net9913));
 sg13g2_nand2_1 _17596_ (.Y(_10638_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][2] ),
    .B(net9908));
 sg13g2_o21ai_1 _17597_ (.B1(_10638_),
    .Y(_01096_),
    .A1(net10225),
    .A2(net9908));
 sg13g2_nand2_1 _17598_ (.Y(_10639_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][30] ),
    .B(net9914));
 sg13g2_o21ai_1 _17599_ (.B1(_10639_),
    .Y(_01097_),
    .A1(net9637),
    .A2(net9914));
 sg13g2_nand2_1 _17600_ (.Y(_10640_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][31] ),
    .B(net9915));
 sg13g2_o21ai_1 _17601_ (.B1(_10640_),
    .Y(_01098_),
    .A1(net9632),
    .A2(net9915));
 sg13g2_nand2_1 _17602_ (.Y(_10641_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][3] ),
    .B(net9907));
 sg13g2_o21ai_1 _17603_ (.B1(_10641_),
    .Y(_01099_),
    .A1(net10219),
    .A2(net9907));
 sg13g2_nand2_1 _17604_ (.Y(_10642_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][4] ),
    .B(net9907));
 sg13g2_o21ai_1 _17605_ (.B1(_10642_),
    .Y(_01100_),
    .A1(net10179),
    .A2(net9907));
 sg13g2_nand2_1 _17606_ (.Y(_10643_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][5] ),
    .B(net9908));
 sg13g2_o21ai_1 _17607_ (.B1(_10643_),
    .Y(_01101_),
    .A1(net10176),
    .A2(net9908));
 sg13g2_nand2_1 _17608_ (.Y(_10644_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][6] ),
    .B(net9910));
 sg13g2_o21ai_1 _17609_ (.B1(_10644_),
    .Y(_01102_),
    .A1(net10173),
    .A2(net9910));
 sg13g2_nand2_1 _17610_ (.Y(_10645_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][7] ),
    .B(net9910));
 sg13g2_o21ai_1 _17611_ (.B1(_10645_),
    .Y(_01103_),
    .A1(net10168),
    .A2(net9910));
 sg13g2_nand2_1 _17612_ (.Y(_10646_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][8] ),
    .B(net9914));
 sg13g2_o21ai_1 _17613_ (.B1(_10646_),
    .Y(_01104_),
    .A1(net10129),
    .A2(net9911));
 sg13g2_nand2_1 _17614_ (.Y(_10647_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][9] ),
    .B(net9910));
 sg13g2_o21ai_1 _17615_ (.B1(_10647_),
    .Y(_01105_),
    .A1(net9977),
    .A2(net9910));
 sg13g2_nand2_2 _17616_ (.Y(_10648_),
    .A(_09850_),
    .B(_10567_));
 sg13g2_buf_2 place10550 (.A(net10549),
    .X(net10550));
 sg13g2_buf_16 clkbuf_leaf_174_clk (.X(clknet_leaf_174_clk),
    .A(clknet_8_88_0_clk));
 sg13g2_buf_2 place10543 (.A(net10542),
    .X(net10543));
 sg13g2_nand2_1 _17620_ (.Y(_10652_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][0] ),
    .B(net10074));
 sg13g2_o21ai_1 _17621_ (.B1(_10652_),
    .Y(_01106_),
    .A1(net10280),
    .A2(net10074));
 sg13g2_nand2_1 _17622_ (.Y(_10653_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][10] ),
    .B(net10078));
 sg13g2_o21ai_1 _17623_ (.B1(_10653_),
    .Y(_01107_),
    .A1(net10132),
    .A2(net10078));
 sg13g2_nand2_1 _17624_ (.Y(_10654_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][11] ),
    .B(net10071));
 sg13g2_o21ai_1 _17625_ (.B1(_10654_),
    .Y(_01108_),
    .A1(net9983),
    .A2(net10071));
 sg13g2_nand2_1 _17626_ (.Y(_10655_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][12] ),
    .B(net10075));
 sg13g2_o21ai_1 _17627_ (.B1(_10655_),
    .Y(_01109_),
    .A1(net9799),
    .A2(net10075));
 sg13g2_nand2_1 _17628_ (.Y(_10656_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][13] ),
    .B(net10075));
 sg13g2_o21ai_1 _17629_ (.B1(_10656_),
    .Y(_01110_),
    .A1(net9980),
    .A2(net10076));
 sg13g2_nand2_1 _17630_ (.Y(_10657_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][14] ),
    .B(net10072));
 sg13g2_o21ai_1 _17631_ (.B1(_10657_),
    .Y(_01111_),
    .A1(net9797),
    .A2(net10072));
 sg13g2_nand2_1 _17632_ (.Y(_10658_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][15] ),
    .B(net10078));
 sg13g2_o21ai_1 _17633_ (.B1(_10658_),
    .Y(_01112_),
    .A1(net9794),
    .A2(net10078));
 sg13g2_nand2_1 _17634_ (.Y(_10659_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][16] ),
    .B(net10074));
 sg13g2_o21ai_1 _17635_ (.B1(_10659_),
    .Y(_01113_),
    .A1(net9743),
    .A2(net10074));
 sg13g2_buf_2 place10544 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[28] ),
    .X(net10544));
 sg13g2_nand2_1 _17637_ (.Y(_10661_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][17] ),
    .B(net10076));
 sg13g2_o21ai_1 _17638_ (.B1(_10661_),
    .Y(_01114_),
    .A1(net9739),
    .A2(net10075));
 sg13g2_nand2_1 _17639_ (.Y(_10662_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][18] ),
    .B(net10069));
 sg13g2_o21ai_1 _17640_ (.B1(_10662_),
    .Y(_01115_),
    .A1(_09938_),
    .A2(net10069));
 sg13g2_buf_16 clkbuf_leaf_176_clk (.X(clknet_leaf_176_clk),
    .A(clknet_8_78_0_clk));
 sg13g2_nand2_1 _17642_ (.Y(_10664_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][19] ),
    .B(net10073));
 sg13g2_o21ai_1 _17643_ (.B1(_10664_),
    .Y(_01116_),
    .A1(_09947_),
    .A2(net10073));
 sg13g2_nand2_1 _17644_ (.Y(_10665_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][1] ),
    .B(net10075));
 sg13g2_o21ai_1 _17645_ (.B1(_10665_),
    .Y(_01117_),
    .A1(net10226),
    .A2(net10075));
 sg13g2_nand2_1 _17646_ (.Y(_10666_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][20] ),
    .B(net10069));
 sg13g2_o21ai_1 _17647_ (.B1(_10666_),
    .Y(_01118_),
    .A1(_09963_),
    .A2(net10069));
 sg13g2_nand2_1 _17648_ (.Y(_10667_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][21] ),
    .B(net10069));
 sg13g2_o21ai_1 _17649_ (.B1(_10667_),
    .Y(_01119_),
    .A1(_09972_),
    .A2(net10069));
 sg13g2_nand2_1 _17650_ (.Y(_10668_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][22] ),
    .B(net10070));
 sg13g2_o21ai_1 _17651_ (.B1(_10668_),
    .Y(_01120_),
    .A1(net9693),
    .A2(net10070));
 sg13g2_nand2_1 _17652_ (.Y(_10669_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][23] ),
    .B(net10070));
 sg13g2_o21ai_1 _17653_ (.B1(_10669_),
    .Y(_01121_),
    .A1(net9690),
    .A2(net10069));
 sg13g2_nand2_1 _17654_ (.Y(_10670_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][24] ),
    .B(net10070));
 sg13g2_o21ai_1 _17655_ (.B1(_10670_),
    .Y(_01122_),
    .A1(net9684),
    .A2(net10070));
 sg13g2_nand2_1 _17656_ (.Y(_10671_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][25] ),
    .B(net10071));
 sg13g2_o21ai_1 _17657_ (.B1(_10671_),
    .Y(_01123_),
    .A1(net9681),
    .A2(net10071));
 sg13g2_buf_2 place10539 (.A(net10538),
    .X(net10539));
 sg13g2_nand2_1 _17659_ (.Y(_10673_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][26] ),
    .B(net10073));
 sg13g2_o21ai_1 _17660_ (.B1(_10673_),
    .Y(_01124_),
    .A1(_10014_),
    .A2(net10073));
 sg13g2_nand2_1 _17661_ (.Y(_10674_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][27] ),
    .B(net10071));
 sg13g2_o21ai_1 _17662_ (.B1(_10674_),
    .Y(_01125_),
    .A1(net9652),
    .A2(net10071));
 sg13g2_buf_16 clkbuf_leaf_177_clk (.X(clknet_leaf_177_clk),
    .A(clknet_8_78_0_clk));
 sg13g2_nand2_1 _17664_ (.Y(_10676_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][28] ),
    .B(net10073));
 sg13g2_o21ai_1 _17665_ (.B1(_10676_),
    .Y(_01126_),
    .A1(_10033_),
    .A2(net10073));
 sg13g2_nand2_1 _17666_ (.Y(_10677_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][29] ),
    .B(net10071));
 sg13g2_o21ai_1 _17667_ (.B1(_10677_),
    .Y(_01127_),
    .A1(net9642),
    .A2(net10071));
 sg13g2_nand2_1 _17668_ (.Y(_10678_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][2] ),
    .B(net10078));
 sg13g2_o21ai_1 _17669_ (.B1(_10678_),
    .Y(_01128_),
    .A1(net10225),
    .A2(net10078));
 sg13g2_nand2_1 _17670_ (.Y(_10679_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][30] ),
    .B(net10072));
 sg13g2_o21ai_1 _17671_ (.B1(_10679_),
    .Y(_01129_),
    .A1(net9637),
    .A2(net10072));
 sg13g2_nand2_1 _17672_ (.Y(_10680_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][31] ),
    .B(net10073));
 sg13g2_o21ai_1 _17673_ (.B1(_10680_),
    .Y(_01130_),
    .A1(_10065_),
    .A2(net10073));
 sg13g2_nand2_1 _17674_ (.Y(_10681_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][3] ),
    .B(net10077));
 sg13g2_o21ai_1 _17675_ (.B1(_10681_),
    .Y(_01131_),
    .A1(net10219),
    .A2(net10077));
 sg13g2_nand2_1 _17676_ (.Y(_10682_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][4] ),
    .B(net10077));
 sg13g2_o21ai_1 _17677_ (.B1(_10682_),
    .Y(_01132_),
    .A1(net10179),
    .A2(net10077));
 sg13g2_nand2_1 _17678_ (.Y(_10683_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][5] ),
    .B(net10078));
 sg13g2_o21ai_1 _17679_ (.B1(_10683_),
    .Y(_01133_),
    .A1(net10176),
    .A2(net10078));
 sg13g2_nand2_1 _17680_ (.Y(_10684_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][6] ),
    .B(net10076));
 sg13g2_o21ai_1 _17681_ (.B1(_10684_),
    .Y(_01134_),
    .A1(net10173),
    .A2(net10076));
 sg13g2_nand2_1 _17682_ (.Y(_10685_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][7] ),
    .B(net10076));
 sg13g2_o21ai_1 _17683_ (.B1(_10685_),
    .Y(_01135_),
    .A1(net10168),
    .A2(net10076));
 sg13g2_nand2_1 _17684_ (.Y(_10686_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][8] ),
    .B(_10648_));
 sg13g2_o21ai_1 _17685_ (.B1(_10686_),
    .Y(_01136_),
    .A1(net10127),
    .A2(net10069));
 sg13g2_nand2_1 _17686_ (.Y(_10687_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][9] ),
    .B(net10076));
 sg13g2_o21ai_1 _17687_ (.B1(_10687_),
    .Y(_01137_),
    .A1(net9977),
    .A2(net10076));
 sg13g2_nand2_2 _17688_ (.Y(_10688_),
    .A(_10124_),
    .B(_10567_));
 sg13g2_buf_2 place10535 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[30] ),
    .X(net10535));
 sg13g2_buf_2 place10538 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[2] ),
    .X(net10538));
 sg13g2_buf_2 place10536 (.A(net10535),
    .X(net10536));
 sg13g2_nand2_1 _17692_ (.Y(_10692_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][0] ),
    .B(_10688_));
 sg13g2_o21ai_1 _17693_ (.B1(_10692_),
    .Y(_01138_),
    .A1(net10280),
    .A2(_10688_));
 sg13g2_nand2_1 _17694_ (.Y(_10693_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][10] ),
    .B(net9901));
 sg13g2_o21ai_1 _17695_ (.B1(_10693_),
    .Y(_01139_),
    .A1(net10132),
    .A2(net9901));
 sg13g2_nand2_1 _17696_ (.Y(_10694_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][11] ),
    .B(net9906));
 sg13g2_o21ai_1 _17697_ (.B1(_10694_),
    .Y(_01140_),
    .A1(net9983),
    .A2(net9906));
 sg13g2_nand2_1 _17698_ (.Y(_10695_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][12] ),
    .B(net9899));
 sg13g2_o21ai_1 _17699_ (.B1(_10695_),
    .Y(_01141_),
    .A1(_09885_),
    .A2(net9899));
 sg13g2_nand2_1 _17700_ (.Y(_10696_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][13] ),
    .B(net9899));
 sg13g2_o21ai_1 _17701_ (.B1(_10696_),
    .Y(_01142_),
    .A1(net9981),
    .A2(net9899));
 sg13g2_nand2_1 _17702_ (.Y(_10697_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][14] ),
    .B(net9902));
 sg13g2_o21ai_1 _17703_ (.B1(_10697_),
    .Y(_01143_),
    .A1(net9797),
    .A2(net9902));
 sg13g2_nand2_1 _17704_ (.Y(_10698_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][15] ),
    .B(net9901));
 sg13g2_o21ai_1 _17705_ (.B1(_10698_),
    .Y(_01144_),
    .A1(net9794),
    .A2(net9901));
 sg13g2_nand2_1 _17706_ (.Y(_10699_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][16] ),
    .B(net9898));
 sg13g2_o21ai_1 _17707_ (.B1(_10699_),
    .Y(_01145_),
    .A1(net9743),
    .A2(net9899));
 sg13g2_buf_2 place10534 (.A(net10533),
    .X(net10534));
 sg13g2_nand2_1 _17709_ (.Y(_10701_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][17] ),
    .B(net9899));
 sg13g2_o21ai_1 _17710_ (.B1(_10701_),
    .Y(_01146_),
    .A1(net9741),
    .A2(net9900));
 sg13g2_nand2_1 _17711_ (.Y(_10702_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][18] ),
    .B(net9904));
 sg13g2_o21ai_1 _17712_ (.B1(_10702_),
    .Y(_01147_),
    .A1(_09938_),
    .A2(net9904));
 sg13g2_buf_16 clkbuf_leaf_179_clk (.X(clknet_leaf_179_clk),
    .A(clknet_8_75_0_clk));
 sg13g2_nand2_1 _17714_ (.Y(_10704_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][19] ),
    .B(net9903));
 sg13g2_o21ai_1 _17715_ (.B1(_10704_),
    .Y(_01148_),
    .A1(_09947_),
    .A2(net9903));
 sg13g2_nand2_1 _17716_ (.Y(_10705_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][1] ),
    .B(net9899));
 sg13g2_o21ai_1 _17717_ (.B1(_10705_),
    .Y(_01149_),
    .A1(net10226),
    .A2(net9899));
 sg13g2_nand2_1 _17718_ (.Y(_10706_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][20] ),
    .B(net9904));
 sg13g2_o21ai_1 _17719_ (.B1(_10706_),
    .Y(_01150_),
    .A1(_09963_),
    .A2(net9904));
 sg13g2_nand2_1 _17720_ (.Y(_10707_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][21] ),
    .B(net9904));
 sg13g2_o21ai_1 _17721_ (.B1(_10707_),
    .Y(_01151_),
    .A1(_09972_),
    .A2(net9904));
 sg13g2_nand2_1 _17722_ (.Y(_10708_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][22] ),
    .B(net9905));
 sg13g2_o21ai_1 _17723_ (.B1(_10708_),
    .Y(_01152_),
    .A1(net9693),
    .A2(net9905));
 sg13g2_nand2_1 _17724_ (.Y(_10709_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][23] ),
    .B(net9905));
 sg13g2_o21ai_1 _17725_ (.B1(_10709_),
    .Y(_01153_),
    .A1(net9690),
    .A2(net9905));
 sg13g2_nand2_1 _17726_ (.Y(_10710_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][24] ),
    .B(net9905));
 sg13g2_o21ai_1 _17727_ (.B1(_10710_),
    .Y(_01154_),
    .A1(net9684),
    .A2(net9905));
 sg13g2_nand2_1 _17728_ (.Y(_10711_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][25] ),
    .B(net9906));
 sg13g2_o21ai_1 _17729_ (.B1(_10711_),
    .Y(_01155_),
    .A1(net9681),
    .A2(net9906));
 sg13g2_buf_2 place10533 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[31] ),
    .X(net10533));
 sg13g2_nand2_1 _17731_ (.Y(_10713_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][26] ),
    .B(net9903));
 sg13g2_o21ai_1 _17732_ (.B1(_10713_),
    .Y(_01156_),
    .A1(_10014_),
    .A2(net9903));
 sg13g2_nand2_1 _17733_ (.Y(_10714_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][27] ),
    .B(net9906));
 sg13g2_o21ai_1 _17734_ (.B1(_10714_),
    .Y(_01157_),
    .A1(net9652),
    .A2(net9906));
 sg13g2_buf_2 place10531 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[3] ),
    .X(net10531));
 sg13g2_nand2_1 _17736_ (.Y(_10716_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][28] ),
    .B(net9903));
 sg13g2_o21ai_1 _17737_ (.B1(_10716_),
    .Y(_01158_),
    .A1(_10033_),
    .A2(net9903));
 sg13g2_nand2_1 _17738_ (.Y(_10717_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][29] ),
    .B(net9906));
 sg13g2_o21ai_1 _17739_ (.B1(_10717_),
    .Y(_01159_),
    .A1(net9642),
    .A2(net9906));
 sg13g2_nand2_1 _17740_ (.Y(_10718_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][2] ),
    .B(net9901));
 sg13g2_o21ai_1 _17741_ (.B1(_10718_),
    .Y(_01160_),
    .A1(net10225),
    .A2(net9901));
 sg13g2_nand2_1 _17742_ (.Y(_10719_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][30] ),
    .B(net9902));
 sg13g2_o21ai_1 _17743_ (.B1(_10719_),
    .Y(_01161_),
    .A1(net9637),
    .A2(net9902));
 sg13g2_nand2_1 _17744_ (.Y(_10720_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][31] ),
    .B(net9903));
 sg13g2_o21ai_1 _17745_ (.B1(_10720_),
    .Y(_01162_),
    .A1(net9632),
    .A2(net9903));
 sg13g2_nand2_1 _17746_ (.Y(_10721_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][3] ),
    .B(net9898));
 sg13g2_o21ai_1 _17747_ (.B1(_10721_),
    .Y(_01163_),
    .A1(net10218),
    .A2(net9898));
 sg13g2_nand2_1 _17748_ (.Y(_10722_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][4] ),
    .B(net9898));
 sg13g2_o21ai_1 _17749_ (.B1(_10722_),
    .Y(_01164_),
    .A1(net10179),
    .A2(net9898));
 sg13g2_nand2_1 _17750_ (.Y(_10723_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][5] ),
    .B(net9901));
 sg13g2_o21ai_1 _17751_ (.B1(_10723_),
    .Y(_01165_),
    .A1(net10176),
    .A2(net9901));
 sg13g2_nand2_1 _17752_ (.Y(_10724_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][6] ),
    .B(net9900));
 sg13g2_o21ai_1 _17753_ (.B1(_10724_),
    .Y(_01166_),
    .A1(net10173),
    .A2(net9900));
 sg13g2_nand2_1 _17754_ (.Y(_10725_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][7] ),
    .B(net9900));
 sg13g2_o21ai_1 _17755_ (.B1(_10725_),
    .Y(_01167_),
    .A1(net10168),
    .A2(net9900));
 sg13g2_nand2_1 _17756_ (.Y(_10726_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][8] ),
    .B(net9904));
 sg13g2_o21ai_1 _17757_ (.B1(_10726_),
    .Y(_01168_),
    .A1(net10129),
    .A2(_10688_));
 sg13g2_nand2_1 _17758_ (.Y(_10727_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][9] ),
    .B(net9900));
 sg13g2_o21ai_1 _17759_ (.B1(_10727_),
    .Y(_01169_),
    .A1(net9977),
    .A2(net9900));
 sg13g2_nand2_2 _17760_ (.Y(_10728_),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[4] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_rd[3] ));
 sg13g2_nor2_2 _17761_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[2] ),
    .B(_10728_),
    .Y(_10729_));
 sg13g2_nand2_2 _17762_ (.Y(_10730_),
    .A(_10169_),
    .B(_10729_));
 sg13g2_buf_16 clkbuf_leaf_182_clk (.X(clknet_leaf_182_clk),
    .A(clknet_8_72_0_clk));
 sg13g2_buf_2 place10532 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[3] ),
    .X(net10532));
 sg13g2_buf_2 place10530 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[4] ),
    .X(net10530));
 sg13g2_nand2_1 _17766_ (.Y(_10734_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][0] ),
    .B(_10730_));
 sg13g2_o21ai_1 _17767_ (.B1(_10734_),
    .Y(_01170_),
    .A1(net10278),
    .A2(_10730_));
 sg13g2_nand2_1 _17768_ (.Y(_10735_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][10] ),
    .B(net10060));
 sg13g2_o21ai_1 _17769_ (.B1(_10735_),
    .Y(_01171_),
    .A1(net10130),
    .A2(net10060));
 sg13g2_nand2_1 _17770_ (.Y(_10736_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][11] ),
    .B(net10066));
 sg13g2_o21ai_1 _17771_ (.B1(_10736_),
    .Y(_01172_),
    .A1(net9984),
    .A2(net10066));
 sg13g2_nand2_1 _17772_ (.Y(_10737_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][12] ),
    .B(net10062));
 sg13g2_o21ai_1 _17773_ (.B1(_10737_),
    .Y(_01173_),
    .A1(net9799),
    .A2(net10062));
 sg13g2_nand2_1 _17774_ (.Y(_10738_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][13] ),
    .B(net10061));
 sg13g2_o21ai_1 _17775_ (.B1(_10738_),
    .Y(_01174_),
    .A1(net9978),
    .A2(net10061));
 sg13g2_nand2_1 _17776_ (.Y(_10739_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][14] ),
    .B(net10065));
 sg13g2_o21ai_1 _17777_ (.B1(_10739_),
    .Y(_01175_),
    .A1(net9795),
    .A2(net10065));
 sg13g2_nand2_1 _17778_ (.Y(_10740_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][15] ),
    .B(net10063));
 sg13g2_o21ai_1 _17779_ (.B1(_10740_),
    .Y(_01176_),
    .A1(net9791),
    .A2(net10063));
 sg13g2_nand2_1 _17780_ (.Y(_10741_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][16] ),
    .B(net10060));
 sg13g2_o21ai_1 _17781_ (.B1(_10741_),
    .Y(_01177_),
    .A1(net9746),
    .A2(net10060));
 sg13g2_buf_2 place10545 (.A(net10544),
    .X(net10545));
 sg13g2_nand2_1 _17783_ (.Y(_10743_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][17] ),
    .B(_10730_));
 sg13g2_o21ai_1 _17784_ (.B1(_10743_),
    .Y(_01178_),
    .A1(net9739),
    .A2(net10062));
 sg13g2_nand2_1 _17785_ (.Y(_10744_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][18] ),
    .B(net10064));
 sg13g2_o21ai_1 _17786_ (.B1(_10744_),
    .Y(_01179_),
    .A1(net9736),
    .A2(net10064));
 sg13g2_buf_2 place10529 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[5] ),
    .X(net10529));
 sg13g2_nand2_1 _17788_ (.Y(_10746_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][19] ),
    .B(net10067));
 sg13g2_o21ai_1 _17789_ (.B1(_10746_),
    .Y(_01180_),
    .A1(net9725),
    .A2(net10067));
 sg13g2_nand2_1 _17790_ (.Y(_10747_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][1] ),
    .B(net10061));
 sg13g2_o21ai_1 _17791_ (.B1(_10747_),
    .Y(_01181_),
    .A1(net10227),
    .A2(net10062));
 sg13g2_nand2_1 _17792_ (.Y(_10748_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][20] ),
    .B(net10068));
 sg13g2_o21ai_1 _17793_ (.B1(_10748_),
    .Y(_01182_),
    .A1(net9718),
    .A2(net10068));
 sg13g2_nand2_1 _17794_ (.Y(_10749_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][21] ),
    .B(net10064));
 sg13g2_o21ai_1 _17795_ (.B1(_10749_),
    .Y(_01183_),
    .A1(net9713),
    .A2(net10064));
 sg13g2_nand2_1 _17796_ (.Y(_10750_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][22] ),
    .B(net10068));
 sg13g2_o21ai_1 _17797_ (.B1(_10750_),
    .Y(_01184_),
    .A1(net9695),
    .A2(net10068));
 sg13g2_nand2_1 _17798_ (.Y(_10751_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][23] ),
    .B(net10068));
 sg13g2_o21ai_1 _17799_ (.B1(_10751_),
    .Y(_01185_),
    .A1(net9692),
    .A2(net10068));
 sg13g2_nand2_1 _17800_ (.Y(_10752_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][24] ),
    .B(net10068));
 sg13g2_o21ai_1 _17801_ (.B1(_10752_),
    .Y(_01186_),
    .A1(net9687),
    .A2(net10068));
 sg13g2_nand2_1 _17802_ (.Y(_10753_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][25] ),
    .B(net10065));
 sg13g2_o21ai_1 _17803_ (.B1(_10753_),
    .Y(_01187_),
    .A1(net9678),
    .A2(net10066));
 sg13g2_buf_2 place10528 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[5] ),
    .X(net10528));
 sg13g2_nand2_1 _17805_ (.Y(_10755_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][26] ),
    .B(net10067));
 sg13g2_o21ai_1 _17806_ (.B1(_10755_),
    .Y(_01188_),
    .A1(net9677),
    .A2(net10067));
 sg13g2_nand2_1 _17807_ (.Y(_10756_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][27] ),
    .B(net10067));
 sg13g2_o21ai_1 _17808_ (.B1(_10756_),
    .Y(_01189_),
    .A1(net9649),
    .A2(net10067));
 sg13g2_buf_2 place10542 (.A(net10541),
    .X(net10542));
 sg13g2_nand2_1 _17810_ (.Y(_10758_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][28] ),
    .B(net10067));
 sg13g2_o21ai_1 _17811_ (.B1(_10758_),
    .Y(_01190_),
    .A1(net9648),
    .A2(net10067));
 sg13g2_nand2_1 _17812_ (.Y(_10759_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][29] ),
    .B(net10066));
 sg13g2_o21ai_1 _17813_ (.B1(_10759_),
    .Y(_01191_),
    .A1(net9644),
    .A2(net10066));
 sg13g2_nand2_1 _17814_ (.Y(_10760_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][2] ),
    .B(net10063));
 sg13g2_o21ai_1 _17815_ (.B1(_10760_),
    .Y(_01192_),
    .A1(net10223),
    .A2(net10063));
 sg13g2_nand2_1 _17816_ (.Y(_10761_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][30] ),
    .B(net10066));
 sg13g2_o21ai_1 _17817_ (.B1(_10761_),
    .Y(_01193_),
    .A1(net9640),
    .A2(net10066));
 sg13g2_nand2_1 _17818_ (.Y(_10762_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][31] ),
    .B(net10066));
 sg13g2_o21ai_1 _17819_ (.B1(_10762_),
    .Y(_01194_),
    .A1(net9634),
    .A2(net10065));
 sg13g2_nand2_1 _17820_ (.Y(_10763_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][3] ),
    .B(net10060));
 sg13g2_o21ai_1 _17821_ (.B1(_10763_),
    .Y(_01195_),
    .A1(net10218),
    .A2(net10060));
 sg13g2_nand2_1 _17822_ (.Y(_10764_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][4] ),
    .B(net10060));
 sg13g2_o21ai_1 _17823_ (.B1(_10764_),
    .Y(_01196_),
    .A1(net10179),
    .A2(net10060));
 sg13g2_nand2_1 _17824_ (.Y(_10765_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][5] ),
    .B(net10063));
 sg13g2_o21ai_1 _17825_ (.B1(_10765_),
    .Y(_01197_),
    .A1(net10178),
    .A2(net10063));
 sg13g2_nand2_1 _17826_ (.Y(_10766_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][6] ),
    .B(net10063));
 sg13g2_o21ai_1 _17827_ (.B1(_10766_),
    .Y(_01198_),
    .A1(net10173),
    .A2(net10063));
 sg13g2_nand2_1 _17828_ (.Y(_10767_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][7] ),
    .B(net10062));
 sg13g2_o21ai_1 _17829_ (.B1(_10767_),
    .Y(_01199_),
    .A1(net10166),
    .A2(net10062));
 sg13g2_nand2_1 _17830_ (.Y(_10768_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][8] ),
    .B(net10065));
 sg13g2_o21ai_1 _17831_ (.B1(_10768_),
    .Y(_01200_),
    .A1(net10127),
    .A2(net10065));
 sg13g2_nand2_1 _17832_ (.Y(_10769_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][9] ),
    .B(net10062));
 sg13g2_o21ai_1 _17833_ (.B1(_10769_),
    .Y(_01201_),
    .A1(net9974),
    .A2(net10062));
 sg13g2_nand2_2 _17834_ (.Y(_10770_),
    .A(_10211_),
    .B(_10729_));
 sg13g2_buf_2 place10526 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[6] ),
    .X(net10526));
 sg13g2_buf_2 place10524 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[7] ),
    .X(net10524));
 sg13g2_buf_2 place10525 (.A(net10524),
    .X(net10525));
 sg13g2_nand2_1 _17838_ (.Y(_10774_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][0] ),
    .B(net9894));
 sg13g2_o21ai_1 _17839_ (.B1(_10774_),
    .Y(_01202_),
    .A1(net10277),
    .A2(net9894));
 sg13g2_nand2_1 _17840_ (.Y(_10775_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][10] ),
    .B(net9897));
 sg13g2_o21ai_1 _17841_ (.B1(_10775_),
    .Y(_01203_),
    .A1(net10130),
    .A2(net9897));
 sg13g2_nand2_1 _17842_ (.Y(_10776_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][11] ),
    .B(net9892));
 sg13g2_o21ai_1 _17843_ (.B1(_10776_),
    .Y(_01204_),
    .A1(net9984),
    .A2(net9892));
 sg13g2_nand2_1 _17844_ (.Y(_10777_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][12] ),
    .B(net9896));
 sg13g2_o21ai_1 _17845_ (.B1(_10777_),
    .Y(_01205_),
    .A1(net9799),
    .A2(net9896));
 sg13g2_nand2_1 _17846_ (.Y(_10778_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][13] ),
    .B(net9894));
 sg13g2_o21ai_1 _17847_ (.B1(_10778_),
    .Y(_01206_),
    .A1(net9978),
    .A2(net9894));
 sg13g2_nand2_1 _17848_ (.Y(_10779_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][14] ),
    .B(net9892));
 sg13g2_o21ai_1 _17849_ (.B1(_10779_),
    .Y(_01207_),
    .A1(net9795),
    .A2(net9892));
 sg13g2_nand2_1 _17850_ (.Y(_10780_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][15] ),
    .B(net9895));
 sg13g2_o21ai_1 _17851_ (.B1(_10780_),
    .Y(_01208_),
    .A1(net9791),
    .A2(net9895));
 sg13g2_nand2_1 _17852_ (.Y(_10781_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][16] ),
    .B(net9897));
 sg13g2_o21ai_1 _17853_ (.B1(_10781_),
    .Y(_01209_),
    .A1(net9746),
    .A2(net9897));
 sg13g2_buf_2 place10522 (.A(net10521),
    .X(net10522));
 sg13g2_nand2_1 _17855_ (.Y(_10783_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][17] ),
    .B(net9894));
 sg13g2_o21ai_1 _17856_ (.B1(_10783_),
    .Y(_01210_),
    .A1(_09928_),
    .A2(net9894));
 sg13g2_nand2_1 _17857_ (.Y(_10784_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][18] ),
    .B(net9889));
 sg13g2_o21ai_1 _17858_ (.B1(_10784_),
    .Y(_01211_),
    .A1(net9736),
    .A2(net9889));
 sg13g2_buf_2 place10519 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[11] ),
    .X(net10519));
 sg13g2_nand2_1 _17860_ (.Y(_10786_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][19] ),
    .B(net9893));
 sg13g2_o21ai_1 _17861_ (.B1(_10786_),
    .Y(_01212_),
    .A1(net9725),
    .A2(net9893));
 sg13g2_nand2_1 _17862_ (.Y(_10787_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][1] ),
    .B(net9896));
 sg13g2_o21ai_1 _17863_ (.B1(_10787_),
    .Y(_01213_),
    .A1(net10226),
    .A2(net9896));
 sg13g2_nand2_1 _17864_ (.Y(_10788_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][20] ),
    .B(net9890));
 sg13g2_o21ai_1 _17865_ (.B1(_10788_),
    .Y(_01214_),
    .A1(net9717),
    .A2(net9889));
 sg13g2_nand2_1 _17866_ (.Y(_10789_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][21] ),
    .B(net9889));
 sg13g2_o21ai_1 _17867_ (.B1(_10789_),
    .Y(_01215_),
    .A1(net9714),
    .A2(net9889));
 sg13g2_nand2_1 _17868_ (.Y(_10790_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][22] ),
    .B(net9890));
 sg13g2_o21ai_1 _17869_ (.B1(_10790_),
    .Y(_01216_),
    .A1(net9695),
    .A2(net9890));
 sg13g2_nand2_1 _17870_ (.Y(_10791_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][23] ),
    .B(net9890));
 sg13g2_o21ai_1 _17871_ (.B1(_10791_),
    .Y(_01217_),
    .A1(net9692),
    .A2(net9890));
 sg13g2_nand2_1 _17872_ (.Y(_10792_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][24] ),
    .B(net9890));
 sg13g2_o21ai_1 _17873_ (.B1(_10792_),
    .Y(_01218_),
    .A1(net9687),
    .A2(net9890));
 sg13g2_nand2_1 _17874_ (.Y(_10793_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][25] ),
    .B(net9891));
 sg13g2_o21ai_1 _17875_ (.B1(_10793_),
    .Y(_01219_),
    .A1(net9678),
    .A2(net9891));
 sg13g2_buf_16 clkbuf_leaf_184_clk (.X(clknet_leaf_184_clk),
    .A(clknet_8_72_0_clk));
 sg13g2_nand2_1 _17877_ (.Y(_10795_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][26] ),
    .B(net9893));
 sg13g2_o21ai_1 _17878_ (.B1(_10795_),
    .Y(_01220_),
    .A1(net9677),
    .A2(net9893));
 sg13g2_nand2_1 _17879_ (.Y(_10796_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][27] ),
    .B(net9893));
 sg13g2_o21ai_1 _17880_ (.B1(_10796_),
    .Y(_01221_),
    .A1(net9649),
    .A2(net9893));
 sg13g2_buf_2 place10518 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[12] ),
    .X(net10518));
 sg13g2_nand2_1 _17882_ (.Y(_10798_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][28] ),
    .B(net9893));
 sg13g2_o21ai_1 _17883_ (.B1(_10798_),
    .Y(_01222_),
    .A1(net9648),
    .A2(net9893));
 sg13g2_nand2_1 _17884_ (.Y(_10799_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][29] ),
    .B(net9892));
 sg13g2_o21ai_1 _17885_ (.B1(_10799_),
    .Y(_01223_),
    .A1(net9644),
    .A2(net9892));
 sg13g2_nand2_1 _17886_ (.Y(_10800_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][2] ),
    .B(net9895));
 sg13g2_o21ai_1 _17887_ (.B1(_10800_),
    .Y(_01224_),
    .A1(net10223),
    .A2(net9895));
 sg13g2_nand2_1 _17888_ (.Y(_10801_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][30] ),
    .B(net9891));
 sg13g2_o21ai_1 _17889_ (.B1(_10801_),
    .Y(_01225_),
    .A1(net9640),
    .A2(net9891));
 sg13g2_nand2_1 _17890_ (.Y(_10802_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][31] ),
    .B(net9892));
 sg13g2_o21ai_1 _17891_ (.B1(_10802_),
    .Y(_01226_),
    .A1(net9635),
    .A2(net9892));
 sg13g2_nand2_1 _17892_ (.Y(_10803_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][3] ),
    .B(net9897));
 sg13g2_o21ai_1 _17893_ (.B1(_10803_),
    .Y(_01227_),
    .A1(net10218),
    .A2(net9897));
 sg13g2_nand2_1 _17894_ (.Y(_10804_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][4] ),
    .B(net9897));
 sg13g2_o21ai_1 _17895_ (.B1(_10804_),
    .Y(_01228_),
    .A1(net10179),
    .A2(net9897));
 sg13g2_nand2_1 _17896_ (.Y(_10805_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][5] ),
    .B(net9895));
 sg13g2_o21ai_1 _17897_ (.B1(_10805_),
    .Y(_01229_),
    .A1(net10178),
    .A2(net9895));
 sg13g2_nand2_1 _17898_ (.Y(_10806_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][6] ),
    .B(net9895));
 sg13g2_o21ai_1 _17899_ (.B1(_10806_),
    .Y(_01230_),
    .A1(net10173),
    .A2(net9895));
 sg13g2_nand2_1 _17900_ (.Y(_10807_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][7] ),
    .B(net9896));
 sg13g2_o21ai_1 _17901_ (.B1(_10807_),
    .Y(_01231_),
    .A1(net10166),
    .A2(net9896));
 sg13g2_nand2_1 _17902_ (.Y(_10808_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][8] ),
    .B(net9891));
 sg13g2_o21ai_1 _17903_ (.B1(_10808_),
    .Y(_01232_),
    .A1(net10127),
    .A2(net9889));
 sg13g2_nand2_1 _17904_ (.Y(_10809_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][9] ),
    .B(net9896));
 sg13g2_o21ai_1 _17905_ (.B1(_10809_),
    .Y(_01233_),
    .A1(net9974),
    .A2(net9896));
 sg13g2_nand2_2 _17906_ (.Y(_10810_),
    .A(_09850_),
    .B(_10729_));
 sg13g2_buf_2 place10523 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[8] ),
    .X(net10523));
 sg13g2_buf_2 place10516 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[14] ),
    .X(net10516));
 sg13g2_buf_2 place10517 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[13] ),
    .X(net10517));
 sg13g2_nand2_1 _17910_ (.Y(_10814_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][0] ),
    .B(_10810_));
 sg13g2_o21ai_1 _17911_ (.B1(_10814_),
    .Y(_01234_),
    .A1(net10276),
    .A2(net10052));
 sg13g2_nand2_1 _17912_ (.Y(_10815_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][10] ),
    .B(net10051));
 sg13g2_o21ai_1 _17913_ (.B1(_10815_),
    .Y(_01235_),
    .A1(_09868_),
    .A2(net10051));
 sg13g2_nand2_1 _17914_ (.Y(_10816_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][11] ),
    .B(net10057));
 sg13g2_o21ai_1 _17915_ (.B1(_10816_),
    .Y(_01236_),
    .A1(net9984),
    .A2(net10057));
 sg13g2_nand2_1 _17916_ (.Y(_10817_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][12] ),
    .B(net10054));
 sg13g2_o21ai_1 _17917_ (.B1(_10817_),
    .Y(_01237_),
    .A1(_09885_),
    .A2(net10054));
 sg13g2_nand2_1 _17918_ (.Y(_10818_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][13] ),
    .B(net10052));
 sg13g2_o21ai_1 _17919_ (.B1(_10818_),
    .Y(_01238_),
    .A1(net9978),
    .A2(net10052));
 sg13g2_nand2_1 _17920_ (.Y(_10819_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][14] ),
    .B(net10056));
 sg13g2_o21ai_1 _17921_ (.B1(_10819_),
    .Y(_01239_),
    .A1(_09902_),
    .A2(net10056));
 sg13g2_nand2_1 _17922_ (.Y(_10820_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][15] ),
    .B(net10053));
 sg13g2_o21ai_1 _17923_ (.B1(_10820_),
    .Y(_01240_),
    .A1(net9791),
    .A2(net10053));
 sg13g2_nand2_1 _17924_ (.Y(_10821_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][16] ),
    .B(net10051));
 sg13g2_o21ai_1 _17925_ (.B1(_10821_),
    .Y(_01241_),
    .A1(_09919_),
    .A2(net10051));
 sg13g2_buf_2 place10515 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[15] ),
    .X(net10515));
 sg13g2_nand2_1 _17927_ (.Y(_10823_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][17] ),
    .B(net10052));
 sg13g2_o21ai_1 _17928_ (.B1(_10823_),
    .Y(_01242_),
    .A1(net9739),
    .A2(net10052));
 sg13g2_nand2_1 _17929_ (.Y(_10824_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][18] ),
    .B(net10055));
 sg13g2_o21ai_1 _17930_ (.B1(_10824_),
    .Y(_01243_),
    .A1(net9738),
    .A2(net10055));
 sg13g2_buf_16 clkbuf_leaf_186_clk (.X(clknet_leaf_186_clk),
    .A(clknet_8_72_0_clk));
 sg13g2_nand2_1 _17932_ (.Y(_10826_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][19] ),
    .B(net10058));
 sg13g2_o21ai_1 _17933_ (.B1(_10826_),
    .Y(_01244_),
    .A1(net9725),
    .A2(net10058));
 sg13g2_nand2_1 _17934_ (.Y(_10827_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][1] ),
    .B(net10054));
 sg13g2_o21ai_1 _17935_ (.B1(_10827_),
    .Y(_01245_),
    .A1(net10226),
    .A2(net10054));
 sg13g2_nand2_1 _17936_ (.Y(_10828_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][20] ),
    .B(net10059));
 sg13g2_o21ai_1 _17937_ (.B1(_10828_),
    .Y(_01246_),
    .A1(net9717),
    .A2(net10055));
 sg13g2_nand2_1 _17938_ (.Y(_10829_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][21] ),
    .B(net10055));
 sg13g2_o21ai_1 _17939_ (.B1(_10829_),
    .Y(_01247_),
    .A1(net9714),
    .A2(net10055));
 sg13g2_nand2_1 _17940_ (.Y(_10830_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][22] ),
    .B(net10059));
 sg13g2_o21ai_1 _17941_ (.B1(_10830_),
    .Y(_01248_),
    .A1(net9695),
    .A2(net10059));
 sg13g2_nand2_1 _17942_ (.Y(_10831_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][23] ),
    .B(net10059));
 sg13g2_o21ai_1 _17943_ (.B1(_10831_),
    .Y(_01249_),
    .A1(net9692),
    .A2(net10059));
 sg13g2_nand2_1 _17944_ (.Y(_10832_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][24] ),
    .B(net10059));
 sg13g2_o21ai_1 _17945_ (.B1(_10832_),
    .Y(_01250_),
    .A1(net9687),
    .A2(net10059));
 sg13g2_nand2_1 _17946_ (.Y(_10833_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][25] ),
    .B(net10056));
 sg13g2_o21ai_1 _17947_ (.B1(_10833_),
    .Y(_01251_),
    .A1(net9678),
    .A2(net10057));
 sg13g2_buf_2 place10514 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[19] ),
    .X(net10514));
 sg13g2_nand2_1 _17949_ (.Y(_10835_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][26] ),
    .B(net10058));
 sg13g2_o21ai_1 _17950_ (.B1(_10835_),
    .Y(_01252_),
    .A1(net9677),
    .A2(net10058));
 sg13g2_nand2_1 _17951_ (.Y(_10836_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][27] ),
    .B(net10058));
 sg13g2_o21ai_1 _17952_ (.B1(_10836_),
    .Y(_01253_),
    .A1(net9649),
    .A2(net10058));
 sg13g2_buf_16 clkbuf_leaf_188_clk (.X(clknet_leaf_188_clk),
    .A(clknet_8_74_0_clk));
 sg13g2_nand2_1 _17954_ (.Y(_10838_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][28] ),
    .B(net10058));
 sg13g2_o21ai_1 _17955_ (.B1(_10838_),
    .Y(_01254_),
    .A1(net9648),
    .A2(net10058));
 sg13g2_nand2_1 _17956_ (.Y(_10839_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][29] ),
    .B(net10057));
 sg13g2_o21ai_1 _17957_ (.B1(_10839_),
    .Y(_01255_),
    .A1(net9644),
    .A2(net10057));
 sg13g2_nand2_1 _17958_ (.Y(_10840_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][2] ),
    .B(net10053));
 sg13g2_o21ai_1 _17959_ (.B1(_10840_),
    .Y(_01256_),
    .A1(net10223),
    .A2(net10053));
 sg13g2_nand2_1 _17960_ (.Y(_10841_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][30] ),
    .B(net10057));
 sg13g2_o21ai_1 _17961_ (.B1(_10841_),
    .Y(_01257_),
    .A1(net9637),
    .A2(net10057));
 sg13g2_nand2_1 _17962_ (.Y(_10842_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][31] ),
    .B(net10057));
 sg13g2_o21ai_1 _17963_ (.B1(_10842_),
    .Y(_01258_),
    .A1(net9634),
    .A2(net10056));
 sg13g2_nand2_1 _17964_ (.Y(_10843_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][3] ),
    .B(net10051));
 sg13g2_o21ai_1 _17965_ (.B1(_10843_),
    .Y(_01259_),
    .A1(net10218),
    .A2(net10051));
 sg13g2_nand2_1 _17966_ (.Y(_10844_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][4] ),
    .B(net10051));
 sg13g2_o21ai_1 _17967_ (.B1(_10844_),
    .Y(_01260_),
    .A1(_10080_),
    .A2(net10051));
 sg13g2_nand2_1 _17968_ (.Y(_10845_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][5] ),
    .B(net10053));
 sg13g2_o21ai_1 _17969_ (.B1(_10845_),
    .Y(_01261_),
    .A1(net10178),
    .A2(net10053));
 sg13g2_nand2_1 _17970_ (.Y(_10846_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][6] ),
    .B(net10053));
 sg13g2_o21ai_1 _17971_ (.B1(_10846_),
    .Y(_01262_),
    .A1(net10173),
    .A2(net10053));
 sg13g2_nand2_1 _17972_ (.Y(_10847_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][7] ),
    .B(net10054));
 sg13g2_o21ai_1 _17973_ (.B1(_10847_),
    .Y(_01263_),
    .A1(net10166),
    .A2(net10054));
 sg13g2_nand2_1 _17974_ (.Y(_10848_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][8] ),
    .B(net10056));
 sg13g2_o21ai_1 _17975_ (.B1(_10848_),
    .Y(_01264_),
    .A1(net10127),
    .A2(net10056));
 sg13g2_nand2_1 _17976_ (.Y(_10849_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][9] ),
    .B(net10054));
 sg13g2_o21ai_1 _17977_ (.B1(_10849_),
    .Y(_01265_),
    .A1(net9974),
    .A2(net10054));
 sg13g2_nand2_2 _17978_ (.Y(_10850_),
    .A(_10124_),
    .B(_10729_));
 sg13g2_buf_2 place10513 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[1] ),
    .X(net10513));
 sg13g2_buf_16 clkbuf_leaf_194_clk (.X(clknet_leaf_194_clk),
    .A(clknet_8_22_0_clk));
 sg13g2_buf_2 place10512 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[20] ),
    .X(net10512));
 sg13g2_nand2_1 _17982_ (.Y(_10854_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][0] ),
    .B(net9881));
 sg13g2_o21ai_1 _17983_ (.B1(_10854_),
    .Y(_01266_),
    .A1(net10276),
    .A2(net9881));
 sg13g2_nand2_1 _17984_ (.Y(_10855_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][10] ),
    .B(net9885));
 sg13g2_o21ai_1 _17985_ (.B1(_10855_),
    .Y(_01267_),
    .A1(_09868_),
    .A2(net9885));
 sg13g2_nand2_1 _17986_ (.Y(_10856_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][11] ),
    .B(net9887));
 sg13g2_o21ai_1 _17987_ (.B1(_10856_),
    .Y(_01268_),
    .A1(net9984),
    .A2(net9887));
 sg13g2_nand2_1 _17988_ (.Y(_10857_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][12] ),
    .B(net9882));
 sg13g2_o21ai_1 _17989_ (.B1(_10857_),
    .Y(_01269_),
    .A1(_09885_),
    .A2(net9882));
 sg13g2_nand2_1 _17990_ (.Y(_10858_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][13] ),
    .B(net9881));
 sg13g2_o21ai_1 _17991_ (.B1(_10858_),
    .Y(_01270_),
    .A1(net9978),
    .A2(net9881));
 sg13g2_nand2_1 _17992_ (.Y(_10859_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][14] ),
    .B(net9886));
 sg13g2_o21ai_1 _17993_ (.B1(_10859_),
    .Y(_01271_),
    .A1(net9795),
    .A2(net9886));
 sg13g2_nand2_1 _17994_ (.Y(_10860_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][15] ),
    .B(net9883));
 sg13g2_o21ai_1 _17995_ (.B1(_10860_),
    .Y(_01272_),
    .A1(net9791),
    .A2(net9883));
 sg13g2_nand2_1 _17996_ (.Y(_10861_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][16] ),
    .B(net9885));
 sg13g2_o21ai_1 _17997_ (.B1(_10861_),
    .Y(_01273_),
    .A1(net9746),
    .A2(net9885));
 sg13g2_buf_16 clkbuf_leaf_195_clk (.X(clknet_leaf_195_clk),
    .A(clknet_8_19_0_clk));
 sg13g2_nand2_1 _17999_ (.Y(_10863_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][17] ),
    .B(net9881));
 sg13g2_o21ai_1 _18000_ (.B1(_10863_),
    .Y(_01274_),
    .A1(net9739),
    .A2(net9881));
 sg13g2_nand2_1 _18001_ (.Y(_10864_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][18] ),
    .B(_10850_));
 sg13g2_o21ai_1 _18002_ (.B1(_10864_),
    .Y(_01275_),
    .A1(net9736),
    .A2(_10850_));
 sg13g2_buf_2 place10511 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[23] ),
    .X(net10511));
 sg13g2_nand2_1 _18004_ (.Y(_10866_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][19] ),
    .B(net9888));
 sg13g2_o21ai_1 _18005_ (.B1(_10866_),
    .Y(_01276_),
    .A1(net9725),
    .A2(net9888));
 sg13g2_nand2_1 _18006_ (.Y(_10867_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][1] ),
    .B(net9882));
 sg13g2_o21ai_1 _18007_ (.B1(_10867_),
    .Y(_01277_),
    .A1(net10226),
    .A2(net9882));
 sg13g2_nand2_1 _18008_ (.Y(_10868_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][20] ),
    .B(net9884));
 sg13g2_o21ai_1 _18009_ (.B1(_10868_),
    .Y(_01278_),
    .A1(net9718),
    .A2(net9884));
 sg13g2_nand2_1 _18010_ (.Y(_10869_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][21] ),
    .B(_10850_));
 sg13g2_o21ai_1 _18011_ (.B1(_10869_),
    .Y(_01279_),
    .A1(net9714),
    .A2(_10850_));
 sg13g2_nand2_1 _18012_ (.Y(_10870_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][22] ),
    .B(net9884));
 sg13g2_o21ai_1 _18013_ (.B1(_10870_),
    .Y(_01280_),
    .A1(net9695),
    .A2(net9884));
 sg13g2_nand2_1 _18014_ (.Y(_10871_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][23] ),
    .B(net9884));
 sg13g2_o21ai_1 _18015_ (.B1(_10871_),
    .Y(_01281_),
    .A1(net9692),
    .A2(net9884));
 sg13g2_nand2_1 _18016_ (.Y(_10872_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][24] ),
    .B(net9884));
 sg13g2_o21ai_1 _18017_ (.B1(_10872_),
    .Y(_01282_),
    .A1(net9687),
    .A2(net9884));
 sg13g2_nand2_1 _18018_ (.Y(_10873_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][25] ),
    .B(net9886));
 sg13g2_o21ai_1 _18019_ (.B1(_10873_),
    .Y(_01283_),
    .A1(net9678),
    .A2(net9886));
 sg13g2_buf_16 clkbuf_leaf_197_clk (.X(clknet_leaf_197_clk),
    .A(clknet_8_19_0_clk));
 sg13g2_nand2_1 _18021_ (.Y(_10875_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][26] ),
    .B(net9888));
 sg13g2_o21ai_1 _18022_ (.B1(_10875_),
    .Y(_01284_),
    .A1(net9677),
    .A2(net9888));
 sg13g2_nand2_1 _18023_ (.Y(_10876_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][27] ),
    .B(net9888));
 sg13g2_o21ai_1 _18024_ (.B1(_10876_),
    .Y(_01285_),
    .A1(net9649),
    .A2(net9888));
 sg13g2_buf_16 clkbuf_leaf_196_clk (.X(clknet_leaf_196_clk),
    .A(clknet_8_19_0_clk));
 sg13g2_nand2_1 _18026_ (.Y(_10878_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][28] ),
    .B(net9888));
 sg13g2_o21ai_1 _18027_ (.B1(_10878_),
    .Y(_01286_),
    .A1(net9648),
    .A2(net9888));
 sg13g2_nand2_1 _18028_ (.Y(_10879_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][29] ),
    .B(net9887));
 sg13g2_o21ai_1 _18029_ (.B1(_10879_),
    .Y(_01287_),
    .A1(net9644),
    .A2(net9887));
 sg13g2_nand2_1 _18030_ (.Y(_10880_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][2] ),
    .B(net9883));
 sg13g2_o21ai_1 _18031_ (.B1(_10880_),
    .Y(_01288_),
    .A1(net10223),
    .A2(net9883));
 sg13g2_nand2_1 _18032_ (.Y(_10881_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][30] ),
    .B(net9887));
 sg13g2_o21ai_1 _18033_ (.B1(_10881_),
    .Y(_01289_),
    .A1(net9640),
    .A2(net9887));
 sg13g2_nand2_1 _18034_ (.Y(_10882_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][31] ),
    .B(net9887));
 sg13g2_o21ai_1 _18035_ (.B1(_10882_),
    .Y(_01290_),
    .A1(net9634),
    .A2(net9887));
 sg13g2_nand2_1 _18036_ (.Y(_10883_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][3] ),
    .B(net9885));
 sg13g2_o21ai_1 _18037_ (.B1(_10883_),
    .Y(_01291_),
    .A1(net10218),
    .A2(net9885));
 sg13g2_nand2_1 _18038_ (.Y(_10884_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][4] ),
    .B(net9885));
 sg13g2_o21ai_1 _18039_ (.B1(_10884_),
    .Y(_01292_),
    .A1(_10080_),
    .A2(net9885));
 sg13g2_nand2_1 _18040_ (.Y(_10885_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][5] ),
    .B(net9883));
 sg13g2_o21ai_1 _18041_ (.B1(_10885_),
    .Y(_01293_),
    .A1(net10178),
    .A2(net9883));
 sg13g2_nand2_1 _18042_ (.Y(_10886_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][6] ),
    .B(net9883));
 sg13g2_o21ai_1 _18043_ (.B1(_10886_),
    .Y(_01294_),
    .A1(net10173),
    .A2(net9883));
 sg13g2_nand2_1 _18044_ (.Y(_10887_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][7] ),
    .B(net9882));
 sg13g2_o21ai_1 _18045_ (.B1(_10887_),
    .Y(_01295_),
    .A1(net10166),
    .A2(net9882));
 sg13g2_nand2_1 _18046_ (.Y(_10888_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][8] ),
    .B(net9886));
 sg13g2_o21ai_1 _18047_ (.B1(_10888_),
    .Y(_01296_),
    .A1(net10127),
    .A2(net9886));
 sg13g2_nand2_1 _18048_ (.Y(_10889_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][9] ),
    .B(net9882));
 sg13g2_o21ai_1 _18049_ (.B1(_10889_),
    .Y(_01297_),
    .A1(net9974),
    .A2(net9882));
 sg13g2_nor2_2 _18050_ (.A(_00084_),
    .B(_10728_),
    .Y(_10890_));
 sg13g2_nand2_2 _18051_ (.Y(_10891_),
    .A(_10169_),
    .B(_10890_));
 sg13g2_buf_2 place10510 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[25] ),
    .X(net10510));
 sg13g2_buf_16 clkbuf_leaf_198_clk (.X(clknet_leaf_198_clk),
    .A(clknet_8_19_0_clk));
 sg13g2_buf_2 place10509 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[26] ),
    .X(net10509));
 sg13g2_nand2_1 _18055_ (.Y(_10895_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][0] ),
    .B(_10891_));
 sg13g2_o21ai_1 _18056_ (.B1(_10895_),
    .Y(_01298_),
    .A1(_09836_),
    .A2(net10049));
 sg13g2_nand2_1 _18057_ (.Y(_10896_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][10] ),
    .B(net10047));
 sg13g2_o21ai_1 _18058_ (.B1(_10896_),
    .Y(_01299_),
    .A1(net10130),
    .A2(net10047));
 sg13g2_nand2_1 _18059_ (.Y(_10897_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][11] ),
    .B(net10043));
 sg13g2_o21ai_1 _18060_ (.B1(_10897_),
    .Y(_01300_),
    .A1(net9984),
    .A2(net10043));
 sg13g2_nand2_1 _18061_ (.Y(_10898_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][12] ),
    .B(net10050));
 sg13g2_o21ai_1 _18062_ (.B1(_10898_),
    .Y(_01301_),
    .A1(net9799),
    .A2(net10050));
 sg13g2_nand2_1 _18063_ (.Y(_10899_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][13] ),
    .B(net10049));
 sg13g2_o21ai_1 _18064_ (.B1(_10899_),
    .Y(_01302_),
    .A1(net9978),
    .A2(net10049));
 sg13g2_nand2_1 _18065_ (.Y(_10900_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][14] ),
    .B(net10042));
 sg13g2_o21ai_1 _18066_ (.B1(_10900_),
    .Y(_01303_),
    .A1(net9798),
    .A2(net10042));
 sg13g2_nand2_1 _18067_ (.Y(_10901_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][15] ),
    .B(net10047));
 sg13g2_o21ai_1 _18068_ (.B1(_10901_),
    .Y(_01304_),
    .A1(_09911_),
    .A2(net10047));
 sg13g2_nand2_1 _18069_ (.Y(_10902_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][16] ),
    .B(net10046));
 sg13g2_o21ai_1 _18070_ (.B1(_10902_),
    .Y(_01305_),
    .A1(_09919_),
    .A2(net10046));
 sg13g2_buf_16 clkbuf_leaf_200_clk (.X(clknet_leaf_200_clk),
    .A(clknet_8_21_0_clk));
 sg13g2_nand2_1 _18072_ (.Y(_10904_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][17] ),
    .B(net10049));
 sg13g2_o21ai_1 _18073_ (.B1(_10904_),
    .Y(_01306_),
    .A1(net9739),
    .A2(net10049));
 sg13g2_nand2_1 _18074_ (.Y(_10905_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][18] ),
    .B(net10045));
 sg13g2_o21ai_1 _18075_ (.B1(_10905_),
    .Y(_01307_),
    .A1(net9737),
    .A2(net10046));
 sg13g2_buf_2 place10508 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[27] ),
    .X(net10508));
 sg13g2_nand2_1 _18077_ (.Y(_10907_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][19] ),
    .B(net10044));
 sg13g2_o21ai_1 _18078_ (.B1(_10907_),
    .Y(_01308_),
    .A1(net9725),
    .A2(net10044));
 sg13g2_nand2_1 _18079_ (.Y(_10908_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][1] ),
    .B(net10049));
 sg13g2_o21ai_1 _18080_ (.B1(_10908_),
    .Y(_01309_),
    .A1(_09954_),
    .A2(net10049));
 sg13g2_nand2_1 _18081_ (.Y(_10909_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][20] ),
    .B(net10048));
 sg13g2_o21ai_1 _18082_ (.B1(_10909_),
    .Y(_01310_),
    .A1(net9717),
    .A2(net10048));
 sg13g2_nand2_1 _18083_ (.Y(_10910_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][21] ),
    .B(net10045));
 sg13g2_o21ai_1 _18084_ (.B1(_10910_),
    .Y(_01311_),
    .A1(net9713),
    .A2(net10045));
 sg13g2_nand2_1 _18085_ (.Y(_10911_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][22] ),
    .B(net10048));
 sg13g2_o21ai_1 _18086_ (.B1(_10911_),
    .Y(_01312_),
    .A1(net9696),
    .A2(net10048));
 sg13g2_nand2_1 _18087_ (.Y(_10912_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][23] ),
    .B(net10048));
 sg13g2_o21ai_1 _18088_ (.B1(_10912_),
    .Y(_01313_),
    .A1(net9691),
    .A2(net10048));
 sg13g2_nand2_1 _18089_ (.Y(_10913_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][24] ),
    .B(net10048));
 sg13g2_o21ai_1 _18090_ (.B1(_10913_),
    .Y(_01314_),
    .A1(net9686),
    .A2(net10048));
 sg13g2_nand2_1 _18091_ (.Y(_10914_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][25] ),
    .B(net10042));
 sg13g2_o21ai_1 _18092_ (.B1(_10914_),
    .Y(_01315_),
    .A1(net9678),
    .A2(net10043));
 sg13g2_buf_2 place10507 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[28] ),
    .X(net10507));
 sg13g2_nand2_1 _18094_ (.Y(_10916_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][26] ),
    .B(net10044));
 sg13g2_o21ai_1 _18095_ (.B1(_10916_),
    .Y(_01316_),
    .A1(net9677),
    .A2(net10044));
 sg13g2_nand2_1 _18096_ (.Y(_10917_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][27] ),
    .B(net10044));
 sg13g2_o21ai_1 _18097_ (.B1(_10917_),
    .Y(_01317_),
    .A1(net9649),
    .A2(net10044));
 sg13g2_buf_2 place10506 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[29] ),
    .X(net10506));
 sg13g2_nand2_1 _18099_ (.Y(_10919_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][28] ),
    .B(net10044));
 sg13g2_o21ai_1 _18100_ (.B1(_10919_),
    .Y(_01318_),
    .A1(net9648),
    .A2(net10044));
 sg13g2_nand2_1 _18101_ (.Y(_10920_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][29] ),
    .B(net10043));
 sg13g2_o21ai_1 _18102_ (.B1(_10920_),
    .Y(_01319_),
    .A1(net9644),
    .A2(net10043));
 sg13g2_nand2_1 _18103_ (.Y(_10921_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][2] ),
    .B(net10047));
 sg13g2_o21ai_1 _18104_ (.B1(_10921_),
    .Y(_01320_),
    .A1(net10223),
    .A2(net10047));
 sg13g2_nand2_1 _18105_ (.Y(_10922_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][30] ),
    .B(net10043));
 sg13g2_o21ai_1 _18106_ (.B1(_10922_),
    .Y(_01321_),
    .A1(net9640),
    .A2(net10043));
 sg13g2_nand2_1 _18107_ (.Y(_10923_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][31] ),
    .B(net10043));
 sg13g2_o21ai_1 _18108_ (.B1(_10923_),
    .Y(_01322_),
    .A1(net9634),
    .A2(net10042));
 sg13g2_nand2_1 _18109_ (.Y(_10924_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][3] ),
    .B(net10046));
 sg13g2_o21ai_1 _18110_ (.B1(_10924_),
    .Y(_01323_),
    .A1(_10072_),
    .A2(net10046));
 sg13g2_nand2_1 _18111_ (.Y(_10925_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][4] ),
    .B(net10045));
 sg13g2_o21ai_1 _18112_ (.B1(_10925_),
    .Y(_01324_),
    .A1(_10080_),
    .A2(net10045));
 sg13g2_nand2_1 _18113_ (.Y(_10926_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][5] ),
    .B(net10047));
 sg13g2_o21ai_1 _18114_ (.B1(_10926_),
    .Y(_01325_),
    .A1(net10174),
    .A2(net10047));
 sg13g2_nand2_1 _18115_ (.Y(_10927_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][6] ),
    .B(net10050));
 sg13g2_o21ai_1 _18116_ (.B1(_10927_),
    .Y(_01326_),
    .A1(_10095_),
    .A2(net10050));
 sg13g2_nand2_1 _18117_ (.Y(_10928_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][7] ),
    .B(net10050));
 sg13g2_o21ai_1 _18118_ (.B1(_10928_),
    .Y(_01327_),
    .A1(_10103_),
    .A2(net10050));
 sg13g2_nand2_1 _18119_ (.Y(_10929_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][8] ),
    .B(net10042));
 sg13g2_o21ai_1 _18120_ (.B1(_10929_),
    .Y(_01328_),
    .A1(_10111_),
    .A2(net10042));
 sg13g2_nand2_1 _18121_ (.Y(_10930_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][9] ),
    .B(net10050));
 sg13g2_o21ai_1 _18122_ (.B1(_10930_),
    .Y(_01329_),
    .A1(net9974),
    .A2(net10050));
 sg13g2_buf_2 place10505 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[2] ),
    .X(net10505));
 sg13g2_nand2_2 _18124_ (.Y(_10932_),
    .A(_10211_),
    .B(_10890_));
 sg13g2_buf_2 place10504 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[4] ),
    .X(net10504));
 sg13g2_buf_2 place10503 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[5] ),
    .X(net10503));
 sg13g2_buf_2 place10502 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[6] ),
    .X(net10502));
 sg13g2_nand2_1 _18128_ (.Y(_10936_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][0] ),
    .B(_10932_));
 sg13g2_o21ai_1 _18129_ (.B1(_10936_),
    .Y(_01330_),
    .A1(net10279),
    .A2(net9872));
 sg13g2_buf_2 place10501 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[7] ),
    .X(net10501));
 sg13g2_nand2_1 _18131_ (.Y(_10938_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][10] ),
    .B(net9875));
 sg13g2_o21ai_1 _18132_ (.B1(_10938_),
    .Y(_01331_),
    .A1(net10130),
    .A2(net9875));
 sg13g2_buf_2 place10500 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[8] ),
    .X(net10500));
 sg13g2_nand2_1 _18134_ (.Y(_10940_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][11] ),
    .B(net9879));
 sg13g2_o21ai_1 _18135_ (.B1(_10940_),
    .Y(_01332_),
    .A1(net9984),
    .A2(net9879));
 sg13g2_buf_2 place10499 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[9] ),
    .X(net10499));
 sg13g2_nand2_1 _18137_ (.Y(_10942_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][12] ),
    .B(net9873));
 sg13g2_o21ai_1 _18138_ (.B1(_10942_),
    .Y(_01333_),
    .A1(net9799),
    .A2(net9873));
 sg13g2_buf_2 place10498 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[10] ),
    .X(net10498));
 sg13g2_nand2_1 _18140_ (.Y(_10944_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][13] ),
    .B(net9872));
 sg13g2_o21ai_1 _18141_ (.B1(_10944_),
    .Y(_01334_),
    .A1(_09894_),
    .A2(net9872));
 sg13g2_buf_2 place10497 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[11] ),
    .X(net10497));
 sg13g2_nand2_1 _18143_ (.Y(_10946_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][14] ),
    .B(net9878));
 sg13g2_o21ai_1 _18144_ (.B1(_10946_),
    .Y(_01335_),
    .A1(net9798),
    .A2(_10932_));
 sg13g2_buf_2 place10496 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[15] ),
    .X(net10496));
 sg13g2_nand2_1 _18146_ (.Y(_10948_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][15] ),
    .B(net9875));
 sg13g2_o21ai_1 _18147_ (.B1(_10948_),
    .Y(_01336_),
    .A1(_09911_),
    .A2(net9875));
 sg13g2_buf_16 clkbuf_leaf_201_clk (.X(clknet_leaf_201_clk),
    .A(clknet_8_17_0_clk));
 sg13g2_nand2_1 _18149_ (.Y(_10950_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][16] ),
    .B(net9874));
 sg13g2_o21ai_1 _18150_ (.B1(_10950_),
    .Y(_01337_),
    .A1(_09919_),
    .A2(net9874));
 sg13g2_buf_2 place10495 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[21] ),
    .X(net10495));
 sg13g2_buf_16 clkbuf_leaf_203_clk (.X(clknet_leaf_203_clk),
    .A(clknet_8_23_0_clk));
 sg13g2_nand2_1 _18153_ (.Y(_10953_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][17] ),
    .B(net9872));
 sg13g2_o21ai_1 _18154_ (.B1(_10953_),
    .Y(_01338_),
    .A1(_09928_),
    .A2(net9872));
 sg13g2_buf_2 place10494 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[22] ),
    .X(net10494));
 sg13g2_nand2_1 _18156_ (.Y(_10955_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][18] ),
    .B(net9874));
 sg13g2_o21ai_1 _18157_ (.B1(_10955_),
    .Y(_01339_),
    .A1(net9736),
    .A2(net9874));
 sg13g2_buf_2 place10493 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[25] ),
    .X(net10493));
 sg13g2_buf_16 clkbuf_leaf_204_clk (.X(clknet_leaf_204_clk),
    .A(clknet_8_72_0_clk));
 sg13g2_nand2_1 _18160_ (.Y(_10958_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][19] ),
    .B(net9880));
 sg13g2_o21ai_1 _18161_ (.B1(_10958_),
    .Y(_01340_),
    .A1(net9725),
    .A2(net9880));
 sg13g2_buf_2 place10521 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[9] ),
    .X(net10521));
 sg13g2_nand2_1 _18163_ (.Y(_10960_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][1] ),
    .B(net9872));
 sg13g2_o21ai_1 _18164_ (.B1(_10960_),
    .Y(_01341_),
    .A1(_09954_),
    .A2(net9872));
 sg13g2_buf_16 clkbuf_leaf_205_clk (.X(clknet_leaf_205_clk),
    .A(clknet_8_23_0_clk));
 sg13g2_nand2_1 _18166_ (.Y(_10962_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][20] ),
    .B(net9877));
 sg13g2_o21ai_1 _18167_ (.B1(_10962_),
    .Y(_01342_),
    .A1(net9717),
    .A2(net9877));
 sg13g2_buf_2 place10491 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[2] ),
    .X(net10491));
 sg13g2_nand2_1 _18169_ (.Y(_10964_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][21] ),
    .B(net9876));
 sg13g2_o21ai_1 _18170_ (.B1(_10964_),
    .Y(_01343_),
    .A1(net9713),
    .A2(net9876));
 sg13g2_buf_2 place10492 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[26] ),
    .X(net10492));
 sg13g2_nand2_1 _18172_ (.Y(_10966_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][22] ),
    .B(net9877));
 sg13g2_o21ai_1 _18173_ (.B1(_10966_),
    .Y(_01344_),
    .A1(net9696),
    .A2(net9877));
 sg13g2_buf_2 place10490 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[3] ),
    .X(net10490));
 sg13g2_nand2_1 _18175_ (.Y(_10968_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][23] ),
    .B(net9877));
 sg13g2_o21ai_1 _18176_ (.B1(_10968_),
    .Y(_01345_),
    .A1(net9691),
    .A2(net9877));
 sg13g2_buf_2 place10541 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[29] ),
    .X(net10541));
 sg13g2_nand2_1 _18178_ (.Y(_10970_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][24] ),
    .B(net9877));
 sg13g2_o21ai_1 _18179_ (.B1(_10970_),
    .Y(_01346_),
    .A1(net9686),
    .A2(net9877));
 sg13g2_buf_2 place10520 (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[0] ),
    .X(net10520));
 sg13g2_nand2_1 _18181_ (.Y(_10972_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][25] ),
    .B(net9879));
 sg13g2_o21ai_1 _18182_ (.B1(_10972_),
    .Y(_01347_),
    .A1(net9679),
    .A2(net9879));
 sg13g2_buf_2 place10537 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[30] ),
    .X(net10537));
 sg13g2_buf_2 place10485 (.A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[31] ),
    .X(net10485));
 sg13g2_nand2_1 _18185_ (.Y(_10975_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][26] ),
    .B(net9880));
 sg13g2_o21ai_1 _18186_ (.B1(_10975_),
    .Y(_01348_),
    .A1(net9677),
    .A2(net9880));
 sg13g2_buf_16 clkbuf_leaf_207_clk (.X(clknet_leaf_207_clk),
    .A(clknet_8_20_0_clk));
 sg13g2_nand2_1 _18188_ (.Y(_10977_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][27] ),
    .B(net9880));
 sg13g2_o21ai_1 _18189_ (.B1(_10977_),
    .Y(_01349_),
    .A1(net9649),
    .A2(net9880));
 sg13g2_buf_2 place10484 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[11] ),
    .X(net10484));
 sg13g2_buf_2 place10483 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[12] ),
    .X(net10483));
 sg13g2_nand2_1 _18192_ (.Y(_10980_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][28] ),
    .B(net9880));
 sg13g2_o21ai_1 _18193_ (.B1(_10980_),
    .Y(_01350_),
    .A1(net9648),
    .A2(net9880));
 sg13g2_buf_2 place10482 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[13] ),
    .X(net10482));
 sg13g2_nand2_1 _18195_ (.Y(_10982_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][29] ),
    .B(net9879));
 sg13g2_o21ai_1 _18196_ (.B1(_10982_),
    .Y(_01351_),
    .A1(net9644),
    .A2(net9879));
 sg13g2_buf_16 clkbuf_leaf_208_clk (.X(clknet_leaf_208_clk),
    .A(clknet_8_20_0_clk));
 sg13g2_nand2_1 _18198_ (.Y(_10984_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][2] ),
    .B(net9875));
 sg13g2_o21ai_1 _18199_ (.B1(_10984_),
    .Y(_01352_),
    .A1(net10223),
    .A2(net9875));
 sg13g2_buf_2 place10487 (.A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[22] ),
    .X(net10487));
 sg13g2_nand2_1 _18201_ (.Y(_10986_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][30] ),
    .B(net9878));
 sg13g2_o21ai_1 _18202_ (.B1(_10986_),
    .Y(_01353_),
    .A1(net9640),
    .A2(net9879));
 sg13g2_buf_2 place10486 (.A(net10485),
    .X(net10486));
 sg13g2_nand2_1 _18204_ (.Y(_10988_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][31] ),
    .B(net9878));
 sg13g2_o21ai_1 _18205_ (.B1(_10988_),
    .Y(_01354_),
    .A1(net9634),
    .A2(net9878));
 sg13g2_buf_16 clkbuf_leaf_212_clk (.X(clknet_leaf_212_clk),
    .A(clknet_8_17_0_clk));
 sg13g2_nand2_1 _18207_ (.Y(_10990_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][3] ),
    .B(net9874));
 sg13g2_o21ai_1 _18208_ (.B1(_10990_),
    .Y(_01355_),
    .A1(_10072_),
    .A2(net9874));
 sg13g2_buf_2 place10479 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2] ),
    .X(net10479));
 sg13g2_nand2_1 _18210_ (.Y(_10992_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][4] ),
    .B(net9876));
 sg13g2_o21ai_1 _18211_ (.B1(_10992_),
    .Y(_01356_),
    .A1(_10080_),
    .A2(net9876));
 sg13g2_buf_2 place10478 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[3] ),
    .X(net10478));
 sg13g2_nand2_1 _18213_ (.Y(_10994_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][5] ),
    .B(net9875));
 sg13g2_o21ai_1 _18214_ (.B1(_10994_),
    .Y(_01357_),
    .A1(net10174),
    .A2(net9875));
 sg13g2_buf_16 clkbuf_leaf_214_clk (.X(clknet_leaf_214_clk),
    .A(clknet_8_16_0_clk));
 sg13g2_nand2_1 _18216_ (.Y(_10996_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][6] ),
    .B(net9873));
 sg13g2_o21ai_1 _18217_ (.B1(_10996_),
    .Y(_01358_),
    .A1(_10095_),
    .A2(net9873));
 sg13g2_buf_2 place10477 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[4] ),
    .X(net10477));
 sg13g2_nand2_1 _18219_ (.Y(_10998_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][7] ),
    .B(net9873));
 sg13g2_o21ai_1 _18220_ (.B1(_10998_),
    .Y(_01359_),
    .A1(_10103_),
    .A2(net9873));
 sg13g2_buf_2 place10489 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[4] ),
    .X(net10489));
 sg13g2_nand2_1 _18222_ (.Y(_11000_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][8] ),
    .B(_10932_));
 sg13g2_o21ai_1 _18223_ (.B1(_11000_),
    .Y(_01360_),
    .A1(_10111_),
    .A2(_10932_));
 sg13g2_buf_2 place10481 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[18] ),
    .X(net10481));
 sg13g2_nand2_1 _18225_ (.Y(_11002_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][9] ),
    .B(net9873));
 sg13g2_o21ai_1 _18226_ (.B1(_11002_),
    .Y(_01361_),
    .A1(_10119_),
    .A2(net9873));
 sg13g2_nand2_1 _18227_ (.Y(_11003_),
    .A(_09850_),
    .B(_10168_));
 sg13g2_buf_2 place10480 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[22] ),
    .X(net10480));
 sg13g2_buf_2 place10476 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[5] ),
    .X(net10476));
 sg13g2_buf_2 place10540 (.A(net10539),
    .X(net10540));
 sg13g2_nand2_1 _18231_ (.Y(_11007_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][0] ),
    .B(net10032));
 sg13g2_o21ai_1 _18232_ (.B1(_11007_),
    .Y(_01362_),
    .A1(net10278),
    .A2(net10032));
 sg13g2_nand2_1 _18233_ (.Y(_11008_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][10] ),
    .B(net10037));
 sg13g2_o21ai_1 _18234_ (.B1(_11008_),
    .Y(_01363_),
    .A1(net10132),
    .A2(net10037));
 sg13g2_nand2_1 _18235_ (.Y(_11009_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][11] ),
    .B(net10041));
 sg13g2_o21ai_1 _18236_ (.B1(_11009_),
    .Y(_01364_),
    .A1(net9983),
    .A2(net10040));
 sg13g2_nand2_1 _18237_ (.Y(_11010_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][12] ),
    .B(net10034));
 sg13g2_o21ai_1 _18238_ (.B1(_11010_),
    .Y(_01365_),
    .A1(net9801),
    .A2(net10034));
 sg13g2_nand2_1 _18239_ (.Y(_11011_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][13] ),
    .B(net10032));
 sg13g2_o21ai_1 _18240_ (.B1(_11011_),
    .Y(_01366_),
    .A1(net9980),
    .A2(net10032));
 sg13g2_nand2_1 _18241_ (.Y(_11012_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][14] ),
    .B(net10038));
 sg13g2_o21ai_1 _18242_ (.B1(_11012_),
    .Y(_01367_),
    .A1(net9796),
    .A2(net10038));
 sg13g2_nand2_1 _18243_ (.Y(_11013_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][15] ),
    .B(net10033));
 sg13g2_o21ai_1 _18244_ (.B1(_11013_),
    .Y(_01368_),
    .A1(net9792),
    .A2(net10033));
 sg13g2_nand2_1 _18245_ (.Y(_11014_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][16] ),
    .B(net10033));
 sg13g2_o21ai_1 _18246_ (.B1(_11014_),
    .Y(_01369_),
    .A1(net9744),
    .A2(net10032));
 sg13g2_buf_2 place10471 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_inc ),
    .X(net10471));
 sg13g2_nand2_1 _18248_ (.Y(_11016_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][17] ),
    .B(net10033));
 sg13g2_o21ai_1 _18249_ (.B1(_11016_),
    .Y(_01370_),
    .A1(net9740),
    .A2(net10033));
 sg13g2_nand2_1 _18250_ (.Y(_11017_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][18] ),
    .B(net10036));
 sg13g2_o21ai_1 _18251_ (.B1(_11017_),
    .Y(_01371_),
    .A1(net9737),
    .A2(net10036));
 sg13g2_buf_16 clkbuf_leaf_221_clk (.X(clknet_leaf_221_clk),
    .A(clknet_8_64_0_clk));
 sg13g2_nand2_1 _18253_ (.Y(_11019_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][19] ),
    .B(net10039));
 sg13g2_o21ai_1 _18254_ (.B1(_11019_),
    .Y(_01372_),
    .A1(_09947_),
    .A2(net10039));
 sg13g2_nand2_1 _18255_ (.Y(_11020_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][1] ),
    .B(net10034));
 sg13g2_o21ai_1 _18256_ (.B1(_11020_),
    .Y(_01373_),
    .A1(net10229),
    .A2(net10034));
 sg13g2_nand2_1 _18257_ (.Y(_11021_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][20] ),
    .B(net10036));
 sg13g2_o21ai_1 _18258_ (.B1(_11021_),
    .Y(_01374_),
    .A1(net9720),
    .A2(net10036));
 sg13g2_nand2_1 _18259_ (.Y(_11022_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][21] ),
    .B(net10036));
 sg13g2_o21ai_1 _18260_ (.B1(_11022_),
    .Y(_01375_),
    .A1(net9715),
    .A2(net10036));
 sg13g2_nand2_1 _18261_ (.Y(_11023_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][22] ),
    .B(net10040));
 sg13g2_o21ai_1 _18262_ (.B1(_11023_),
    .Y(_01376_),
    .A1(_09980_),
    .A2(net10040));
 sg13g2_nand2_1 _18263_ (.Y(_11024_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][23] ),
    .B(net10040));
 sg13g2_o21ai_1 _18264_ (.B1(_11024_),
    .Y(_01377_),
    .A1(_09988_),
    .A2(net10040));
 sg13g2_nand2_1 _18265_ (.Y(_11025_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][24] ),
    .B(net10040));
 sg13g2_o21ai_1 _18266_ (.B1(_11025_),
    .Y(_01378_),
    .A1(_09997_),
    .A2(net10040));
 sg13g2_nand2_1 _18267_ (.Y(_11026_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][25] ),
    .B(net10041));
 sg13g2_o21ai_1 _18268_ (.B1(_11026_),
    .Y(_01379_),
    .A1(net9681),
    .A2(net10041));
 sg13g2_buf_16 clkbuf_leaf_220_clk (.X(clknet_leaf_220_clk),
    .A(clknet_8_64_0_clk));
 sg13g2_nand2_1 _18270_ (.Y(_11028_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][26] ),
    .B(net10039));
 sg13g2_o21ai_1 _18271_ (.B1(_11028_),
    .Y(_01380_),
    .A1(net9674),
    .A2(net10039));
 sg13g2_nand2_1 _18272_ (.Y(_11029_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][27] ),
    .B(net10041));
 sg13g2_o21ai_1 _18273_ (.B1(_11029_),
    .Y(_01381_),
    .A1(net9652),
    .A2(net10041));
 sg13g2_buf_16 clkbuf_leaf_218_clk (.X(clknet_leaf_218_clk),
    .A(clknet_8_21_0_clk));
 sg13g2_nand2_1 _18275_ (.Y(_11031_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][28] ),
    .B(net10039));
 sg13g2_o21ai_1 _18276_ (.B1(_11031_),
    .Y(_01382_),
    .A1(_10033_),
    .A2(net10039));
 sg13g2_nand2_1 _18277_ (.Y(_11032_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][29] ),
    .B(net10041));
 sg13g2_o21ai_1 _18278_ (.B1(_11032_),
    .Y(_01383_),
    .A1(net9642),
    .A2(net10041));
 sg13g2_nand2_1 _18279_ (.Y(_11033_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][2] ),
    .B(net10033));
 sg13g2_o21ai_1 _18280_ (.B1(_11033_),
    .Y(_01384_),
    .A1(net10225),
    .A2(net10033));
 sg13g2_nand2_1 _18281_ (.Y(_11034_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][30] ),
    .B(net10038));
 sg13g2_o21ai_1 _18282_ (.B1(_11034_),
    .Y(_01385_),
    .A1(_10056_),
    .A2(net10038));
 sg13g2_nand2_1 _18283_ (.Y(_11035_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][31] ),
    .B(net10039));
 sg13g2_o21ai_1 _18284_ (.B1(_11035_),
    .Y(_01386_),
    .A1(net9632),
    .A2(net10039));
 sg13g2_nand2_1 _18285_ (.Y(_11036_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][3] ),
    .B(net10037));
 sg13g2_o21ai_1 _18286_ (.B1(_11036_),
    .Y(_01387_),
    .A1(net10221),
    .A2(net10037));
 sg13g2_nand2_1 _18287_ (.Y(_11037_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][4] ),
    .B(net10037));
 sg13g2_o21ai_1 _18288_ (.B1(_11037_),
    .Y(_01388_),
    .A1(net10180),
    .A2(net10037));
 sg13g2_nand2_1 _18289_ (.Y(_11038_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][5] ),
    .B(net10037));
 sg13g2_o21ai_1 _18290_ (.B1(_11038_),
    .Y(_01389_),
    .A1(net10177),
    .A2(net10037));
 sg13g2_nand2_1 _18291_ (.Y(_11039_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][6] ),
    .B(net10035));
 sg13g2_o21ai_1 _18292_ (.B1(_11039_),
    .Y(_01390_),
    .A1(net10172),
    .A2(net10035));
 sg13g2_nand2_1 _18293_ (.Y(_11040_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][7] ),
    .B(net10035));
 sg13g2_o21ai_1 _18294_ (.B1(_11040_),
    .Y(_01391_),
    .A1(net10169),
    .A2(net10035));
 sg13g2_nand2_1 _18295_ (.Y(_11041_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][8] ),
    .B(net10038));
 sg13g2_o21ai_1 _18296_ (.B1(_11041_),
    .Y(_01392_),
    .A1(net10126),
    .A2(net10038));
 sg13g2_nand2_1 _18297_ (.Y(_11042_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][9] ),
    .B(net10035));
 sg13g2_o21ai_1 _18298_ (.B1(_11042_),
    .Y(_01393_),
    .A1(net9977),
    .A2(net10035));
 sg13g2_nand2_2 _18299_ (.Y(_11043_),
    .A(_09850_),
    .B(_10890_));
 sg13g2_buf_16 clkbuf_leaf_216_clk (.X(clknet_leaf_216_clk),
    .A(clknet_8_20_0_clk));
 sg13g2_buf_2 place10470 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[1] ),
    .X(net10470));
 sg13g2_buf_2 place10562 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[21] ),
    .X(net10562));
 sg13g2_nand2_1 _18303_ (.Y(_11047_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][0] ),
    .B(_11043_));
 sg13g2_o21ai_1 _18304_ (.B1(_11047_),
    .Y(_01394_),
    .A1(net10276),
    .A2(net10023));
 sg13g2_nand2_1 _18305_ (.Y(_11048_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][10] ),
    .B(net10026));
 sg13g2_o21ai_1 _18306_ (.B1(_11048_),
    .Y(_01395_),
    .A1(net10130),
    .A2(net10026));
 sg13g2_nand2_1 _18307_ (.Y(_11049_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][11] ),
    .B(net10030));
 sg13g2_o21ai_1 _18308_ (.B1(_11049_),
    .Y(_01396_),
    .A1(net9984),
    .A2(net10030));
 sg13g2_nand2_1 _18309_ (.Y(_11050_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][12] ),
    .B(net10024));
 sg13g2_o21ai_1 _18310_ (.B1(_11050_),
    .Y(_01397_),
    .A1(net9799),
    .A2(net10024));
 sg13g2_nand2_1 _18311_ (.Y(_11051_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][13] ),
    .B(net10023));
 sg13g2_o21ai_1 _18312_ (.B1(_11051_),
    .Y(_01398_),
    .A1(_09894_),
    .A2(net10023));
 sg13g2_nand2_1 _18313_ (.Y(_11052_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][14] ),
    .B(net10029));
 sg13g2_o21ai_1 _18314_ (.B1(_11052_),
    .Y(_01399_),
    .A1(net9798),
    .A2(net10029));
 sg13g2_nand2_1 _18315_ (.Y(_11053_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][15] ),
    .B(net10026));
 sg13g2_o21ai_1 _18316_ (.B1(_11053_),
    .Y(_01400_),
    .A1(_09911_),
    .A2(net10026));
 sg13g2_nand2_1 _18317_ (.Y(_11054_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][16] ),
    .B(net10025));
 sg13g2_o21ai_1 _18318_ (.B1(_11054_),
    .Y(_01401_),
    .A1(_09919_),
    .A2(net10025));
 sg13g2_buf_2 place10576 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[18] ),
    .X(net10576));
 sg13g2_nand2_1 _18320_ (.Y(_11056_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][17] ),
    .B(net10023));
 sg13g2_o21ai_1 _18321_ (.B1(_11056_),
    .Y(_01402_),
    .A1(net9741),
    .A2(net10023));
 sg13g2_nand2_1 _18322_ (.Y(_11057_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][18] ),
    .B(net10027));
 sg13g2_o21ai_1 _18323_ (.B1(_11057_),
    .Y(_01403_),
    .A1(net9737),
    .A2(net10025));
 sg13g2_buf_2 place10720 (.A(net10719),
    .X(net10720));
 sg13g2_nand2_1 _18325_ (.Y(_11059_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][19] ),
    .B(net10031));
 sg13g2_o21ai_1 _18326_ (.B1(_11059_),
    .Y(_01404_),
    .A1(net9725),
    .A2(net10031));
 sg13g2_nand2_1 _18327_ (.Y(_11060_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][1] ),
    .B(net10023));
 sg13g2_o21ai_1 _18328_ (.B1(_11060_),
    .Y(_01405_),
    .A1(_09954_),
    .A2(net10023));
 sg13g2_nand2_1 _18329_ (.Y(_11061_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][20] ),
    .B(net10028));
 sg13g2_o21ai_1 _18330_ (.B1(_11061_),
    .Y(_01406_),
    .A1(net9717),
    .A2(net10028));
 sg13g2_nand2_1 _18331_ (.Y(_11062_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][21] ),
    .B(net10027));
 sg13g2_o21ai_1 _18332_ (.B1(_11062_),
    .Y(_01407_),
    .A1(net9712),
    .A2(net10027));
 sg13g2_nand2_1 _18333_ (.Y(_11063_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][22] ),
    .B(net10028));
 sg13g2_o21ai_1 _18334_ (.B1(_11063_),
    .Y(_01408_),
    .A1(net9694),
    .A2(net10028));
 sg13g2_nand2_1 _18335_ (.Y(_11064_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][23] ),
    .B(net10028));
 sg13g2_o21ai_1 _18336_ (.B1(_11064_),
    .Y(_01409_),
    .A1(net9691),
    .A2(net10028));
 sg13g2_nand2_1 _18337_ (.Y(_11065_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][24] ),
    .B(net10028));
 sg13g2_o21ai_1 _18338_ (.B1(_11065_),
    .Y(_01410_),
    .A1(net9686),
    .A2(net10028));
 sg13g2_nand2_1 _18339_ (.Y(_11066_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][25] ),
    .B(net10030));
 sg13g2_o21ai_1 _18340_ (.B1(_11066_),
    .Y(_01411_),
    .A1(net9680),
    .A2(net10030));
 sg13g2_buf_16 clkbuf_leaf_226_clk (.X(clknet_leaf_226_clk),
    .A(clknet_8_66_0_clk));
 sg13g2_nand2_1 _18342_ (.Y(_11068_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][26] ),
    .B(net10031));
 sg13g2_o21ai_1 _18343_ (.B1(_11068_),
    .Y(_01412_),
    .A1(net9677),
    .A2(net10031));
 sg13g2_nand2_1 _18344_ (.Y(_11069_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][27] ),
    .B(net10031));
 sg13g2_o21ai_1 _18345_ (.B1(_11069_),
    .Y(_01413_),
    .A1(net9649),
    .A2(net10031));
 sg13g2_buf_2 place10475 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[6] ),
    .X(net10475));
 sg13g2_nand2_1 _18347_ (.Y(_11071_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][28] ),
    .B(net10031));
 sg13g2_o21ai_1 _18348_ (.B1(_11071_),
    .Y(_01414_),
    .A1(net9648),
    .A2(net10031));
 sg13g2_nand2_1 _18349_ (.Y(_11072_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][29] ),
    .B(net10030));
 sg13g2_o21ai_1 _18350_ (.B1(_11072_),
    .Y(_01415_),
    .A1(net9644),
    .A2(net10030));
 sg13g2_nand2_1 _18351_ (.Y(_11073_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][2] ),
    .B(net10026));
 sg13g2_o21ai_1 _18352_ (.B1(_11073_),
    .Y(_01416_),
    .A1(net10223),
    .A2(net10026));
 sg13g2_nand2_1 _18353_ (.Y(_11074_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][30] ),
    .B(net10029));
 sg13g2_o21ai_1 _18354_ (.B1(_11074_),
    .Y(_01417_),
    .A1(net9640),
    .A2(net10029));
 sg13g2_nand2_1 _18355_ (.Y(_11075_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][31] ),
    .B(net10029));
 sg13g2_o21ai_1 _18356_ (.B1(_11075_),
    .Y(_01418_),
    .A1(net9634),
    .A2(net10029));
 sg13g2_nand2_1 _18357_ (.Y(_11076_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][3] ),
    .B(net10025));
 sg13g2_o21ai_1 _18358_ (.B1(_11076_),
    .Y(_01419_),
    .A1(net10218),
    .A2(net10025));
 sg13g2_nand2_1 _18359_ (.Y(_11077_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][4] ),
    .B(net10027));
 sg13g2_o21ai_1 _18360_ (.B1(_11077_),
    .Y(_01420_),
    .A1(_10080_),
    .A2(net10027));
 sg13g2_nand2_1 _18361_ (.Y(_11078_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][5] ),
    .B(net10026));
 sg13g2_o21ai_1 _18362_ (.B1(_11078_),
    .Y(_01421_),
    .A1(net10174),
    .A2(net10026));
 sg13g2_nand2_1 _18363_ (.Y(_11079_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][6] ),
    .B(net10024));
 sg13g2_o21ai_1 _18364_ (.B1(_11079_),
    .Y(_01422_),
    .A1(_10095_),
    .A2(net10024));
 sg13g2_nand2_1 _18365_ (.Y(_11080_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][7] ),
    .B(net10024));
 sg13g2_o21ai_1 _18366_ (.B1(_11080_),
    .Y(_01423_),
    .A1(_10103_),
    .A2(net10024));
 sg13g2_nand2_1 _18367_ (.Y(_11081_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][8] ),
    .B(_11043_));
 sg13g2_o21ai_1 _18368_ (.B1(_11081_),
    .Y(_01424_),
    .A1(_10111_),
    .A2(_11043_));
 sg13g2_nand2_1 _18369_ (.Y(_11082_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][9] ),
    .B(net10024));
 sg13g2_o21ai_1 _18370_ (.B1(_11082_),
    .Y(_01425_),
    .A1(_10119_),
    .A2(net10024));
 sg13g2_nand2_2 _18371_ (.Y(_11083_),
    .A(_10124_),
    .B(_10890_));
 sg13g2_buf_2 place10473 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[9] ),
    .X(net10473));
 sg13g2_buf_2 place10527 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[6] ),
    .X(net10527));
 sg13g2_buf_2 place10571 (.A(net10568),
    .X(net10571));
 sg13g2_nand2_1 _18375_ (.Y(_11087_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][0] ),
    .B(_11083_));
 sg13g2_o21ai_1 _18376_ (.B1(_11087_),
    .Y(_01426_),
    .A1(net10279),
    .A2(_11083_));
 sg13g2_nand2_1 _18377_ (.Y(_11088_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][10] ),
    .B(net9866));
 sg13g2_o21ai_1 _18378_ (.B1(_11088_),
    .Y(_01427_),
    .A1(net10130),
    .A2(net9866));
 sg13g2_nand2_1 _18379_ (.Y(_11089_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][11] ),
    .B(net9869));
 sg13g2_o21ai_1 _18380_ (.B1(_11089_),
    .Y(_01428_),
    .A1(net9984),
    .A2(net9869));
 sg13g2_nand2_1 _18381_ (.Y(_11090_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][12] ),
    .B(net9863));
 sg13g2_o21ai_1 _18382_ (.B1(_11090_),
    .Y(_01429_),
    .A1(_09885_),
    .A2(net9863));
 sg13g2_nand2_1 _18383_ (.Y(_11091_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][13] ),
    .B(net9862));
 sg13g2_o21ai_1 _18384_ (.B1(_11091_),
    .Y(_01430_),
    .A1(_09894_),
    .A2(net9862));
 sg13g2_nand2_1 _18385_ (.Y(_11092_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][14] ),
    .B(net9868));
 sg13g2_o21ai_1 _18386_ (.B1(_11092_),
    .Y(_01431_),
    .A1(net9798),
    .A2(net9868));
 sg13g2_nand2_1 _18387_ (.Y(_11093_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][15] ),
    .B(net9866));
 sg13g2_o21ai_1 _18388_ (.B1(_11093_),
    .Y(_01432_),
    .A1(_09911_),
    .A2(net9866));
 sg13g2_nand2_1 _18389_ (.Y(_11094_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][16] ),
    .B(net9865));
 sg13g2_o21ai_1 _18390_ (.B1(_11094_),
    .Y(_01433_),
    .A1(_09919_),
    .A2(net9865));
 sg13g2_buf_2 place10488 (.A(\u_ac_controller_soc_inst.u_picorv32.reg_pc[8] ),
    .X(net10488));
 sg13g2_nand2_1 _18392_ (.Y(_11096_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][17] ),
    .B(net9862));
 sg13g2_o21ai_1 _18393_ (.B1(_11096_),
    .Y(_01434_),
    .A1(_09928_),
    .A2(net9862));
 sg13g2_nand2_1 _18394_ (.Y(_11097_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][18] ),
    .B(net9864));
 sg13g2_o21ai_1 _18395_ (.B1(_11097_),
    .Y(_01435_),
    .A1(net9737),
    .A2(net9864));
 sg13g2_buf_16 clkbuf_leaf_231_clk (.X(clknet_leaf_231_clk),
    .A(clknet_8_65_0_clk));
 sg13g2_nand2_1 _18397_ (.Y(_11099_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][19] ),
    .B(net9871));
 sg13g2_o21ai_1 _18398_ (.B1(_11099_),
    .Y(_01436_),
    .A1(net9725),
    .A2(net9871));
 sg13g2_nand2_1 _18399_ (.Y(_11100_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][1] ),
    .B(net9862));
 sg13g2_o21ai_1 _18400_ (.B1(_11100_),
    .Y(_01437_),
    .A1(_09954_),
    .A2(net9862));
 sg13g2_nand2_1 _18401_ (.Y(_11101_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][20] ),
    .B(net9867));
 sg13g2_o21ai_1 _18402_ (.B1(_11101_),
    .Y(_01438_),
    .A1(net9716),
    .A2(net9867));
 sg13g2_nand2_1 _18403_ (.Y(_11102_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][21] ),
    .B(net9864));
 sg13g2_o21ai_1 _18404_ (.B1(_11102_),
    .Y(_01439_),
    .A1(net9712),
    .A2(net9864));
 sg13g2_nand2_1 _18405_ (.Y(_11103_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][22] ),
    .B(net9867));
 sg13g2_o21ai_1 _18406_ (.B1(_11103_),
    .Y(_01440_),
    .A1(net9694),
    .A2(net9867));
 sg13g2_nand2_1 _18407_ (.Y(_11104_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][23] ),
    .B(net9867));
 sg13g2_o21ai_1 _18408_ (.B1(_11104_),
    .Y(_01441_),
    .A1(net9691),
    .A2(net9867));
 sg13g2_nand2_1 _18409_ (.Y(_11105_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][24] ),
    .B(net9867));
 sg13g2_o21ai_1 _18410_ (.B1(_11105_),
    .Y(_01442_),
    .A1(net9686),
    .A2(net9867));
 sg13g2_nand2_1 _18411_ (.Y(_11106_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][25] ),
    .B(net9870));
 sg13g2_o21ai_1 _18412_ (.B1(_11106_),
    .Y(_01443_),
    .A1(net9680),
    .A2(net9870));
 sg13g2_buf_16 clkbuf_leaf_229_clk (.X(clknet_leaf_229_clk),
    .A(clknet_8_67_0_clk));
 sg13g2_nand2_1 _18414_ (.Y(_11108_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][26] ),
    .B(net9871));
 sg13g2_o21ai_1 _18415_ (.B1(_11108_),
    .Y(_01444_),
    .A1(net9677),
    .A2(net9871));
 sg13g2_nand2_1 _18416_ (.Y(_11109_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][27] ),
    .B(net9871));
 sg13g2_o21ai_1 _18417_ (.B1(_11109_),
    .Y(_01445_),
    .A1(net9649),
    .A2(net9871));
 sg13g2_buf_2 place10468 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[6] ),
    .X(net10468));
 sg13g2_nand2_1 _18419_ (.Y(_11111_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][28] ),
    .B(net9871));
 sg13g2_o21ai_1 _18420_ (.B1(_11111_),
    .Y(_01446_),
    .A1(net9648),
    .A2(net9871));
 sg13g2_nand2_1 _18421_ (.Y(_11112_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][29] ),
    .B(net9869));
 sg13g2_o21ai_1 _18422_ (.B1(_11112_),
    .Y(_01447_),
    .A1(net9644),
    .A2(net9869));
 sg13g2_nand2_1 _18423_ (.Y(_11113_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][2] ),
    .B(net9866));
 sg13g2_o21ai_1 _18424_ (.B1(_11113_),
    .Y(_01448_),
    .A1(net10222),
    .A2(net9866));
 sg13g2_nand2_1 _18425_ (.Y(_11114_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][30] ),
    .B(net9869));
 sg13g2_o21ai_1 _18426_ (.B1(_11114_),
    .Y(_01449_),
    .A1(net9639),
    .A2(net9868));
 sg13g2_nand2_1 _18427_ (.Y(_11115_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][31] ),
    .B(net9868));
 sg13g2_o21ai_1 _18428_ (.B1(_11115_),
    .Y(_01450_),
    .A1(net9634),
    .A2(net9868));
 sg13g2_nand2_1 _18429_ (.Y(_11116_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][3] ),
    .B(net9865));
 sg13g2_o21ai_1 _18430_ (.B1(_11116_),
    .Y(_01451_),
    .A1(net10218),
    .A2(net9865));
 sg13g2_nand2_1 _18431_ (.Y(_11117_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][4] ),
    .B(net9864));
 sg13g2_o21ai_1 _18432_ (.B1(_11117_),
    .Y(_01452_),
    .A1(_10080_),
    .A2(net9864));
 sg13g2_nand2_1 _18433_ (.Y(_11118_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][5] ),
    .B(net9866));
 sg13g2_o21ai_1 _18434_ (.B1(_11118_),
    .Y(_01453_),
    .A1(net10176),
    .A2(net9866));
 sg13g2_nand2_1 _18435_ (.Y(_11119_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][6] ),
    .B(net9863));
 sg13g2_o21ai_1 _18436_ (.B1(_11119_),
    .Y(_01454_),
    .A1(_10095_),
    .A2(net9863));
 sg13g2_nand2_1 _18437_ (.Y(_11120_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][7] ),
    .B(net9863));
 sg13g2_o21ai_1 _18438_ (.B1(_11120_),
    .Y(_01455_),
    .A1(_10103_),
    .A2(net9863));
 sg13g2_nand2_1 _18439_ (.Y(_11121_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][8] ),
    .B(net9868));
 sg13g2_o21ai_1 _18440_ (.B1(_11121_),
    .Y(_01456_),
    .A1(_10111_),
    .A2(_11083_));
 sg13g2_nand2_1 _18441_ (.Y(_11122_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][9] ),
    .B(net9863));
 sg13g2_o21ai_1 _18442_ (.B1(_11122_),
    .Y(_01457_),
    .A1(_10119_),
    .A2(net9863));
 sg13g2_nand2_2 _18443_ (.Y(_11123_),
    .A(_10124_),
    .B(_10168_));
 sg13g2_buf_2 place10634 (.A(net10633),
    .X(net10634));
 sg13g2_buf_16 clkbuf_leaf_228_clk (.X(clknet_leaf_228_clk),
    .A(clknet_8_67_0_clk));
 sg13g2_buf_16 clkbuf_leaf_227_clk (.X(clknet_leaf_227_clk),
    .A(clknet_8_66_0_clk));
 sg13g2_nand2_1 _18447_ (.Y(_11127_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][0] ),
    .B(net9858));
 sg13g2_o21ai_1 _18448_ (.B1(_11127_),
    .Y(_01458_),
    .A1(net10279),
    .A2(_11123_));
 sg13g2_nand2_1 _18449_ (.Y(_11128_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][10] ),
    .B(net9857));
 sg13g2_o21ai_1 _18450_ (.B1(_11128_),
    .Y(_01459_),
    .A1(net10132),
    .A2(net9857));
 sg13g2_nand2_1 _18451_ (.Y(_11129_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][11] ),
    .B(net9855));
 sg13g2_o21ai_1 _18452_ (.B1(_11129_),
    .Y(_01460_),
    .A1(net9983),
    .A2(net9855));
 sg13g2_nand2_1 _18453_ (.Y(_11130_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][12] ),
    .B(net9860));
 sg13g2_o21ai_1 _18454_ (.B1(_11130_),
    .Y(_01461_),
    .A1(net9803),
    .A2(net9860));
 sg13g2_nand2_1 _18455_ (.Y(_11131_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][13] ),
    .B(net9859));
 sg13g2_o21ai_1 _18456_ (.B1(_11131_),
    .Y(_01462_),
    .A1(net9980),
    .A2(net9859));
 sg13g2_nand2_1 _18457_ (.Y(_11132_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][14] ),
    .B(net9853));
 sg13g2_o21ai_1 _18458_ (.B1(_11132_),
    .Y(_01463_),
    .A1(net9796),
    .A2(net9853));
 sg13g2_nand2_1 _18459_ (.Y(_11133_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][15] ),
    .B(net9861));
 sg13g2_o21ai_1 _18460_ (.B1(_11133_),
    .Y(_01464_),
    .A1(net9792),
    .A2(net9861));
 sg13g2_nand2_1 _18461_ (.Y(_11134_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][16] ),
    .B(net9858));
 sg13g2_o21ai_1 _18462_ (.B1(_11134_),
    .Y(_01465_),
    .A1(net9745),
    .A2(net9858));
 sg13g2_buf_2 place10462 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_qspi ),
    .X(net10462));
 sg13g2_nand2_1 _18464_ (.Y(_11136_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][17] ),
    .B(net9858));
 sg13g2_o21ai_1 _18465_ (.B1(_11136_),
    .Y(_01466_),
    .A1(net9739),
    .A2(net9858));
 sg13g2_nand2_1 _18466_ (.Y(_11137_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][18] ),
    .B(_11123_));
 sg13g2_o21ai_1 _18467_ (.B1(_11137_),
    .Y(_01467_),
    .A1(net9737),
    .A2(_11123_));
 sg13g2_buf_16 clkbuf_leaf_233_clk (.X(clknet_leaf_233_clk),
    .A(clknet_8_64_0_clk));
 sg13g2_nand2_1 _18469_ (.Y(_11139_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][19] ),
    .B(net9856));
 sg13g2_o21ai_1 _18470_ (.B1(_11139_),
    .Y(_01468_),
    .A1(net9721),
    .A2(net9856));
 sg13g2_nand2_1 _18471_ (.Y(_11140_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][1] ),
    .B(net9859));
 sg13g2_o21ai_1 _18472_ (.B1(_11140_),
    .Y(_01469_),
    .A1(net10229),
    .A2(net9859));
 sg13g2_nand2_1 _18473_ (.Y(_11141_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][20] ),
    .B(net9857));
 sg13g2_o21ai_1 _18474_ (.B1(_11141_),
    .Y(_01470_),
    .A1(net9720),
    .A2(net9857));
 sg13g2_nand2_1 _18475_ (.Y(_11142_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][21] ),
    .B(net9857));
 sg13g2_o21ai_1 _18476_ (.B1(_11142_),
    .Y(_01471_),
    .A1(net9715),
    .A2(net9857));
 sg13g2_nand2_1 _18477_ (.Y(_11143_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][22] ),
    .B(net9854));
 sg13g2_o21ai_1 _18478_ (.B1(_11143_),
    .Y(_01472_),
    .A1(_09980_),
    .A2(net9854));
 sg13g2_nand2_1 _18479_ (.Y(_11144_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][23] ),
    .B(net9854));
 sg13g2_o21ai_1 _18480_ (.B1(_11144_),
    .Y(_01473_),
    .A1(_09988_),
    .A2(net9854));
 sg13g2_nand2_1 _18481_ (.Y(_11145_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][24] ),
    .B(net9854));
 sg13g2_o21ai_1 _18482_ (.B1(_11145_),
    .Y(_01474_),
    .A1(_09997_),
    .A2(net9854));
 sg13g2_nand2_1 _18483_ (.Y(_11146_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][25] ),
    .B(net9855));
 sg13g2_o21ai_1 _18484_ (.B1(_11146_),
    .Y(_01475_),
    .A1(net9681),
    .A2(net9855));
 sg13g2_buf_16 clkbuf_leaf_232_clk (.X(clknet_leaf_232_clk),
    .A(clknet_8_64_0_clk));
 sg13g2_nand2_1 _18486_ (.Y(_11148_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][26] ),
    .B(net9856));
 sg13g2_o21ai_1 _18487_ (.B1(_11148_),
    .Y(_01476_),
    .A1(net9674),
    .A2(net9856));
 sg13g2_nand2_1 _18488_ (.Y(_11149_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][27] ),
    .B(net9855));
 sg13g2_o21ai_1 _18489_ (.B1(_11149_),
    .Y(_01477_),
    .A1(net9652),
    .A2(net9855));
 sg13g2_buf_2 place10469 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[2] ),
    .X(net10469));
 sg13g2_nand2_1 _18491_ (.Y(_11151_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][28] ),
    .B(net9856));
 sg13g2_o21ai_1 _18492_ (.B1(_11151_),
    .Y(_01478_),
    .A1(net9647),
    .A2(net9856));
 sg13g2_nand2_1 _18493_ (.Y(_11152_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][29] ),
    .B(net9855));
 sg13g2_o21ai_1 _18494_ (.B1(_11152_),
    .Y(_01479_),
    .A1(net9641),
    .A2(net9855));
 sg13g2_nand2_1 _18495_ (.Y(_11153_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][2] ),
    .B(net9861));
 sg13g2_o21ai_1 _18496_ (.B1(_11153_),
    .Y(_01480_),
    .A1(_10047_),
    .A2(net9861));
 sg13g2_nand2_1 _18497_ (.Y(_11154_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][30] ),
    .B(net9853));
 sg13g2_o21ai_1 _18498_ (.B1(_11154_),
    .Y(_01481_),
    .A1(_10056_),
    .A2(net9853));
 sg13g2_nand2_1 _18499_ (.Y(_11155_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][31] ),
    .B(net9856));
 sg13g2_o21ai_1 _18500_ (.B1(_11155_),
    .Y(_01482_),
    .A1(net9632),
    .A2(net9856));
 sg13g2_nand2_1 _18501_ (.Y(_11156_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][3] ),
    .B(net9861));
 sg13g2_o21ai_1 _18502_ (.B1(_11156_),
    .Y(_01483_),
    .A1(net10221),
    .A2(net9861));
 sg13g2_nand2_1 _18503_ (.Y(_11157_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][4] ),
    .B(net9857));
 sg13g2_o21ai_1 _18504_ (.B1(_11157_),
    .Y(_01484_),
    .A1(net10181),
    .A2(net9857));
 sg13g2_nand2_1 _18505_ (.Y(_11158_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][5] ),
    .B(net9861));
 sg13g2_o21ai_1 _18506_ (.B1(_11158_),
    .Y(_01485_),
    .A1(net10177),
    .A2(net9861));
 sg13g2_nand2_1 _18507_ (.Y(_11159_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][6] ),
    .B(net9860));
 sg13g2_o21ai_1 _18508_ (.B1(_11159_),
    .Y(_01486_),
    .A1(net10172),
    .A2(net9860));
 sg13g2_nand2_1 _18509_ (.Y(_11160_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][7] ),
    .B(net9860));
 sg13g2_o21ai_1 _18510_ (.B1(_11160_),
    .Y(_01487_),
    .A1(net10169),
    .A2(net9860));
 sg13g2_nand2_1 _18511_ (.Y(_11161_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][8] ),
    .B(net9853));
 sg13g2_o21ai_1 _18512_ (.B1(_11161_),
    .Y(_01488_),
    .A1(net10126),
    .A2(net9853));
 sg13g2_nand2_1 _18513_ (.Y(_11162_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][9] ),
    .B(net9860));
 sg13g2_o21ai_1 _18514_ (.B1(_11162_),
    .Y(_01489_),
    .A1(net9977),
    .A2(net9860));
 sg13g2_nor3_2 _18515_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[4] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_rd[3] ),
    .C(_00084_),
    .Y(_11163_));
 sg13g2_nand2_2 _18516_ (.Y(_11164_),
    .A(_10169_),
    .B(_11163_));
 sg13g2_buf_2 place10474 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[8] ),
    .X(net10474));
 sg13g2_buf_2 place10461 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.resetn ),
    .X(net10461));
 sg13g2_buf_2 place10467 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk ),
    .X(net10467));
 sg13g2_nand2_1 _18520_ (.Y(_11168_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][0] ),
    .B(_11164_));
 sg13g2_o21ai_1 _18521_ (.B1(_11168_),
    .Y(_01490_),
    .A1(net10279),
    .A2(_11164_));
 sg13g2_nand2_1 _18522_ (.Y(_11169_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][10] ),
    .B(net10017));
 sg13g2_o21ai_1 _18523_ (.B1(_11169_),
    .Y(_01491_),
    .A1(net10133),
    .A2(net10017));
 sg13g2_nand2_1 _18524_ (.Y(_11170_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][11] ),
    .B(net10021));
 sg13g2_o21ai_1 _18525_ (.B1(_11170_),
    .Y(_01492_),
    .A1(net9982),
    .A2(net10019));
 sg13g2_nand2_1 _18526_ (.Y(_11171_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][12] ),
    .B(net10014));
 sg13g2_o21ai_1 _18527_ (.B1(_11171_),
    .Y(_01493_),
    .A1(net9803),
    .A2(net10015));
 sg13g2_nand2_1 _18528_ (.Y(_11172_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][13] ),
    .B(net10014));
 sg13g2_o21ai_1 _18529_ (.B1(_11172_),
    .Y(_01494_),
    .A1(net9979),
    .A2(net10014));
 sg13g2_nand2_1 _18530_ (.Y(_11173_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][14] ),
    .B(net10018));
 sg13g2_o21ai_1 _18531_ (.B1(_11173_),
    .Y(_01495_),
    .A1(net9796),
    .A2(net10018));
 sg13g2_nand2_1 _18532_ (.Y(_11174_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][15] ),
    .B(net10017));
 sg13g2_o21ai_1 _18533_ (.B1(_11174_),
    .Y(_01496_),
    .A1(net9794),
    .A2(net10017));
 sg13g2_nand2_1 _18534_ (.Y(_11175_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][16] ),
    .B(_11164_));
 sg13g2_o21ai_1 _18535_ (.B1(_11175_),
    .Y(_01497_),
    .A1(net9743),
    .A2(net10013));
 sg13g2_buf_2 place10565 (.A(net10564),
    .X(net10565));
 sg13g2_nand2_1 _18537_ (.Y(_11177_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][17] ),
    .B(net10013));
 sg13g2_o21ai_1 _18538_ (.B1(_11177_),
    .Y(_01498_),
    .A1(net9740),
    .A2(net10013));
 sg13g2_nand2_1 _18539_ (.Y(_11178_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][18] ),
    .B(_11164_));
 sg13g2_o21ai_1 _18540_ (.B1(_11178_),
    .Y(_01499_),
    .A1(net9737),
    .A2(_11164_));
 sg13g2_buf_2 place10597 (.A(net10596),
    .X(net10597));
 sg13g2_nand2_1 _18542_ (.Y(_11180_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][19] ),
    .B(net10022));
 sg13g2_o21ai_1 _18543_ (.B1(_11180_),
    .Y(_01500_),
    .A1(net9722),
    .A2(net10022));
 sg13g2_nand2_1 _18544_ (.Y(_11181_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][1] ),
    .B(net10014));
 sg13g2_o21ai_1 _18545_ (.B1(_11181_),
    .Y(_01501_),
    .A1(net10228),
    .A2(net10014));
 sg13g2_nand2_1 _18546_ (.Y(_11182_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][20] ),
    .B(net10016));
 sg13g2_o21ai_1 _18547_ (.B1(_11182_),
    .Y(_01502_),
    .A1(net9720),
    .A2(net10016));
 sg13g2_nand2_1 _18548_ (.Y(_11183_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][21] ),
    .B(net10016));
 sg13g2_o21ai_1 _18549_ (.B1(_11183_),
    .Y(_01503_),
    .A1(net9715),
    .A2(net10016));
 sg13g2_nand2_1 _18550_ (.Y(_11184_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][22] ),
    .B(net10019));
 sg13g2_o21ai_1 _18551_ (.B1(_11184_),
    .Y(_01504_),
    .A1(net9693),
    .A2(net10019));
 sg13g2_nand2_1 _18552_ (.Y(_11185_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][23] ),
    .B(net10019));
 sg13g2_o21ai_1 _18553_ (.B1(_11185_),
    .Y(_01505_),
    .A1(net9689),
    .A2(net10019));
 sg13g2_nand2_1 _18554_ (.Y(_11186_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][24] ),
    .B(net10019));
 sg13g2_o21ai_1 _18555_ (.B1(_11186_),
    .Y(_01506_),
    .A1(net9688),
    .A2(net10019));
 sg13g2_nand2_1 _18556_ (.Y(_11187_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][25] ),
    .B(net10020));
 sg13g2_o21ai_1 _18557_ (.B1(_11187_),
    .Y(_01507_),
    .A1(_10005_),
    .A2(net10020));
 sg13g2_buf_2 place10466 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr ),
    .X(net10466));
 sg13g2_nand2_1 _18559_ (.Y(_11189_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][26] ),
    .B(net10021));
 sg13g2_o21ai_1 _18560_ (.B1(_11189_),
    .Y(_01508_),
    .A1(net9676),
    .A2(net10021));
 sg13g2_nand2_1 _18561_ (.Y(_11190_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][27] ),
    .B(net10020));
 sg13g2_o21ai_1 _18562_ (.B1(_11190_),
    .Y(_01509_),
    .A1(net9650),
    .A2(net10020));
 sg13g2_buf_2 place10464 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_qspi ),
    .X(net10464));
 sg13g2_nand2_1 _18564_ (.Y(_11192_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][28] ),
    .B(net10022));
 sg13g2_o21ai_1 _18565_ (.B1(_11192_),
    .Y(_01510_),
    .A1(net9645),
    .A2(net10022));
 sg13g2_nand2_1 _18566_ (.Y(_11193_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][29] ),
    .B(net10020));
 sg13g2_o21ai_1 _18567_ (.B1(_11193_),
    .Y(_01511_),
    .A1(net9642),
    .A2(net10020));
 sg13g2_nand2_1 _18568_ (.Y(_11194_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][2] ),
    .B(net10013));
 sg13g2_o21ai_1 _18569_ (.B1(_11194_),
    .Y(_01512_),
    .A1(_10047_),
    .A2(net10013));
 sg13g2_nand2_1 _18570_ (.Y(_11195_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][30] ),
    .B(net10021));
 sg13g2_o21ai_1 _18571_ (.B1(_11195_),
    .Y(_01513_),
    .A1(_10056_),
    .A2(net10022));
 sg13g2_nand2_1 _18572_ (.Y(_11196_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][31] ),
    .B(net10022));
 sg13g2_o21ai_1 _18573_ (.B1(_11196_),
    .Y(_01514_),
    .A1(net9633),
    .A2(net10022));
 sg13g2_nand2_1 _18574_ (.Y(_11197_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][3] ),
    .B(net10017));
 sg13g2_o21ai_1 _18575_ (.B1(_11197_),
    .Y(_01515_),
    .A1(net10221),
    .A2(net10017));
 sg13g2_nand2_1 _18576_ (.Y(_11198_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][4] ),
    .B(net10016));
 sg13g2_o21ai_1 _18577_ (.B1(_11198_),
    .Y(_01516_),
    .A1(net10180),
    .A2(net10016));
 sg13g2_nand2_1 _18578_ (.Y(_11199_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][5] ),
    .B(net10017));
 sg13g2_o21ai_1 _18579_ (.B1(_11199_),
    .Y(_01517_),
    .A1(net10175),
    .A2(net10017));
 sg13g2_nand2_1 _18580_ (.Y(_11200_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][6] ),
    .B(net10015));
 sg13g2_o21ai_1 _18581_ (.B1(_11200_),
    .Y(_01518_),
    .A1(net10172),
    .A2(net10015));
 sg13g2_nand2_1 _18582_ (.Y(_11201_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][7] ),
    .B(net10015));
 sg13g2_o21ai_1 _18583_ (.B1(_11201_),
    .Y(_01519_),
    .A1(net10169),
    .A2(net10015));
 sg13g2_nand2_1 _18584_ (.Y(_11202_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][8] ),
    .B(net10018));
 sg13g2_o21ai_1 _18585_ (.B1(_11202_),
    .Y(_01520_),
    .A1(net10129),
    .A2(net10018));
 sg13g2_nand2_1 _18586_ (.Y(_11203_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][9] ),
    .B(net10015));
 sg13g2_o21ai_1 _18587_ (.B1(_11203_),
    .Y(_01521_),
    .A1(net9976),
    .A2(net10015));
 sg13g2_nand2_2 _18588_ (.Y(_11204_),
    .A(_10211_),
    .B(_11163_));
 sg13g2_buf_16 clkbuf_leaf_234_clk (.X(clknet_leaf_234_clk),
    .A(clknet_8_65_0_clk));
 sg13g2_buf_2 place10460 (.A(_07949_),
    .X(net10460));
 sg13g2_buf_2 place10472 (.A(net10471),
    .X(net10472));
 sg13g2_nand2_1 _18592_ (.Y(_11208_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][0] ),
    .B(net9844));
 sg13g2_o21ai_1 _18593_ (.B1(_11208_),
    .Y(_01522_),
    .A1(net10280),
    .A2(net9844));
 sg13g2_nand2_1 _18594_ (.Y(_11209_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][10] ),
    .B(net9848));
 sg13g2_o21ai_1 _18595_ (.B1(_11209_),
    .Y(_01523_),
    .A1(net10133),
    .A2(net9848));
 sg13g2_nand2_1 _18596_ (.Y(_11210_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][11] ),
    .B(net9850));
 sg13g2_o21ai_1 _18597_ (.B1(_11210_),
    .Y(_01524_),
    .A1(net9982),
    .A2(net9850));
 sg13g2_nand2_1 _18598_ (.Y(_11211_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][12] ),
    .B(net9846));
 sg13g2_o21ai_1 _18599_ (.B1(_11211_),
    .Y(_01525_),
    .A1(net9803),
    .A2(net9846));
 sg13g2_nand2_1 _18600_ (.Y(_11212_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][13] ),
    .B(net9844));
 sg13g2_o21ai_1 _18601_ (.B1(_11212_),
    .Y(_01526_),
    .A1(net9981),
    .A2(net9844));
 sg13g2_nand2_1 _18602_ (.Y(_11213_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][14] ),
    .B(net9851));
 sg13g2_o21ai_1 _18603_ (.B1(_11213_),
    .Y(_01527_),
    .A1(net9796),
    .A2(net9851));
 sg13g2_nand2_1 _18604_ (.Y(_11214_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][15] ),
    .B(net9848));
 sg13g2_o21ai_1 _18605_ (.B1(_11214_),
    .Y(_01528_),
    .A1(net9794),
    .A2(net9848));
 sg13g2_nand2_1 _18606_ (.Y(_11215_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][16] ),
    .B(net9844));
 sg13g2_o21ai_1 _18607_ (.B1(_11215_),
    .Y(_01529_),
    .A1(net9743),
    .A2(net9844));
 sg13g2_buf_2 place10575 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[18] ),
    .X(net10575));
 sg13g2_nand2_1 _18609_ (.Y(_11217_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][17] ),
    .B(net9845));
 sg13g2_o21ai_1 _18610_ (.B1(_11217_),
    .Y(_01530_),
    .A1(net9740),
    .A2(net9845));
 sg13g2_nand2_1 _18611_ (.Y(_11218_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][18] ),
    .B(_11204_));
 sg13g2_o21ai_1 _18612_ (.B1(_11218_),
    .Y(_01531_),
    .A1(net9736),
    .A2(net9844));
 sg13g2_buf_2 place10646 (.A(net10645),
    .X(net10646));
 sg13g2_nand2_1 _18614_ (.Y(_11220_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][19] ),
    .B(net9852));
 sg13g2_o21ai_1 _18615_ (.B1(_11220_),
    .Y(_01532_),
    .A1(net9722),
    .A2(net9852));
 sg13g2_nand2_1 _18616_ (.Y(_11221_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][1] ),
    .B(net9845));
 sg13g2_o21ai_1 _18617_ (.B1(_11221_),
    .Y(_01533_),
    .A1(net10228),
    .A2(net9845));
 sg13g2_nand2_1 _18618_ (.Y(_11222_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][20] ),
    .B(net9847));
 sg13g2_o21ai_1 _18619_ (.B1(_11222_),
    .Y(_01534_),
    .A1(net9720),
    .A2(net9847));
 sg13g2_nand2_1 _18620_ (.Y(_11223_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][21] ),
    .B(net9847));
 sg13g2_o21ai_1 _18621_ (.B1(_11223_),
    .Y(_01535_),
    .A1(net9715),
    .A2(net9847));
 sg13g2_nand2_1 _18622_ (.Y(_11224_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][22] ),
    .B(net9851));
 sg13g2_o21ai_1 _18623_ (.B1(_11224_),
    .Y(_01536_),
    .A1(net9693),
    .A2(net9851));
 sg13g2_nand2_1 _18624_ (.Y(_11225_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][23] ),
    .B(net9851));
 sg13g2_o21ai_1 _18625_ (.B1(_11225_),
    .Y(_01537_),
    .A1(net9689),
    .A2(net9851));
 sg13g2_nand2_1 _18626_ (.Y(_11226_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][24] ),
    .B(net9851));
 sg13g2_o21ai_1 _18627_ (.B1(_11226_),
    .Y(_01538_),
    .A1(net9685),
    .A2(net9851));
 sg13g2_nand2_1 _18628_ (.Y(_11227_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][25] ),
    .B(net9850));
 sg13g2_o21ai_1 _18629_ (.B1(_11227_),
    .Y(_01539_),
    .A1(_10005_),
    .A2(net9850));
 sg13g2_buf_2 place10463 (.A(net10462),
    .X(net10463));
 sg13g2_nand2_1 _18631_ (.Y(_11229_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][26] ),
    .B(net9849));
 sg13g2_o21ai_1 _18632_ (.B1(_11229_),
    .Y(_01540_),
    .A1(net9676),
    .A2(net9849));
 sg13g2_nand2_1 _18633_ (.Y(_11230_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][27] ),
    .B(net9850));
 sg13g2_o21ai_1 _18634_ (.B1(_11230_),
    .Y(_01541_),
    .A1(net9650),
    .A2(net9850));
 sg13g2_buf_2 place10465 (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_qspi ),
    .X(net10465));
 sg13g2_nand2_1 _18636_ (.Y(_11232_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][28] ),
    .B(net9852));
 sg13g2_o21ai_1 _18637_ (.B1(_11232_),
    .Y(_01542_),
    .A1(net9645),
    .A2(net9852));
 sg13g2_nand2_1 _18638_ (.Y(_11233_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][29] ),
    .B(net9850));
 sg13g2_o21ai_1 _18639_ (.B1(_11233_),
    .Y(_01543_),
    .A1(net9642),
    .A2(net9850));
 sg13g2_nand2_1 _18640_ (.Y(_11234_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][2] ),
    .B(net9845));
 sg13g2_o21ai_1 _18641_ (.B1(_11234_),
    .Y(_01544_),
    .A1(_10047_),
    .A2(net9845));
 sg13g2_nand2_1 _18642_ (.Y(_11235_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][30] ),
    .B(net9849));
 sg13g2_o21ai_1 _18643_ (.B1(_11235_),
    .Y(_01545_),
    .A1(_10056_),
    .A2(net9852));
 sg13g2_nand2_1 _18644_ (.Y(_11236_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][31] ),
    .B(net9852));
 sg13g2_o21ai_1 _18645_ (.B1(_11236_),
    .Y(_01546_),
    .A1(net9632),
    .A2(net9852));
 sg13g2_nand2_1 _18646_ (.Y(_11237_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][3] ),
    .B(net9848));
 sg13g2_o21ai_1 _18647_ (.B1(_11237_),
    .Y(_01547_),
    .A1(net10221),
    .A2(net9848));
 sg13g2_nand2_1 _18648_ (.Y(_11238_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][4] ),
    .B(net9847));
 sg13g2_o21ai_1 _18649_ (.B1(_11238_),
    .Y(_01548_),
    .A1(net10181),
    .A2(net9847));
 sg13g2_nand2_1 _18650_ (.Y(_11239_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][5] ),
    .B(net9848));
 sg13g2_o21ai_1 _18651_ (.B1(_11239_),
    .Y(_01549_),
    .A1(net10177),
    .A2(net9848));
 sg13g2_nand2_1 _18652_ (.Y(_11240_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][6] ),
    .B(net9846));
 sg13g2_o21ai_1 _18653_ (.B1(_11240_),
    .Y(_01550_),
    .A1(net10172),
    .A2(net9846));
 sg13g2_nand2_1 _18654_ (.Y(_11241_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][7] ),
    .B(net9846));
 sg13g2_o21ai_1 _18655_ (.B1(_11241_),
    .Y(_01551_),
    .A1(net10169),
    .A2(net9846));
 sg13g2_nand2_1 _18656_ (.Y(_11242_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][8] ),
    .B(net9849));
 sg13g2_o21ai_1 _18657_ (.B1(_11242_),
    .Y(_01552_),
    .A1(net10129),
    .A2(net9849));
 sg13g2_nand2_1 _18658_ (.Y(_11243_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][9] ),
    .B(net9846));
 sg13g2_o21ai_1 _18659_ (.B1(_11243_),
    .Y(_01553_),
    .A1(net9976),
    .A2(net9846));
 sg13g2_nand2_2 _18660_ (.Y(_11244_),
    .A(_09850_),
    .B(_11163_));
 sg13g2_buf_16 clkbuf_leaf_241_clk (.X(clknet_leaf_241_clk),
    .A(clknet_8_70_0_clk));
 sg13g2_buf_16 clkbuf_leaf_240_clk (.X(clknet_leaf_240_clk),
    .A(clknet_8_65_0_clk));
 sg13g2_buf_2 place10457 (.A(net10456),
    .X(net10457));
 sg13g2_nand2_1 _18664_ (.Y(_11248_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][0] ),
    .B(_11244_));
 sg13g2_o21ai_1 _18665_ (.B1(_11248_),
    .Y(_01554_),
    .A1(net10279),
    .A2(_11244_));
 sg13g2_nand2_1 _18666_ (.Y(_11249_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][10] ),
    .B(net10006));
 sg13g2_o21ai_1 _18667_ (.B1(_11249_),
    .Y(_01555_),
    .A1(net10133),
    .A2(net10006));
 sg13g2_nand2_1 _18668_ (.Y(_11250_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][11] ),
    .B(net10007));
 sg13g2_o21ai_1 _18669_ (.B1(_11250_),
    .Y(_01556_),
    .A1(net9982),
    .A2(net10007));
 sg13g2_nand2_1 _18670_ (.Y(_11251_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][12] ),
    .B(net10012));
 sg13g2_o21ai_1 _18671_ (.B1(_11251_),
    .Y(_01557_),
    .A1(net9803),
    .A2(net10012));
 sg13g2_nand2_1 _18672_ (.Y(_11252_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][13] ),
    .B(_11244_));
 sg13g2_o21ai_1 _18673_ (.B1(_11252_),
    .Y(_01558_),
    .A1(net9981),
    .A2(_11244_));
 sg13g2_nand2_1 _18674_ (.Y(_11253_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][14] ),
    .B(net10007));
 sg13g2_o21ai_1 _18675_ (.B1(_11253_),
    .Y(_01559_),
    .A1(net9796),
    .A2(net10007));
 sg13g2_nand2_1 _18676_ (.Y(_11254_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][15] ),
    .B(net10006));
 sg13g2_o21ai_1 _18677_ (.B1(_11254_),
    .Y(_01560_),
    .A1(net9794),
    .A2(net10006));
 sg13g2_nand2_1 _18678_ (.Y(_11255_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][16] ),
    .B(_11244_));
 sg13g2_o21ai_1 _18679_ (.B1(_11255_),
    .Y(_01561_),
    .A1(net9743),
    .A2(_11244_));
 sg13g2_buf_2 place10665 (.A(net10664),
    .X(net10665));
 sg13g2_nand2_1 _18681_ (.Y(_11257_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][17] ),
    .B(net10011));
 sg13g2_o21ai_1 _18682_ (.B1(_11257_),
    .Y(_01562_),
    .A1(net9740),
    .A2(net10011));
 sg13g2_nand2_1 _18683_ (.Y(_11258_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][18] ),
    .B(net10005));
 sg13g2_o21ai_1 _18684_ (.B1(_11258_),
    .Y(_01563_),
    .A1(net9736),
    .A2(net10005));
 sg13g2_buf_2 place10458 (.A(net10456),
    .X(net10458));
 sg13g2_nand2_1 _18686_ (.Y(_11260_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][19] ),
    .B(net10009));
 sg13g2_o21ai_1 _18687_ (.B1(_11260_),
    .Y(_01564_),
    .A1(net9721),
    .A2(net10009));
 sg13g2_nand2_1 _18688_ (.Y(_11261_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][1] ),
    .B(net10011));
 sg13g2_o21ai_1 _18689_ (.B1(_11261_),
    .Y(_01565_),
    .A1(net10228),
    .A2(net10011));
 sg13g2_nand2_1 _18690_ (.Y(_11262_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][20] ),
    .B(net10005));
 sg13g2_o21ai_1 _18691_ (.B1(_11262_),
    .Y(_01566_),
    .A1(net9720),
    .A2(net10005));
 sg13g2_nand2_1 _18692_ (.Y(_11263_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][21] ),
    .B(net10005));
 sg13g2_o21ai_1 _18693_ (.B1(_11263_),
    .Y(_01567_),
    .A1(net9715),
    .A2(net10004));
 sg13g2_nand2_1 _18694_ (.Y(_11264_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][22] ),
    .B(net10008));
 sg13g2_o21ai_1 _18695_ (.B1(_11264_),
    .Y(_01568_),
    .A1(net9693),
    .A2(net10008));
 sg13g2_nand2_1 _18696_ (.Y(_11265_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][23] ),
    .B(net10008));
 sg13g2_o21ai_1 _18697_ (.B1(_11265_),
    .Y(_01569_),
    .A1(net9689),
    .A2(net10008));
 sg13g2_nand2_1 _18698_ (.Y(_11266_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][24] ),
    .B(net10008));
 sg13g2_o21ai_1 _18699_ (.B1(_11266_),
    .Y(_01570_),
    .A1(net9688),
    .A2(net10008));
 sg13g2_nand2_1 _18700_ (.Y(_11267_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][25] ),
    .B(net10010));
 sg13g2_o21ai_1 _18701_ (.B1(_11267_),
    .Y(_01571_),
    .A1(_10005_),
    .A2(net10010));
 sg13g2_buf_2 place10455 (.A(_08231_),
    .X(net10455));
 sg13g2_nand2_1 _18703_ (.Y(_11269_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][26] ),
    .B(net10004));
 sg13g2_o21ai_1 _18704_ (.B1(_11269_),
    .Y(_01572_),
    .A1(net9676),
    .A2(net10004));
 sg13g2_nand2_1 _18705_ (.Y(_11270_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][27] ),
    .B(net10010));
 sg13g2_o21ai_1 _18706_ (.B1(_11270_),
    .Y(_01573_),
    .A1(net9650),
    .A2(net10010));
 sg13g2_buf_16 clkbuf_leaf_238_clk (.X(clknet_leaf_238_clk),
    .A(clknet_8_70_0_clk));
 sg13g2_nand2_1 _18708_ (.Y(_11272_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][28] ),
    .B(net10009));
 sg13g2_o21ai_1 _18709_ (.B1(_11272_),
    .Y(_01574_),
    .A1(net9645),
    .A2(net10009));
 sg13g2_nand2_1 _18710_ (.Y(_11273_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][29] ),
    .B(net10010));
 sg13g2_o21ai_1 _18711_ (.B1(_11273_),
    .Y(_01575_),
    .A1(net9642),
    .A2(net10010));
 sg13g2_nand2_1 _18712_ (.Y(_11274_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][2] ),
    .B(net10011));
 sg13g2_o21ai_1 _18713_ (.B1(_11274_),
    .Y(_01576_),
    .A1(_10047_),
    .A2(net10011));
 sg13g2_nand2_1 _18714_ (.Y(_11275_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][30] ),
    .B(net10009));
 sg13g2_o21ai_1 _18715_ (.B1(_11275_),
    .Y(_01577_),
    .A1(net9639),
    .A2(net10004));
 sg13g2_nand2_1 _18716_ (.Y(_11276_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][31] ),
    .B(net10009));
 sg13g2_o21ai_1 _18717_ (.B1(_11276_),
    .Y(_01578_),
    .A1(net9633),
    .A2(net10009));
 sg13g2_nand2_1 _18718_ (.Y(_11277_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][3] ),
    .B(net10006));
 sg13g2_o21ai_1 _18719_ (.B1(_11277_),
    .Y(_01579_),
    .A1(net10221),
    .A2(net10006));
 sg13g2_nand2_1 _18720_ (.Y(_11278_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][4] ),
    .B(net10005));
 sg13g2_o21ai_1 _18721_ (.B1(_11278_),
    .Y(_01580_),
    .A1(net10180),
    .A2(net10005));
 sg13g2_nand2_1 _18722_ (.Y(_11279_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][5] ),
    .B(net10006));
 sg13g2_o21ai_1 _18723_ (.B1(_11279_),
    .Y(_01581_),
    .A1(net10177),
    .A2(net10006));
 sg13g2_nand2_1 _18724_ (.Y(_11280_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][6] ),
    .B(net10012));
 sg13g2_o21ai_1 _18725_ (.B1(_11280_),
    .Y(_01582_),
    .A1(net10172),
    .A2(net10012));
 sg13g2_nand2_1 _18726_ (.Y(_11281_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][7] ),
    .B(net10012));
 sg13g2_o21ai_1 _18727_ (.B1(_11281_),
    .Y(_01583_),
    .A1(net10169),
    .A2(net10012));
 sg13g2_nand2_1 _18728_ (.Y(_11282_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][8] ),
    .B(net10007));
 sg13g2_o21ai_1 _18729_ (.B1(_11282_),
    .Y(_01584_),
    .A1(net10129),
    .A2(net10007));
 sg13g2_nand2_1 _18730_ (.Y(_11283_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][9] ),
    .B(net10012));
 sg13g2_o21ai_1 _18731_ (.B1(_11283_),
    .Y(_01585_),
    .A1(net9976),
    .A2(net10012));
 sg13g2_nand2_2 _18732_ (.Y(_11284_),
    .A(_10124_),
    .B(_11163_));
 sg13g2_buf_16 clkbuf_leaf_235_clk (.X(clknet_leaf_235_clk),
    .A(clknet_8_65_0_clk));
 sg13g2_buf_16 clkbuf_leaf_236_clk (.X(clknet_leaf_236_clk),
    .A(clknet_8_68_0_clk));
 sg13g2_buf_16 clkbuf_leaf_244_clk (.X(clknet_leaf_244_clk),
    .A(clknet_8_76_0_clk));
 sg13g2_nand2_1 _18736_ (.Y(_11288_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][0] ),
    .B(net9835));
 sg13g2_o21ai_1 _18737_ (.B1(_11288_),
    .Y(_01586_),
    .A1(net10280),
    .A2(net9835));
 sg13g2_nand2_1 _18738_ (.Y(_11289_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][10] ),
    .B(net9839));
 sg13g2_o21ai_1 _18739_ (.B1(_11289_),
    .Y(_01587_),
    .A1(net10133),
    .A2(net9839));
 sg13g2_nand2_1 _18740_ (.Y(_11290_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][11] ),
    .B(net9842));
 sg13g2_o21ai_1 _18741_ (.B1(_11290_),
    .Y(_01588_),
    .A1(_09877_),
    .A2(net9842));
 sg13g2_nand2_1 _18742_ (.Y(_11291_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][12] ),
    .B(net9837));
 sg13g2_o21ai_1 _18743_ (.B1(_11291_),
    .Y(_01589_),
    .A1(net9803),
    .A2(net9837));
 sg13g2_nand2_1 _18744_ (.Y(_11292_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][13] ),
    .B(net9835));
 sg13g2_o21ai_1 _18745_ (.B1(_11292_),
    .Y(_01590_),
    .A1(net9981),
    .A2(net9835));
 sg13g2_nand2_1 _18746_ (.Y(_11293_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][14] ),
    .B(net9841));
 sg13g2_o21ai_1 _18747_ (.B1(_11293_),
    .Y(_01591_),
    .A1(net9796),
    .A2(net9841));
 sg13g2_nand2_1 _18748_ (.Y(_11294_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][15] ),
    .B(net9839));
 sg13g2_o21ai_1 _18749_ (.B1(_11294_),
    .Y(_01592_),
    .A1(net9794),
    .A2(net9839));
 sg13g2_nand2_1 _18750_ (.Y(_11295_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][16] ),
    .B(net9835));
 sg13g2_o21ai_1 _18751_ (.B1(_11295_),
    .Y(_01593_),
    .A1(net9743),
    .A2(net9835));
 sg13g2_buf_2 place10578 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[17] ),
    .X(net10578));
 sg13g2_nand2_1 _18753_ (.Y(_11297_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][17] ),
    .B(net9836));
 sg13g2_o21ai_1 _18754_ (.B1(_11297_),
    .Y(_01594_),
    .A1(net9740),
    .A2(net9836));
 sg13g2_nand2_1 _18755_ (.Y(_11298_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][18] ),
    .B(_11284_));
 sg13g2_o21ai_1 _18756_ (.B1(_11298_),
    .Y(_01595_),
    .A1(net9736),
    .A2(_11284_));
 sg13g2_buf_16 clkbuf_leaf_243_clk (.X(clknet_leaf_243_clk),
    .A(clknet_8_70_0_clk));
 sg13g2_nand2_1 _18758_ (.Y(_11300_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][19] ),
    .B(net9843));
 sg13g2_o21ai_1 _18759_ (.B1(_11300_),
    .Y(_01596_),
    .A1(net9721),
    .A2(net9843));
 sg13g2_nand2_1 _18760_ (.Y(_11301_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][1] ),
    .B(net9836));
 sg13g2_o21ai_1 _18761_ (.B1(_11301_),
    .Y(_01597_),
    .A1(net10229),
    .A2(net9836));
 sg13g2_nand2_1 _18762_ (.Y(_11302_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][20] ),
    .B(_11284_));
 sg13g2_o21ai_1 _18763_ (.B1(_11302_),
    .Y(_01598_),
    .A1(net9720),
    .A2(_11284_));
 sg13g2_nand2_1 _18764_ (.Y(_11303_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][21] ),
    .B(_11284_));
 sg13g2_o21ai_1 _18765_ (.B1(_11303_),
    .Y(_01599_),
    .A1(net9715),
    .A2(_11284_));
 sg13g2_nand2_1 _18766_ (.Y(_11304_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][22] ),
    .B(net9841));
 sg13g2_o21ai_1 _18767_ (.B1(_11304_),
    .Y(_01600_),
    .A1(net9694),
    .A2(net9841));
 sg13g2_nand2_1 _18768_ (.Y(_11305_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][23] ),
    .B(net9841));
 sg13g2_o21ai_1 _18769_ (.B1(_11305_),
    .Y(_01601_),
    .A1(net9689),
    .A2(net9841));
 sg13g2_nand2_1 _18770_ (.Y(_11306_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][24] ),
    .B(net9841));
 sg13g2_o21ai_1 _18771_ (.B1(_11306_),
    .Y(_01602_),
    .A1(net9688),
    .A2(net9841));
 sg13g2_nand2_1 _18772_ (.Y(_11307_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][25] ),
    .B(net9842));
 sg13g2_o21ai_1 _18773_ (.B1(_11307_),
    .Y(_01603_),
    .A1(net9681),
    .A2(net9842));
 sg13g2_buf_16 clkbuf_leaf_242_clk (.X(clknet_leaf_242_clk),
    .A(clknet_8_70_0_clk));
 sg13g2_nand2_1 _18775_ (.Y(_11309_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][26] ),
    .B(net9840));
 sg13g2_o21ai_1 _18776_ (.B1(_11309_),
    .Y(_01604_),
    .A1(net9676),
    .A2(net9840));
 sg13g2_nand2_1 _18777_ (.Y(_11310_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][27] ),
    .B(net9842));
 sg13g2_o21ai_1 _18778_ (.B1(_11310_),
    .Y(_01605_),
    .A1(net9651),
    .A2(net9842));
 sg13g2_buf_2 place10577 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[17] ),
    .X(net10577));
 sg13g2_nand2_1 _18780_ (.Y(_11312_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][28] ),
    .B(net9843));
 sg13g2_o21ai_1 _18781_ (.B1(_11312_),
    .Y(_01606_),
    .A1(net9647),
    .A2(net9843));
 sg13g2_nand2_1 _18782_ (.Y(_11313_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][29] ),
    .B(net9842));
 sg13g2_o21ai_1 _18783_ (.B1(_11313_),
    .Y(_01607_),
    .A1(net9642),
    .A2(net9842));
 sg13g2_nand2_1 _18784_ (.Y(_11314_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][2] ),
    .B(net9836));
 sg13g2_o21ai_1 _18785_ (.B1(_11314_),
    .Y(_01608_),
    .A1(_10047_),
    .A2(net9836));
 sg13g2_nand2_1 _18786_ (.Y(_11315_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][30] ),
    .B(net9843));
 sg13g2_o21ai_1 _18787_ (.B1(_11315_),
    .Y(_01609_),
    .A1(net9639),
    .A2(net9843));
 sg13g2_nand2_1 _18788_ (.Y(_11316_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][31] ),
    .B(net9843));
 sg13g2_o21ai_1 _18789_ (.B1(_11316_),
    .Y(_01610_),
    .A1(net9633),
    .A2(net9843));
 sg13g2_nand2_1 _18790_ (.Y(_11317_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][3] ),
    .B(net9839));
 sg13g2_o21ai_1 _18791_ (.B1(_11317_),
    .Y(_01611_),
    .A1(net10221),
    .A2(net9839));
 sg13g2_nand2_1 _18792_ (.Y(_11318_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][4] ),
    .B(net9838));
 sg13g2_o21ai_1 _18793_ (.B1(_11318_),
    .Y(_01612_),
    .A1(net10181),
    .A2(net9838));
 sg13g2_nand2_1 _18794_ (.Y(_11319_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][5] ),
    .B(net9839));
 sg13g2_o21ai_1 _18795_ (.B1(_11319_),
    .Y(_01613_),
    .A1(net10177),
    .A2(net9839));
 sg13g2_nand2_1 _18796_ (.Y(_11320_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][6] ),
    .B(net9837));
 sg13g2_o21ai_1 _18797_ (.B1(_11320_),
    .Y(_01614_),
    .A1(net10172),
    .A2(net9837));
 sg13g2_nand2_1 _18798_ (.Y(_11321_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][7] ),
    .B(net9837));
 sg13g2_o21ai_1 _18799_ (.B1(_11321_),
    .Y(_01615_),
    .A1(net10169),
    .A2(net9837));
 sg13g2_nand2_1 _18800_ (.Y(_11322_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][8] ),
    .B(net9840));
 sg13g2_o21ai_1 _18801_ (.B1(_11322_),
    .Y(_01616_),
    .A1(net10129),
    .A2(net9840));
 sg13g2_nand2_1 _18802_ (.Y(_11323_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][9] ),
    .B(net9837));
 sg13g2_o21ai_1 _18803_ (.B1(_11323_),
    .Y(_01617_),
    .A1(net9976),
    .A2(net9837));
 sg13g2_nand2_1 _18804_ (.Y(_11324_),
    .A(_09843_),
    .B(_10169_));
 sg13g2_buf_2 place10572 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[1] ),
    .X(net10572));
 sg13g2_buf_2 place10447 (.A(net10446),
    .X(net10447));
 sg13g2_buf_2 place10452 (.A(_08292_),
    .X(net10452));
 sg13g2_nand2_1 _18808_ (.Y(_11328_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][0] ),
    .B(net9994));
 sg13g2_o21ai_1 _18809_ (.B1(_11328_),
    .Y(_01618_),
    .A1(net10276),
    .A2(net9994));
 sg13g2_nand2_1 _18810_ (.Y(_11329_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][10] ),
    .B(net9997));
 sg13g2_o21ai_1 _18811_ (.B1(_11329_),
    .Y(_01619_),
    .A1(net10131),
    .A2(net9997));
 sg13g2_nand2_1 _18812_ (.Y(_11330_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][11] ),
    .B(net10000));
 sg13g2_o21ai_1 _18813_ (.B1(_11330_),
    .Y(_01620_),
    .A1(_09877_),
    .A2(net10000));
 sg13g2_nand2_1 _18814_ (.Y(_11331_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][12] ),
    .B(net9995));
 sg13g2_o21ai_1 _18815_ (.B1(_11331_),
    .Y(_01621_),
    .A1(net9801),
    .A2(net9995));
 sg13g2_nand2_1 _18816_ (.Y(_11332_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][13] ),
    .B(net9994));
 sg13g2_o21ai_1 _18817_ (.B1(_11332_),
    .Y(_01622_),
    .A1(net9979),
    .A2(net9994));
 sg13g2_nand2_1 _18818_ (.Y(_11333_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][14] ),
    .B(net9998));
 sg13g2_o21ai_1 _18819_ (.B1(_11333_),
    .Y(_01623_),
    .A1(net9795),
    .A2(net9998));
 sg13g2_nand2_1 _18820_ (.Y(_11334_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][15] ),
    .B(net9997));
 sg13g2_o21ai_1 _18821_ (.B1(_11334_),
    .Y(_01624_),
    .A1(net9792),
    .A2(net9997));
 sg13g2_nand2_1 _18822_ (.Y(_11335_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][16] ),
    .B(net9997));
 sg13g2_o21ai_1 _18823_ (.B1(_11335_),
    .Y(_01625_),
    .A1(net9745),
    .A2(net9997));
 sg13g2_buf_2 place10459 (.A(_08082_),
    .X(net10459));
 sg13g2_nand2_1 _18825_ (.Y(_11337_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][17] ),
    .B(net9996));
 sg13g2_o21ai_1 _18826_ (.B1(_11337_),
    .Y(_01626_),
    .A1(net9742),
    .A2(net9996));
 sg13g2_nand2_1 _18827_ (.Y(_11338_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][18] ),
    .B(net9998));
 sg13g2_o21ai_1 _18828_ (.B1(_11338_),
    .Y(_01627_),
    .A1(net9738),
    .A2(net9998));
 sg13g2_buf_2 place10453 (.A(net10452),
    .X(net10453));
 sg13g2_nand2_1 _18830_ (.Y(_11340_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][19] ),
    .B(net10001));
 sg13g2_o21ai_1 _18831_ (.B1(_11340_),
    .Y(_01628_),
    .A1(net9724),
    .A2(net10001));
 sg13g2_nand2_1 _18832_ (.Y(_11341_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][1] ),
    .B(net9994));
 sg13g2_o21ai_1 _18833_ (.B1(_11341_),
    .Y(_01629_),
    .A1(net10228),
    .A2(net9994));
 sg13g2_nand2_1 _18834_ (.Y(_11342_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][20] ),
    .B(net10003));
 sg13g2_o21ai_1 _18835_ (.B1(_11342_),
    .Y(_01630_),
    .A1(net9718),
    .A2(net10003));
 sg13g2_nand2_1 _18836_ (.Y(_11343_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][21] ),
    .B(net10003));
 sg13g2_o21ai_1 _18837_ (.B1(_11343_),
    .Y(_01631_),
    .A1(net9714),
    .A2(net10003));
 sg13g2_nand2_1 _18838_ (.Y(_11344_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][22] ),
    .B(net10002));
 sg13g2_o21ai_1 _18839_ (.B1(_11344_),
    .Y(_01632_),
    .A1(net9696),
    .A2(net10002));
 sg13g2_nand2_1 _18840_ (.Y(_11345_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][23] ),
    .B(net10002));
 sg13g2_o21ai_1 _18841_ (.B1(_11345_),
    .Y(_01633_),
    .A1(net9691),
    .A2(net10002));
 sg13g2_nand2_1 _18842_ (.Y(_11346_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][24] ),
    .B(net10002));
 sg13g2_o21ai_1 _18843_ (.B1(_11346_),
    .Y(_01634_),
    .A1(net9685),
    .A2(net10002));
 sg13g2_nand2_1 _18844_ (.Y(_11347_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][25] ),
    .B(net9999));
 sg13g2_o21ai_1 _18845_ (.B1(_11347_),
    .Y(_01635_),
    .A1(net9678),
    .A2(net9999));
 sg13g2_buf_2 place10456 (.A(_08197_),
    .X(net10456));
 sg13g2_nand2_1 _18847_ (.Y(_11349_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][26] ),
    .B(net10001));
 sg13g2_o21ai_1 _18848_ (.B1(_11349_),
    .Y(_01636_),
    .A1(net9675),
    .A2(net10001));
 sg13g2_nand2_1 _18849_ (.Y(_11350_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][27] ),
    .B(net10001));
 sg13g2_o21ai_1 _18850_ (.B1(_11350_),
    .Y(_01637_),
    .A1(net9651),
    .A2(net10001));
 sg13g2_buf_2 place10719 (.A(net10718),
    .X(net10719));
 sg13g2_nand2_1 _18852_ (.Y(_11352_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][28] ),
    .B(net10001));
 sg13g2_o21ai_1 _18853_ (.B1(_11352_),
    .Y(_01638_),
    .A1(net9646),
    .A2(net10001));
 sg13g2_nand2_1 _18854_ (.Y(_11353_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][29] ),
    .B(net10000));
 sg13g2_o21ai_1 _18855_ (.B1(_11353_),
    .Y(_01639_),
    .A1(net9643),
    .A2(net10000));
 sg13g2_nand2_1 _18856_ (.Y(_11354_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][2] ),
    .B(net9996));
 sg13g2_o21ai_1 _18857_ (.B1(_11354_),
    .Y(_01640_),
    .A1(net10222),
    .A2(net9996));
 sg13g2_nand2_1 _18858_ (.Y(_11355_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][30] ),
    .B(net9999));
 sg13g2_o21ai_1 _18859_ (.B1(_11355_),
    .Y(_01641_),
    .A1(net9638),
    .A2(net9999));
 sg13g2_nand2_1 _18860_ (.Y(_11356_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][31] ),
    .B(net10000));
 sg13g2_o21ai_1 _18861_ (.B1(_11356_),
    .Y(_01642_),
    .A1(net9636),
    .A2(net10000));
 sg13g2_nand2_1 _18862_ (.Y(_11357_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][3] ),
    .B(net9997));
 sg13g2_o21ai_1 _18863_ (.B1(_11357_),
    .Y(_01643_),
    .A1(net10220),
    .A2(net9997));
 sg13g2_nand2_1 _18864_ (.Y(_11358_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][4] ),
    .B(net10003));
 sg13g2_o21ai_1 _18865_ (.B1(_11358_),
    .Y(_01644_),
    .A1(net10181),
    .A2(net10003));
 sg13g2_nand2_1 _18866_ (.Y(_11359_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][5] ),
    .B(net9996));
 sg13g2_o21ai_1 _18867_ (.B1(_11359_),
    .Y(_01645_),
    .A1(net10178),
    .A2(net9996));
 sg13g2_nand2_1 _18868_ (.Y(_11360_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][6] ),
    .B(net9995));
 sg13g2_o21ai_1 _18869_ (.B1(_11360_),
    .Y(_01646_),
    .A1(net10170),
    .A2(net9995));
 sg13g2_nand2_1 _18870_ (.Y(_11361_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][7] ),
    .B(net9995));
 sg13g2_o21ai_1 _18871_ (.B1(_11361_),
    .Y(_01647_),
    .A1(net10167),
    .A2(net9995));
 sg13g2_nand2_1 _18872_ (.Y(_11362_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][8] ),
    .B(net9998));
 sg13g2_o21ai_1 _18873_ (.B1(_11362_),
    .Y(_01648_),
    .A1(net10128),
    .A2(net9998));
 sg13g2_nand2_1 _18874_ (.Y(_11363_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][9] ),
    .B(net9995));
 sg13g2_o21ai_1 _18875_ (.B1(_11363_),
    .Y(_01649_),
    .A1(net9975),
    .A2(net9995));
 sg13g2_nand2_2 _18876_ (.Y(_11364_),
    .A(_09843_),
    .B(_10211_));
 sg13g2_buf_2 place10664 (.A(_00133_),
    .X(net10664));
 sg13g2_buf_2 place10445 (.A(net10444),
    .X(net10445));
 sg13g2_buf_2 place10744 (.A(net10741),
    .X(net10744));
 sg13g2_nand2_1 _18880_ (.Y(_11368_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][0] ),
    .B(net9826));
 sg13g2_o21ai_1 _18881_ (.B1(_11368_),
    .Y(_01650_),
    .A1(net10276),
    .A2(net9826));
 sg13g2_nand2_1 _18882_ (.Y(_11369_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][10] ),
    .B(net9829));
 sg13g2_o21ai_1 _18883_ (.B1(_11369_),
    .Y(_01651_),
    .A1(net10131),
    .A2(net9829));
 sg13g2_nand2_1 _18884_ (.Y(_11370_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][11] ),
    .B(net9832));
 sg13g2_o21ai_1 _18885_ (.B1(_11370_),
    .Y(_01652_),
    .A1(net9985),
    .A2(net9832));
 sg13g2_nand2_1 _18886_ (.Y(_11371_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][12] ),
    .B(net9827));
 sg13g2_o21ai_1 _18887_ (.B1(_11371_),
    .Y(_01653_),
    .A1(net9800),
    .A2(net9827));
 sg13g2_nand2_1 _18888_ (.Y(_11372_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][13] ),
    .B(net9826));
 sg13g2_o21ai_1 _18889_ (.B1(_11372_),
    .Y(_01654_),
    .A1(net9979),
    .A2(net9826));
 sg13g2_nand2_1 _18890_ (.Y(_11373_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][14] ),
    .B(_11364_));
 sg13g2_o21ai_1 _18891_ (.B1(_11373_),
    .Y(_01655_),
    .A1(net9795),
    .A2(_11364_));
 sg13g2_nand2_1 _18892_ (.Y(_11374_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][15] ),
    .B(net9829));
 sg13g2_o21ai_1 _18893_ (.B1(_11374_),
    .Y(_01656_),
    .A1(net9793),
    .A2(net9829));
 sg13g2_nand2_1 _18894_ (.Y(_11375_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][16] ),
    .B(net9829));
 sg13g2_o21ai_1 _18895_ (.B1(_11375_),
    .Y(_01657_),
    .A1(net9745),
    .A2(net9829));
 sg13g2_buf_2 place10450 (.A(_08297_),
    .X(net10450));
 sg13g2_nand2_1 _18897_ (.Y(_11377_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][17] ),
    .B(net9828));
 sg13g2_o21ai_1 _18898_ (.B1(_11377_),
    .Y(_01658_),
    .A1(net9740),
    .A2(net9828));
 sg13g2_nand2_1 _18899_ (.Y(_11378_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][18] ),
    .B(net9830));
 sg13g2_o21ai_1 _18900_ (.B1(_11378_),
    .Y(_01659_),
    .A1(net9738),
    .A2(net9830));
 sg13g2_buf_2 place10763 (.A(net10762),
    .X(net10763));
 sg13g2_nand2_1 _18902_ (.Y(_11380_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][19] ),
    .B(net9834));
 sg13g2_o21ai_1 _18903_ (.B1(_11380_),
    .Y(_01660_),
    .A1(net9724),
    .A2(net9834));
 sg13g2_nand2_1 _18904_ (.Y(_11381_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][1] ),
    .B(net9826));
 sg13g2_o21ai_1 _18905_ (.B1(_11381_),
    .Y(_01661_),
    .A1(net10227),
    .A2(net9826));
 sg13g2_nand2_1 _18906_ (.Y(_11382_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][20] ),
    .B(net9831));
 sg13g2_o21ai_1 _18907_ (.B1(_11382_),
    .Y(_01662_),
    .A1(net9718),
    .A2(net9831));
 sg13g2_nand2_1 _18908_ (.Y(_11383_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][21] ),
    .B(net9831));
 sg13g2_o21ai_1 _18909_ (.B1(_11383_),
    .Y(_01663_),
    .A1(net9714),
    .A2(net9831));
 sg13g2_nand2_1 _18910_ (.Y(_11384_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][22] ),
    .B(net9830));
 sg13g2_o21ai_1 _18911_ (.B1(_11384_),
    .Y(_01664_),
    .A1(net9696),
    .A2(net9830));
 sg13g2_nand2_1 _18912_ (.Y(_11385_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][23] ),
    .B(net9831));
 sg13g2_o21ai_1 _18913_ (.B1(_11385_),
    .Y(_01665_),
    .A1(net9691),
    .A2(net9831));
 sg13g2_nand2_1 _18914_ (.Y(_11386_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][24] ),
    .B(net9830));
 sg13g2_o21ai_1 _18915_ (.B1(_11386_),
    .Y(_01666_),
    .A1(net9686),
    .A2(net9830));
 sg13g2_nand2_1 _18916_ (.Y(_11387_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][25] ),
    .B(net9833));
 sg13g2_o21ai_1 _18917_ (.B1(_11387_),
    .Y(_01667_),
    .A1(net9678),
    .A2(net9833));
 sg13g2_buf_2 place10446 (.A(_08297_),
    .X(net10446));
 sg13g2_nand2_1 _18919_ (.Y(_11389_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][26] ),
    .B(net9834));
 sg13g2_o21ai_1 _18920_ (.B1(_11389_),
    .Y(_01668_),
    .A1(net9675),
    .A2(net9834));
 sg13g2_nand2_1 _18921_ (.Y(_11390_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][27] ),
    .B(net9834));
 sg13g2_o21ai_1 _18922_ (.B1(_11390_),
    .Y(_01669_),
    .A1(_10023_),
    .A2(net9834));
 sg13g2_buf_2 place10717 (.A(net10716),
    .X(net10717));
 sg13g2_nand2_1 _18924_ (.Y(_11392_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][28] ),
    .B(net9834));
 sg13g2_o21ai_1 _18925_ (.B1(_11392_),
    .Y(_01670_),
    .A1(net9646),
    .A2(net9834));
 sg13g2_nand2_1 _18926_ (.Y(_11393_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][29] ),
    .B(net9833));
 sg13g2_o21ai_1 _18927_ (.B1(_11393_),
    .Y(_01671_),
    .A1(net9643),
    .A2(net9833));
 sg13g2_nand2_1 _18928_ (.Y(_11394_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][2] ),
    .B(net9828));
 sg13g2_o21ai_1 _18929_ (.B1(_11394_),
    .Y(_01672_),
    .A1(net10222),
    .A2(net9828));
 sg13g2_nand2_1 _18930_ (.Y(_11395_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][30] ),
    .B(net9833));
 sg13g2_o21ai_1 _18931_ (.B1(_11395_),
    .Y(_01673_),
    .A1(net9638),
    .A2(net9833));
 sg13g2_nand2_1 _18932_ (.Y(_11396_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][31] ),
    .B(net9832));
 sg13g2_o21ai_1 _18933_ (.B1(_11396_),
    .Y(_01674_),
    .A1(net9636),
    .A2(net9832));
 sg13g2_nand2_1 _18934_ (.Y(_11397_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][3] ),
    .B(net9829));
 sg13g2_o21ai_1 _18935_ (.B1(_11397_),
    .Y(_01675_),
    .A1(net10220),
    .A2(net9829));
 sg13g2_nand2_1 _18936_ (.Y(_11398_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][4] ),
    .B(net9831));
 sg13g2_o21ai_1 _18937_ (.B1(_11398_),
    .Y(_01676_),
    .A1(net10182),
    .A2(net9831));
 sg13g2_nand2_1 _18938_ (.Y(_11399_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][5] ),
    .B(net9828));
 sg13g2_o21ai_1 _18939_ (.B1(_11399_),
    .Y(_01677_),
    .A1(net10174),
    .A2(net9828));
 sg13g2_nand2_1 _18940_ (.Y(_11400_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][6] ),
    .B(net9827));
 sg13g2_o21ai_1 _18941_ (.B1(_11400_),
    .Y(_01678_),
    .A1(net10170),
    .A2(net9827));
 sg13g2_nand2_1 _18942_ (.Y(_11401_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][7] ),
    .B(net9827));
 sg13g2_o21ai_1 _18943_ (.B1(_11401_),
    .Y(_01679_),
    .A1(net10167),
    .A2(net9827));
 sg13g2_nand2_1 _18944_ (.Y(_11402_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][8] ),
    .B(_11364_));
 sg13g2_o21ai_1 _18945_ (.B1(_11402_),
    .Y(_01680_),
    .A1(net10126),
    .A2(_11364_));
 sg13g2_nand2_1 _18946_ (.Y(_11403_),
    .A(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][9] ),
    .B(net9827));
 sg13g2_o21ai_1 _18947_ (.B1(_11403_),
    .Y(_01681_),
    .A1(net9975),
    .A2(net9827));
 sg13g2_inv_4 _18948_ (.A(\u_ac_controller_soc_inst.u_picorv32.is_alu_reg_imm ),
    .Y(_11404_));
 sg13g2_nand3b_1 _18949_ (.B(_00101_),
    .C(_11404_),
    .Y(_11405_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.instr_jalr ));
 sg13g2_buf_2 place10712 (.A(net10710),
    .X(net10712));
 sg13g2_nand2_2 _18951_ (.Y(_11407_),
    .A(_08861_),
    .B(_08341_));
 sg13g2_or2_1 _18952_ (.X(_11408_),
    .B(_11407_),
    .A(_11405_));
 sg13g2_buf_2 place10441 (.A(net10440),
    .X(net10441));
 sg13g2_inv_2 _18954_ (.Y(_11410_),
    .A(net10660));
 sg13g2_nor2_2 _18955_ (.A(net10380),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoder_pseudo_trigger ),
    .Y(_11411_));
 sg13g2_buf_2 place10711 (.A(net10710),
    .X(net10711));
 sg13g2_o21ai_1 _18957_ (.B1(_11411_),
    .Y(_11413_),
    .A1(_00045_),
    .A2(_11408_));
 sg13g2_buf_2 place10748 (.A(net10747),
    .X(net10748));
 sg13g2_buf_2 place10752 (.A(net10747),
    .X(net10752));
 sg13g2_a22oi_1 _18960_ (.Y(_11416_),
    .B1(_11405_),
    .B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.is_sb_sh_sw ));
 sg13g2_buf_2 place10440 (.A(_08310_),
    .X(net10440));
 sg13g2_nand2b_2 _18962_ (.Y(_11418_),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoder_trigger ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.decoder_pseudo_trigger ));
 sg13g2_buf_2 place10723 (.A(net10722),
    .X(net10723));
 sg13g2_buf_2 place10713 (.A(net10709),
    .X(net10713));
 sg13g2_buf_2 place10439 (.A(_08312_),
    .X(net10439));
 sg13g2_nand2_2 _18966_ (.Y(_11422_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[0] ),
    .B(net10369));
 sg13g2_o21ai_1 _18967_ (.B1(_11422_),
    .Y(_01682_),
    .A1(_11413_),
    .A2(_11416_));
 sg13g2_buf_2 place10739 (.A(net10738),
    .X(net10739));
 sg13g2_buf_2 place10444 (.A(_08306_),
    .X(net10444));
 sg13g2_buf_2 place10442 (.A(net10441),
    .X(net10442));
 sg13g2_buf_2 place10433 (.A(_08320_),
    .X(net10433));
 sg13g2_a22oi_1 _18972_ (.Y(_11427_),
    .B1(net10217),
    .B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[10] ),
    .A1(net10653));
 sg13g2_nand2_1 _18973_ (.Y(_11428_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[10] ),
    .B(net10369));
 sg13g2_o21ai_1 _18974_ (.B1(_11428_),
    .Y(_01683_),
    .A1(net10369),
    .A2(_11427_));
 sg13g2_buf_2 place10727 (.A(net10725),
    .X(net10727));
 sg13g2_a22oi_1 _18976_ (.Y(_11430_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11] ),
    .B2(net10654),
    .A2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.is_beq_bne_blt_bge_bltu_bgeu ));
 sg13g2_buf_2 place10432 (.A(net10431),
    .X(net10432));
 sg13g2_o21ai_1 _18978_ (.B1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[31] ),
    .Y(_11432_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.is_sb_sh_sw ),
    .A2(_11405_));
 sg13g2_a21oi_2 _18979_ (.B1(_11413_),
    .Y(_11433_),
    .A2(_11432_),
    .A1(_11430_));
 sg13g2_a21o_1 _18980_ (.A2(net10368),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[11] ),
    .B1(_11433_),
    .X(_01684_));
 sg13g2_buf_2 place10425 (.A(net10424),
    .X(net10425));
 sg13g2_buf_2 place10729 (.A(net10725),
    .X(net10729));
 sg13g2_and2_1 _18983_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[31] ),
    .B(net10217),
    .X(_11436_));
 sg13g2_buf_2 place10431 (.A(net10430),
    .X(net10431));
 sg13g2_a221oi_1 _18985_ (.B2(net10608),
    .C1(_11436_),
    .B1(_08306_),
    .A1(net10654),
    .Y(_11438_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12] ));
 sg13g2_nand2_1 _18986_ (.Y(_11439_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[12] ),
    .B(net10368));
 sg13g2_o21ai_1 _18987_ (.B1(_11439_),
    .Y(_01685_),
    .A1(net10163),
    .A2(_11438_));
 sg13g2_buf_2 place10420 (.A(_08345_),
    .X(net10420));
 sg13g2_a221oi_1 _18989_ (.B2(net10607),
    .C1(_11436_),
    .B1(_08306_),
    .A1(net10654),
    .Y(_11441_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[13] ));
 sg13g2_nand2_1 _18990_ (.Y(_11442_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[13] ),
    .B(net10368));
 sg13g2_o21ai_1 _18991_ (.B1(_11442_),
    .Y(_01686_),
    .A1(net10163),
    .A2(_11441_));
 sg13g2_a221oi_1 _18992_ (.B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[14] ),
    .C1(net10162),
    .B1(_08306_),
    .A1(net10654),
    .Y(_11443_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[14] ));
 sg13g2_nand2_1 _18993_ (.Y(_11444_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[14] ),
    .B(net10368));
 sg13g2_o21ai_1 _18994_ (.B1(_11444_),
    .Y(_01687_),
    .A1(net10163),
    .A2(_11443_));
 sg13g2_a221oi_1 _18995_ (.B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[15] ),
    .C1(net10162),
    .B1(_08306_),
    .A1(net10652),
    .Y(_11445_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15] ));
 sg13g2_nand2_1 _18996_ (.Y(_11446_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[15] ),
    .B(net10367));
 sg13g2_o21ai_1 _18997_ (.B1(_11446_),
    .Y(_01688_),
    .A1(net10163),
    .A2(_11445_));
 sg13g2_a221oi_1 _18998_ (.B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[16] ),
    .C1(net10162),
    .B1(_08306_),
    .A1(net10652),
    .Y(_11447_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[16] ));
 sg13g2_nand2_1 _18999_ (.Y(_11448_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[16] ),
    .B(net10367));
 sg13g2_o21ai_1 _19000_ (.B1(_11448_),
    .Y(_01689_),
    .A1(net10164),
    .A2(_11447_));
 sg13g2_a221oi_1 _19001_ (.B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[17] ),
    .C1(net10162),
    .B1(net10444),
    .A1(net10652),
    .Y(_11449_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17] ));
 sg13g2_nand2_1 _19002_ (.Y(_11450_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[17] ),
    .B(net10367));
 sg13g2_o21ai_1 _19003_ (.B1(_11450_),
    .Y(_01690_),
    .A1(net10164),
    .A2(_11449_));
 sg13g2_a221oi_1 _19004_ (.B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[18] ),
    .C1(net10162),
    .B1(_08306_),
    .A1(net10652),
    .Y(_11451_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18] ));
 sg13g2_buf_2 place10419 (.A(net10417),
    .X(net10419));
 sg13g2_nand2_1 _19006_ (.Y(_11453_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[18] ),
    .B(net10367));
 sg13g2_o21ai_1 _19007_ (.B1(_11453_),
    .Y(_01691_),
    .A1(net10164),
    .A2(_11451_));
 sg13g2_a221oi_1 _19008_ (.B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[19] ),
    .C1(net10162),
    .B1(net10444),
    .A1(net10657),
    .Y(_11454_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[19] ));
 sg13g2_nand2_1 _19009_ (.Y(_11455_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[19] ),
    .B(net10365));
 sg13g2_o21ai_1 _19010_ (.B1(_11455_),
    .Y(_01692_),
    .A1(net10165),
    .A2(_11454_));
 sg13g2_nand2_1 _19011_ (.Y(_11456_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[21] ),
    .B(_11405_));
 sg13g2_a22oi_1 _19012_ (.Y(_11457_),
    .B1(_11407_),
    .B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1] ),
    .A1(net10653));
 sg13g2_a21oi_1 _19013_ (.A1(_11456_),
    .A2(_11457_),
    .Y(_11458_),
    .B1(_11413_));
 sg13g2_a21o_1 _19014_ (.A2(net10369),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[1] ),
    .B1(_11458_),
    .X(_01693_));
 sg13g2_buf_2 place10422 (.A(net10421),
    .X(net10422));
 sg13g2_buf_2 place10409 (.A(net10408),
    .X(net10409));
 sg13g2_buf_2 place10404 (.A(net10403),
    .X(net10404));
 sg13g2_a21o_2 _19018_ (.A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20] ),
    .A1(net10657),
    .B1(net10162),
    .X(_11462_));
 sg13g2_buf_2 place10417 (.A(net10416),
    .X(net10417));
 sg13g2_buf_16 clkbuf_leaf_248_clk (.X(clknet_leaf_248_clk),
    .A(clknet_8_73_0_clk));
 sg13g2_a21oi_1 _19021_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[20] ),
    .A2(net10444),
    .Y(_11465_),
    .B1(net9993));
 sg13g2_nand2_1 _19022_ (.Y(_11466_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[20] ),
    .B(net10366));
 sg13g2_o21ai_1 _19023_ (.B1(_11466_),
    .Y(_01694_),
    .A1(net10164),
    .A2(_11465_));
 sg13g2_buf_2 place10714 (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[2] ),
    .X(net10714));
 sg13g2_a21oi_1 _19025_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[21] ),
    .A2(net10445),
    .Y(_11468_),
    .B1(net9993));
 sg13g2_nand2_1 _19026_ (.Y(_11469_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[21] ),
    .B(net10366));
 sg13g2_o21ai_1 _19027_ (.B1(_11469_),
    .Y(_01695_),
    .A1(net10163),
    .A2(_11468_));
 sg13g2_a21oi_1 _19028_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[22] ),
    .A2(net10445),
    .Y(_11470_),
    .B1(net9993));
 sg13g2_nand2_1 _19029_ (.Y(_11471_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[22] ),
    .B(net10366));
 sg13g2_o21ai_1 _19030_ (.B1(_11471_),
    .Y(_01696_),
    .A1(net10164),
    .A2(_11470_));
 sg13g2_a21oi_1 _19031_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[23] ),
    .A2(net10445),
    .Y(_11472_),
    .B1(net9993));
 sg13g2_nand2_1 _19032_ (.Y(_11473_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[23] ),
    .B(net10367));
 sg13g2_o21ai_1 _19033_ (.B1(_11473_),
    .Y(_01697_),
    .A1(net10163),
    .A2(_11472_));
 sg13g2_a21oi_1 _19034_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[24] ),
    .A2(net10445),
    .Y(_11474_),
    .B1(net9993));
 sg13g2_nand2_1 _19035_ (.Y(_11475_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[24] ),
    .B(net10367));
 sg13g2_o21ai_1 _19036_ (.B1(_11475_),
    .Y(_01698_),
    .A1(net10164),
    .A2(_11474_));
 sg13g2_buf_2 place10416 (.A(_08348_),
    .X(net10416));
 sg13g2_a21oi_1 _19038_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[25] ),
    .A2(net10445),
    .Y(_11477_),
    .B1(net9993));
 sg13g2_nand2_1 _19039_ (.Y(_11478_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[25] ),
    .B(net10366));
 sg13g2_o21ai_1 _19040_ (.B1(_11478_),
    .Y(_01699_),
    .A1(net10165),
    .A2(_11477_));
 sg13g2_buf_2 place10396 (.A(_08971_),
    .X(net10396));
 sg13g2_a21oi_1 _19042_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[26] ),
    .A2(net10445),
    .Y(_11480_),
    .B1(net9993));
 sg13g2_nand2_1 _19043_ (.Y(_11481_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[26] ),
    .B(net10366));
 sg13g2_o21ai_1 _19044_ (.B1(_11481_),
    .Y(_01700_),
    .A1(net10163),
    .A2(_11480_));
 sg13g2_buf_16 clkbuf_leaf_247_clk (.X(clknet_leaf_247_clk),
    .A(clknet_8_73_0_clk));
 sg13g2_a21oi_1 _19046_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27] ),
    .A2(net10444),
    .Y(_11483_),
    .B1(_11462_));
 sg13g2_nand2_1 _19047_ (.Y(_11484_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[27] ),
    .B(net10366));
 sg13g2_o21ai_1 _19048_ (.B1(_11484_),
    .Y(_01701_),
    .A1(net10165),
    .A2(_11483_));
 sg13g2_buf_16 clkbuf_leaf_246_clk (.X(clknet_leaf_246_clk),
    .A(clknet_8_67_0_clk));
 sg13g2_a21oi_1 _19050_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[28] ),
    .A2(net10445),
    .Y(_11486_),
    .B1(net9993));
 sg13g2_buf_16 clkbuf_leaf_245_clk (.X(clknet_leaf_245_clk),
    .A(clknet_8_67_0_clk));
 sg13g2_nand2_1 _19052_ (.Y(_11488_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[28] ),
    .B(net10366));
 sg13g2_o21ai_1 _19053_ (.B1(_11488_),
    .Y(_01702_),
    .A1(net10165),
    .A2(_11486_));
 sg13g2_buf_2 place10448 (.A(net10447),
    .X(net10448));
 sg13g2_a21oi_1 _19055_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[29] ),
    .A2(net10444),
    .Y(_11490_),
    .B1(_11462_));
 sg13g2_nand2_1 _19056_ (.Y(_11491_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[29] ),
    .B(net10365));
 sg13g2_o21ai_1 _19057_ (.B1(_11491_),
    .Y(_01703_),
    .A1(net10165),
    .A2(_11490_));
 sg13g2_and2_1 _19058_ (.A(net10655),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2] ),
    .X(_11492_));
 sg13g2_a221oi_1 _19059_ (.B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[9] ),
    .C1(_11492_),
    .B1(_11407_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[22] ),
    .Y(_11493_),
    .A2(_11405_));
 sg13g2_nand2_1 _19060_ (.Y(_11494_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[2] ),
    .B(net10370));
 sg13g2_o21ai_1 _19061_ (.B1(_11494_),
    .Y(_01704_),
    .A1(_11413_),
    .A2(_11493_));
 sg13g2_a21oi_1 _19062_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[30] ),
    .A2(net10444),
    .Y(_11495_),
    .B1(_11462_));
 sg13g2_nand2_1 _19063_ (.Y(_11496_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[30] ),
    .B(net10365));
 sg13g2_o21ai_1 _19064_ (.B1(_11496_),
    .Y(_01705_),
    .A1(net10165),
    .A2(_11495_));
 sg13g2_inv_4 _19065_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[31] ),
    .Y(_11497_));
 sg13g2_o21ai_1 _19066_ (.B1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[31] ),
    .Y(_11498_),
    .A1(net10444),
    .A2(net10217));
 sg13g2_buf_2 place10430 (.A(_08320_),
    .X(net10430));
 sg13g2_a21oi_1 _19068_ (.A1(net10657),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20] ),
    .Y(_11500_),
    .B1(net10365));
 sg13g2_a22oi_1 _19069_ (.Y(_01706_),
    .B1(_11498_),
    .B2(_11500_),
    .A2(net10365),
    .A1(_11497_));
 sg13g2_inv_2 _19070_ (.Y(_11501_),
    .A(net10657));
 sg13g2_buf_2 place10728 (.A(net10725),
    .X(net10728));
 sg13g2_nor2_1 _19072_ (.A(net10363),
    .B(_08548_),
    .Y(_11503_));
 sg13g2_a221oi_1 _19073_ (.B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[10] ),
    .C1(_11503_),
    .B1(_11407_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[23] ),
    .Y(_11504_),
    .A2(_11405_));
 sg13g2_nand2_1 _19074_ (.Y(_11505_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[3] ),
    .B(net10370));
 sg13g2_o21ai_1 _19075_ (.B1(_11505_),
    .Y(_01707_),
    .A1(_11413_),
    .A2(_11504_));
 sg13g2_nand2_1 _19076_ (.Y(_11506_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[24] ),
    .B(_11405_));
 sg13g2_a22oi_1 _19077_ (.Y(_11507_),
    .B1(_11407_),
    .B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[4] ),
    .A1(net10656));
 sg13g2_a21oi_1 _19078_ (.A1(_11506_),
    .A2(_11507_),
    .Y(_11508_),
    .B1(_11413_));
 sg13g2_a21o_1 _19079_ (.A2(net10371),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[4] ),
    .B1(_11508_),
    .X(_01708_));
 sg13g2_buf_2 place10454 (.A(net10453),
    .X(net10454));
 sg13g2_a22oi_1 _19081_ (.Y(_11510_),
    .B1(net10217),
    .B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[5] ),
    .A1(net10656));
 sg13g2_nand2_1 _19082_ (.Y(_11511_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[5] ),
    .B(net10371));
 sg13g2_o21ai_1 _19083_ (.B1(_11511_),
    .Y(_01709_),
    .A1(net10371),
    .A2(_11510_));
 sg13g2_buf_2 place10449 (.A(net10448),
    .X(net10449));
 sg13g2_a22oi_1 _19085_ (.Y(_11513_),
    .B1(net10217),
    .B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[6] ),
    .A1(net10656));
 sg13g2_nand2_1 _19086_ (.Y(_11514_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[6] ),
    .B(net10371));
 sg13g2_o21ai_1 _19087_ (.B1(_11514_),
    .Y(_01710_),
    .A1(net10371),
    .A2(_11513_));
 sg13g2_buf_2 place10423 (.A(net10422),
    .X(net10423));
 sg13g2_a22oi_1 _19089_ (.Y(_11516_),
    .B1(net10217),
    .B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[7] ),
    .A1(net10655));
 sg13g2_nand2_1 _19090_ (.Y(_11517_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[7] ),
    .B(net10370));
 sg13g2_o21ai_1 _19091_ (.B1(_11517_),
    .Y(_01711_),
    .A1(net10371),
    .A2(_11516_));
 sg13g2_buf_2 place10397 (.A(net10396),
    .X(net10397));
 sg13g2_a22oi_1 _19093_ (.Y(_11519_),
    .B1(net10217),
    .B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[28] ),
    .A2(net10663),
    .A1(net10655));
 sg13g2_nand2_1 _19094_ (.Y(_11520_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[8] ),
    .B(net10370));
 sg13g2_o21ai_1 _19095_ (.B1(_11520_),
    .Y(_01712_),
    .A1(net10370),
    .A2(_11519_));
 sg13g2_buf_2 place10418 (.A(net10417),
    .X(net10418));
 sg13g2_a22oi_1 _19097_ (.Y(_11522_),
    .B1(net10217),
    .B2(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[9] ),
    .A1(net10655));
 sg13g2_nand2_1 _19098_ (.Y(_11523_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[9] ),
    .B(net10370));
 sg13g2_o21ai_1 _19099_ (.B1(_11523_),
    .Y(_01713_),
    .A1(net10370),
    .A2(_11522_));
 sg13g2_buf_2 place10403 (.A(_08963_),
    .X(net10403));
 sg13g2_nor2_1 _19101_ (.A(net10607),
    .B(net10608),
    .Y(_11525_));
 sg13g2_nand2_2 _19102_ (.Y(_11526_),
    .A(_00121_),
    .B(_11525_));
 sg13g2_nand2_2 _19103_ (.Y(_11527_),
    .A(_08344_),
    .B(_11411_));
 sg13g2_buf_16 clkbuf_leaf_266_clk (.X(clknet_leaf_266_clk),
    .A(clknet_8_82_0_clk));
 sg13g2_nand2_1 _19105_ (.Y(_11529_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_lb ),
    .B(net10377));
 sg13g2_o21ai_1 _19106_ (.B1(_11529_),
    .Y(_01744_),
    .A1(_11526_),
    .A2(_11527_));
 sg13g2_inv_1 _19107_ (.Y(_11530_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_lbu ));
 sg13g2_buf_16 clkbuf_leaf_254_clk (.X(clknet_leaf_254_clk),
    .A(clknet_8_77_0_clk));
 sg13g2_nor3_2 _19109_ (.A(net10607),
    .B(net10608),
    .C(_00121_),
    .Y(_11532_));
 sg13g2_nand3_1 _19110_ (.B(net10274),
    .C(_11532_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_lb_lh_lw_lbu_lhu ),
    .Y(_11533_));
 sg13g2_o21ai_1 _19111_ (.B1(_11533_),
    .Y(_01745_),
    .A1(_11530_),
    .A2(net10274));
 sg13g2_inv_1 _19112_ (.Y(_11534_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_lh ));
 sg13g2_nor2b_2 _19113_ (.A(net10607),
    .B_N(net10608),
    .Y(_11535_));
 sg13g2_buf_2 place10424 (.A(net10421),
    .X(net10424));
 sg13g2_nor2b_2 _19115_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[14] ),
    .B_N(_11535_),
    .Y(_11537_));
 sg13g2_nand3_1 _19116_ (.B(net10274),
    .C(_11537_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_lb_lh_lw_lbu_lhu ),
    .Y(_11538_));
 sg13g2_o21ai_1 _19117_ (.B1(_11538_),
    .Y(_01746_),
    .A1(_11534_),
    .A2(net10274));
 sg13g2_nand2_2 _19118_ (.Y(_11539_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[14] ),
    .B(_11535_));
 sg13g2_nand2_1 _19119_ (.Y(_11540_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_lhu ),
    .B(net10377));
 sg13g2_o21ai_1 _19120_ (.B1(_11540_),
    .Y(_01747_),
    .A1(_11527_),
    .A2(_11539_));
 sg13g2_nand3b_1 _19121_ (.B(_00121_),
    .C(net10607),
    .Y(_11541_),
    .A_N(net10608));
 sg13g2_buf_2 place10410 (.A(net10406),
    .X(net10410));
 sg13g2_nand2_1 _19123_ (.Y(_11543_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_lw ),
    .B(net10377));
 sg13g2_o21ai_1 _19124_ (.B1(_11543_),
    .Y(_01749_),
    .A1(_11527_),
    .A2(_11541_));
 sg13g2_nand2b_2 _19125_ (.Y(_11544_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[13] ),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[12] ));
 sg13g2_nand2_2 _19126_ (.Y(_11545_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[0] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[1] ));
 sg13g2_nor3_2 _19127_ (.A(_11418_),
    .B(_11544_),
    .C(_11545_),
    .Y(_11546_));
 sg13g2_inv_1 _19128_ (.Y(_11547_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[31] ));
 sg13g2_nor4_1 _19129_ (.A(_11547_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[14] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[16] ),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[24] ),
    .Y(_11548_));
 sg13g2_nor4_1 _19130_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[17] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[18] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[19] ),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[22] ),
    .Y(_11549_));
 sg13g2_nand3_1 _19131_ (.B(_11548_),
    .C(_11549_),
    .A(_11546_),
    .Y(_11550_));
 sg13g2_inv_1 _19132_ (.Y(_11551_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[3] ));
 sg13g2_nand4_1 _19133_ (.B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[4] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[5] ),
    .A(_11551_),
    .Y(_11552_),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[6] ));
 sg13g2_or4_1 _19134_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[25] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[26] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[28] ),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[29] ),
    .X(_11553_));
 sg13g2_buf_2 place10405 (.A(net10404),
    .X(net10405));
 sg13g2_inv_1 _19136_ (.Y(_11555_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[30] ));
 sg13g2_or4_1 _19137_ (.A(_11555_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[23] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[15] ),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[2] ),
    .X(_11556_));
 sg13g2_nor4_2 _19138_ (.A(_11550_),
    .B(_11552_),
    .C(_11553_),
    .Y(_11557_),
    .D(_11556_));
 sg13g2_nand2b_2 _19139_ (.Y(_11558_),
    .B(_11557_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[21] ));
 sg13g2_nand2_1 _19140_ (.Y(_11559_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycle ),
    .B(net10365));
 sg13g2_o21ai_1 _19141_ (.B1(_11559_),
    .Y(_01752_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27] ),
    .A2(_11558_));
 sg13g2_inv_1 _19142_ (.Y(_11560_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27] ));
 sg13g2_nand2_1 _19143_ (.Y(_11561_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycleh ),
    .B(net10375));
 sg13g2_o21ai_1 _19144_ (.B1(_11561_),
    .Y(_01753_),
    .A1(_11560_),
    .A2(_11558_));
 sg13g2_nand3b_1 _19145_ (.B(_11557_),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[21] ),
    .Y(_11562_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[20] ));
 sg13g2_nand2_1 _19146_ (.Y(_11563_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstr ),
    .B(net10375));
 sg13g2_o21ai_1 _19147_ (.B1(_11563_),
    .Y(_01754_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27] ),
    .A2(_11562_));
 sg13g2_nand2_1 _19148_ (.Y(_11564_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh ),
    .B(net10375));
 sg13g2_o21ai_1 _19149_ (.B1(_11564_),
    .Y(_01755_),
    .A1(_11560_),
    .A2(_11562_));
 sg13g2_nand2_2 _19150_ (.Y(_11565_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_sb_sh_sw ),
    .B(net10274));
 sg13g2_nand2_1 _19151_ (.Y(_11566_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_sb ),
    .B(net10377));
 sg13g2_o21ai_1 _19152_ (.B1(_11566_),
    .Y(_01756_),
    .A1(_11526_),
    .A2(_11565_));
 sg13g2_nand2b_2 _19153_ (.Y(_11567_),
    .B(_11535_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[14] ));
 sg13g2_nand2_1 _19154_ (.Y(_11568_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_sh ),
    .B(net10377));
 sg13g2_o21ai_1 _19155_ (.B1(_11568_),
    .Y(_01757_),
    .A1(_11567_),
    .A2(_11565_));
 sg13g2_inv_1 _19156_ (.Y(_11569_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_slli ));
 sg13g2_nor4_2 _19157_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[30] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[31] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27] ),
    .Y(_11570_),
    .D(_11553_));
 sg13g2_nor2_2 _19158_ (.A(_11404_),
    .B(net10378),
    .Y(_11571_));
 sg13g2_nand3_1 _19159_ (.B(_11570_),
    .C(_11571_),
    .A(_11537_),
    .Y(_11572_));
 sg13g2_o21ai_1 _19160_ (.B1(_11572_),
    .Y(_01759_),
    .A1(_11569_),
    .A2(net10273));
 sg13g2_or4_1 _19161_ (.A(_11555_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[31] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27] ),
    .D(_11553_),
    .X(_11573_));
 sg13g2_nor2_2 _19162_ (.A(_11539_),
    .B(_11573_),
    .Y(_11574_));
 sg13g2_nor2_2 _19163_ (.A(_00122_),
    .B(net10378),
    .Y(_11575_));
 sg13g2_a22oi_1 _19164_ (.Y(_11576_),
    .B1(_11574_),
    .B2(_11575_),
    .A2(net10372),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_srai ));
 sg13g2_inv_1 _19165_ (.Y(_01765_),
    .A(_11576_));
 sg13g2_inv_2 _19166_ (.Y(_11577_),
    .A(_11575_));
 sg13g2_nor2_1 _19167_ (.A(_11539_),
    .B(_11577_),
    .Y(_11578_));
 sg13g2_a22oi_1 _19168_ (.Y(_11579_),
    .B1(_11570_),
    .B2(_11578_),
    .A2(net10373),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_srli ));
 sg13g2_inv_1 _19169_ (.Y(_01767_),
    .A(_11579_));
 sg13g2_nand2_1 _19170_ (.Y(_11580_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_sw ),
    .B(net10377));
 sg13g2_o21ai_1 _19171_ (.B1(_11580_),
    .Y(_01769_),
    .A1(_11541_),
    .A2(_11565_));
 sg13g2_inv_1 _19172_ (.Y(_11581_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_jalr_addi_slti_sltiu_xori_ori_andi ));
 sg13g2_nor2_1 _19173_ (.A(_11404_),
    .B(_11535_),
    .Y(_11582_));
 sg13g2_o21ai_1 _19174_ (.B1(_11411_),
    .Y(_11583_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_jalr ),
    .A2(_11582_));
 sg13g2_o21ai_1 _19175_ (.B1(_11583_),
    .Y(_01776_),
    .A1(_11581_),
    .A2(_11411_));
 sg13g2_a21oi_1 _19176_ (.A1(_11535_),
    .A2(_11570_),
    .Y(_11584_),
    .B1(_11574_));
 sg13g2_nand2_2 _19177_ (.Y(_11585_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_alu_reg_reg ),
    .B(net10274));
 sg13g2_nand2_1 _19178_ (.Y(_11586_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_sll_srl_sra ),
    .B(_11418_));
 sg13g2_o21ai_1 _19179_ (.B1(_11586_),
    .Y(_01779_),
    .A1(_11584_),
    .A2(_11585_));
 sg13g2_nor3_1 _19180_ (.A(_11404_),
    .B(_11418_),
    .C(_11584_),
    .Y(_11587_));
 sg13g2_a21o_1 _19181_ (.A2(_11418_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.is_slli_srli_srai ),
    .B1(_11587_),
    .X(_01780_));
 sg13g2_buf_2 place10414 (.A(_08348_),
    .X(net10414));
 sg13g2_buf_16 clkbuf_leaf_250_clk (.X(clknet_leaf_250_clk),
    .A(clknet_8_76_0_clk));
 sg13g2_buf_2 place10402 (.A(net10401),
    .X(net10402));
 sg13g2_a22oi_1 _19185_ (.Y(_11591_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[0] ),
    .B2(net10275),
    .A2(\u_ac_controller_soc_inst.u_picorv32.latched_rd[0] ),
    .A1(net10383));
 sg13g2_nand2_1 _19186_ (.Y(_11592_),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[0] ),
    .B(_08397_));
 sg13g2_o21ai_1 _19187_ (.B1(_11592_),
    .Y(_01784_),
    .A1(net10712),
    .A2(_11591_));
 sg13g2_a22oi_1 _19188_ (.Y(_11593_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[1] ),
    .B2(net10275),
    .A2(\u_ac_controller_soc_inst.u_picorv32.latched_rd[1] ),
    .A1(net10383));
 sg13g2_nand2_1 _19189_ (.Y(_11594_),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[1] ),
    .B(_08397_));
 sg13g2_o21ai_1 _19190_ (.B1(_11594_),
    .Y(_01785_),
    .A1(net10712),
    .A2(_11593_));
 sg13g2_a22oi_1 _19191_ (.Y(_11595_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[2] ),
    .B2(net10275),
    .A2(\u_ac_controller_soc_inst.u_picorv32.latched_rd[2] ),
    .A1(net10383));
 sg13g2_nand2_1 _19192_ (.Y(_11596_),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[2] ),
    .B(_08397_));
 sg13g2_o21ai_1 _19193_ (.B1(_11596_),
    .Y(_01786_),
    .A1(net10712),
    .A2(_11595_));
 sg13g2_a22oi_1 _19194_ (.Y(_11597_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[3] ),
    .B2(net10275),
    .A2(\u_ac_controller_soc_inst.u_picorv32.latched_rd[3] ),
    .A1(net10383));
 sg13g2_nand2_1 _19195_ (.Y(_11598_),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[3] ),
    .B(_08397_));
 sg13g2_o21ai_1 _19196_ (.B1(_11598_),
    .Y(_01787_),
    .A1(net10712),
    .A2(_11597_));
 sg13g2_a22oi_1 _19197_ (.Y(_11599_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[4] ),
    .B2(net10275),
    .A2(\u_ac_controller_soc_inst.u_picorv32.latched_rd[4] ),
    .A1(net10383));
 sg13g2_nand2_1 _19198_ (.Y(_11600_),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_rd[4] ),
    .B(_08397_));
 sg13g2_o21ai_1 _19199_ (.B1(_11600_),
    .Y(_01788_),
    .A1(net10712),
    .A2(_11599_));
 sg13g2_buf_16 clkbuf_leaf_265_clk (.X(clknet_leaf_265_clk),
    .A(clknet_8_82_0_clk));
 sg13g2_nor2_2 _19201_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_do_rinst ),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_do_prefetch ),
    .Y(_11602_));
 sg13g2_buf_16 clkbuf_leaf_262_clk (.X(clknet_leaf_262_clk),
    .A(clknet_8_82_0_clk));
 sg13g2_buf_16 clkbuf_leaf_256_clk (.X(clknet_leaf_256_clk),
    .A(clknet_8_79_0_clk));
 sg13g2_and2_1 _19204_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_store ),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_branch ),
    .X(_11605_));
 sg13g2_buf_16 clkbuf_leaf_255_clk (.X(clknet_leaf_255_clk),
    .A(clknet_8_77_0_clk));
 sg13g2_buf_16 clkbuf_leaf_261_clk (.X(clknet_leaf_261_clk),
    .A(clknet_8_82_0_clk));
 sg13g2_buf_16 clkbuf_leaf_258_clk (.X(clknet_leaf_258_clk),
    .A(clknet_8_88_0_clk));
 sg13g2_buf_16 clkbuf_leaf_257_clk (.X(clknet_leaf_257_clk),
    .A(clknet_8_88_0_clk));
 sg13g2_buf_2 place10407 (.A(net10406),
    .X(net10407));
 sg13g2_nand2_1 _19210_ (.Y(_11611_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[10] ),
    .B(net10350));
 sg13g2_nand2_2 _19211_ (.Y(_11612_),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_store ),
    .B(\u_ac_controller_soc_inst.u_picorv32.latched_branch ));
 sg13g2_buf_2 place10401 (.A(_08963_),
    .X(net10401));
 sg13g2_buf_2 place10863 (.A(net10862),
    .X(net10863));
 sg13g2_buf_2 place10395 (.A(_09117_),
    .X(net10395));
 sg13g2_nand2_1 _19215_ (.Y(_11616_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[10] ),
    .B(net10344));
 sg13g2_buf_2 place10747 (.A(spi_sensor_clk),
    .X(net10747));
 sg13g2_a21oi_1 _19217_ (.A1(_11611_),
    .A2(_11616_),
    .Y(_11618_),
    .B1(net10355));
 sg13g2_a21oi_2 _19218_ (.B1(_11618_),
    .Y(_11619_),
    .A2(net10355),
    .A1(net10594));
 sg13g2_nor3_2 _19219_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_do_rinst ),
    .B(net10610),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_do_prefetch ),
    .Y(_11620_));
 sg13g2_inv_1 _19220_ (.Y(_11621_),
    .A(_11620_));
 sg13g2_nand2b_2 _19221_ (.Y(_11622_),
    .B(net11048),
    .A_N(\u_ac_controller_soc_inst.trap ));
 sg13g2_nor3_2 _19222_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_state[1] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_state[0] ),
    .C(_11622_),
    .Y(_11623_));
 sg13g2_buf_2 place10400 (.A(_08969_),
    .X(net10400));
 sg13g2_o21ai_1 _19224_ (.B1(_11623_),
    .Y(_11625_),
    .A1(net10609),
    .A2(_11621_));
 sg13g2_buf_2 place10799 (.A(net10795),
    .X(net10799));
 sg13g2_buf_2 place10864 (.A(net10863),
    .X(net10864));
 sg13g2_buf_2 place10408 (.A(net10407),
    .X(net10408));
 sg13g2_buf_2 place10394 (.A(_09263_),
    .X(net10394));
 sg13g2_nand2_1 _19229_ (.Y(_11630_),
    .A(\u_ac_controller_soc_inst.cbus_addr[10] ),
    .B(net10215));
 sg13g2_o21ai_1 _19230_ (.B1(_11630_),
    .Y(_01791_),
    .A1(_11619_),
    .A2(net10215));
 sg13g2_buf_2 place10438 (.A(_08312_),
    .X(net10438));
 sg13g2_buf_2 place10443 (.A(_08310_),
    .X(net10443));
 sg13g2_nand2_1 _19233_ (.Y(_11633_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[11] ),
    .B(_11605_));
 sg13g2_nand2_1 _19234_ (.Y(_11634_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[11] ),
    .B(net10340));
 sg13g2_buf_2 place10385 (.A(_09828_),
    .X(net10385));
 sg13g2_a21oi_1 _19236_ (.A1(_11633_),
    .A2(_11634_),
    .Y(_11636_),
    .B1(_11602_));
 sg13g2_a21oi_2 _19237_ (.B1(_11636_),
    .Y(_11637_),
    .A2(net10355),
    .A1(net10592));
 sg13g2_nand2_1 _19238_ (.Y(_11638_),
    .A(\u_ac_controller_soc_inst.cbus_addr[11] ),
    .B(net10215));
 sg13g2_o21ai_1 _19239_ (.B1(_11638_),
    .Y(_01792_),
    .A1(net10215),
    .A2(_11637_));
 sg13g2_nand2_1 _19240_ (.Y(_11639_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[12] ),
    .B(net10350));
 sg13g2_buf_2 place10427 (.A(net10420),
    .X(net10427));
 sg13g2_nand2_1 _19242_ (.Y(_11641_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[12] ),
    .B(net10344));
 sg13g2_a21oi_1 _19243_ (.A1(_11639_),
    .A2(_11641_),
    .Y(_11642_),
    .B1(net10355));
 sg13g2_a21oi_2 _19244_ (.B1(_11642_),
    .Y(_11643_),
    .A2(net10355),
    .A1(net10589));
 sg13g2_nand2_1 _19245_ (.Y(_11644_),
    .A(\u_ac_controller_soc_inst.cbus_addr[12] ),
    .B(net10214));
 sg13g2_o21ai_1 _19246_ (.B1(_11644_),
    .Y(_01793_),
    .A1(net10214),
    .A2(_11643_));
 sg13g2_nand2_1 _19247_ (.Y(_11645_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[13] ),
    .B(_11605_));
 sg13g2_nand2_1 _19248_ (.Y(_11646_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[13] ),
    .B(net10340));
 sg13g2_a21oi_1 _19249_ (.A1(_11645_),
    .A2(_11646_),
    .Y(_11647_),
    .B1(_11602_));
 sg13g2_a21oi_2 _19250_ (.B1(_11647_),
    .Y(_11648_),
    .A2(_11602_),
    .A1(net10587));
 sg13g2_nand2_1 _19251_ (.Y(_11649_),
    .A(net10625),
    .B(net10215));
 sg13g2_o21ai_1 _19252_ (.B1(_11649_),
    .Y(_01794_),
    .A1(net10213),
    .A2(_11648_));
 sg13g2_nand2_1 _19253_ (.Y(_11650_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[14] ),
    .B(net10349));
 sg13g2_nand2_2 _19254_ (.Y(_11651_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[14] ),
    .B(net10340));
 sg13g2_a21oi_1 _19255_ (.A1(_11650_),
    .A2(_11651_),
    .Y(_11652_),
    .B1(net10354));
 sg13g2_a21oi_2 _19256_ (.B1(_11652_),
    .Y(_11653_),
    .A2(net10354),
    .A1(net10585));
 sg13g2_nand2_1 _19257_ (.Y(_11654_),
    .A(\u_ac_controller_soc_inst.cbus_addr[14] ),
    .B(net10216));
 sg13g2_o21ai_1 _19258_ (.B1(_11654_),
    .Y(_01795_),
    .A1(net10216),
    .A2(_11653_));
 sg13g2_nand2_1 _19259_ (.Y(_11655_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[15] ),
    .B(net10349));
 sg13g2_nand2_1 _19260_ (.Y(_11656_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[15] ),
    .B(net10340));
 sg13g2_a21oi_1 _19261_ (.A1(_11655_),
    .A2(_11656_),
    .Y(_11657_),
    .B1(net10354));
 sg13g2_a21oi_2 _19262_ (.B1(_11657_),
    .Y(_11658_),
    .A2(net10354),
    .A1(net10583));
 sg13g2_nand2_1 _19263_ (.Y(_11659_),
    .A(\u_ac_controller_soc_inst.cbus_addr[15] ),
    .B(net10216));
 sg13g2_o21ai_1 _19264_ (.B1(_11659_),
    .Y(_01796_),
    .A1(net10216),
    .A2(_11658_));
 sg13g2_nand2_1 _19265_ (.Y(_11660_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[16] ),
    .B(net10349));
 sg13g2_nand2_1 _19266_ (.Y(_11661_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[16] ),
    .B(net10341));
 sg13g2_a21oi_1 _19267_ (.A1(_11660_),
    .A2(_11661_),
    .Y(_11662_),
    .B1(net10354));
 sg13g2_a21oi_2 _19268_ (.B1(_11662_),
    .Y(_11663_),
    .A2(net10354),
    .A1(net10581));
 sg13g2_nand2_1 _19269_ (.Y(_11664_),
    .A(\u_ac_controller_soc_inst.cbus_addr[16] ),
    .B(net10216));
 sg13g2_o21ai_1 _19270_ (.B1(_11664_),
    .Y(_01797_),
    .A1(net10216),
    .A2(_11663_));
 sg13g2_nand2_1 _19271_ (.Y(_11665_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[17] ),
    .B(net10349));
 sg13g2_nand2_1 _19272_ (.Y(_11666_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[17] ),
    .B(net10341));
 sg13g2_a21oi_1 _19273_ (.A1(_11665_),
    .A2(_11666_),
    .Y(_11667_),
    .B1(net10354));
 sg13g2_a21oi_2 _19274_ (.B1(_11667_),
    .Y(_11668_),
    .A2(net10354),
    .A1(net10578));
 sg13g2_nand2_1 _19275_ (.Y(_11669_),
    .A(\u_ac_controller_soc_inst.cbus_addr[17] ),
    .B(net10214));
 sg13g2_o21ai_1 _19276_ (.B1(_11669_),
    .Y(_01798_),
    .A1(net10214),
    .A2(_11668_));
 sg13g2_nand2_1 _19277_ (.Y(_11670_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[18] ),
    .B(net10346));
 sg13g2_nand2_1 _19278_ (.Y(_11671_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[18] ),
    .B(net10341));
 sg13g2_a21oi_1 _19279_ (.A1(_11670_),
    .A2(_11671_),
    .Y(_11672_),
    .B1(net10358));
 sg13g2_a21oi_2 _19280_ (.B1(_11672_),
    .Y(_11673_),
    .A2(net10358),
    .A1(net10576));
 sg13g2_nand2_1 _19281_ (.Y(_11674_),
    .A(\u_ac_controller_soc_inst.cbus_addr[18] ),
    .B(net10212));
 sg13g2_o21ai_1 _19282_ (.B1(_11674_),
    .Y(_01799_),
    .A1(net10212),
    .A2(_11673_));
 sg13g2_nand2_1 _19283_ (.Y(_11675_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[19] ),
    .B(net10346));
 sg13g2_nand2_2 _19284_ (.Y(_11676_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[19] ),
    .B(net10341));
 sg13g2_a21oi_2 _19285_ (.B1(net10359),
    .Y(_11677_),
    .A2(_11676_),
    .A1(_11675_));
 sg13g2_a21oi_2 _19286_ (.B1(_11677_),
    .Y(_11678_),
    .A2(net10358),
    .A1(net10574));
 sg13g2_buf_2 place10801 (.A(net10799),
    .X(net10801));
 sg13g2_nand2_1 _19288_ (.Y(_11680_),
    .A(\u_ac_controller_soc_inst.cbus_addr[19] ),
    .B(net10213));
 sg13g2_o21ai_1 _19289_ (.B1(_11680_),
    .Y(_01800_),
    .A1(net10213),
    .A2(_11678_));
 sg13g2_buf_2 place10413 (.A(net10410),
    .X(net10413));
 sg13g2_nand2_1 _19291_ (.Y(_11682_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[20] ),
    .B(net10346));
 sg13g2_nand2_2 _19292_ (.Y(_11683_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[20] ),
    .B(net10342));
 sg13g2_a21oi_2 _19293_ (.B1(net10360),
    .Y(_11684_),
    .A2(_11683_),
    .A1(_11682_));
 sg13g2_a21oi_2 _19294_ (.B1(_11684_),
    .Y(_11685_),
    .A2(net10358),
    .A1(net10567));
 sg13g2_nand2_1 _19295_ (.Y(_11686_),
    .A(net10624),
    .B(_11625_));
 sg13g2_o21ai_1 _19296_ (.B1(_11686_),
    .Y(_01801_),
    .A1(_11625_),
    .A2(_11685_));
 sg13g2_buf_2 place10426 (.A(net10420),
    .X(net10426));
 sg13g2_buf_2 place10412 (.A(net10410),
    .X(net10412));
 sg13g2_nand2_1 _19299_ (.Y(_11689_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[21] ),
    .B(net10346));
 sg13g2_nand2_2 _19300_ (.Y(_11690_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[21] ),
    .B(net10342));
 sg13g2_buf_2 place10599 (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[0] ),
    .X(net10599));
 sg13g2_a21oi_2 _19302_ (.B1(net10360),
    .Y(_11692_),
    .A2(_11690_),
    .A1(_11689_));
 sg13g2_a21oi_2 _19303_ (.B1(_11692_),
    .Y(_11693_),
    .A2(net10358),
    .A1(net10565));
 sg13g2_nand2_1 _19304_ (.Y(_11694_),
    .A(net10623),
    .B(net10210));
 sg13g2_o21ai_1 _19305_ (.B1(_11694_),
    .Y(_01802_),
    .A1(net10210),
    .A2(_11693_));
 sg13g2_nand2_1 _19306_ (.Y(_11695_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[22] ),
    .B(net10347));
 sg13g2_nand2_2 _19307_ (.Y(_11696_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[22] ),
    .B(net10342));
 sg13g2_a21oi_2 _19308_ (.B1(net10361),
    .Y(_11697_),
    .A2(_11696_),
    .A1(_11695_));
 sg13g2_a21oi_2 _19309_ (.B1(_11697_),
    .Y(_11698_),
    .A2(net10358),
    .A1(net10561));
 sg13g2_nand2_1 _19310_ (.Y(_11699_),
    .A(\u_ac_controller_soc_inst.cbus_addr[22] ),
    .B(net10209));
 sg13g2_o21ai_1 _19311_ (.B1(_11699_),
    .Y(_01803_),
    .A1(net10209),
    .A2(_11698_));
 sg13g2_nand2_1 _19312_ (.Y(_11700_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[23] ),
    .B(net10347));
 sg13g2_nand2_2 _19313_ (.Y(_11701_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[23] ),
    .B(net10343));
 sg13g2_a21oi_2 _19314_ (.B1(net10361),
    .Y(_11702_),
    .A2(_11701_),
    .A1(_11700_));
 sg13g2_a21oi_2 _19315_ (.B1(_11702_),
    .Y(_11703_),
    .A2(net10358),
    .A1(net10559));
 sg13g2_nand2_1 _19316_ (.Y(_11704_),
    .A(net10622),
    .B(net10210));
 sg13g2_o21ai_1 _19317_ (.B1(_11704_),
    .Y(_01804_),
    .A1(net10210),
    .A2(_11703_));
 sg13g2_nand2_1 _19318_ (.Y(_11705_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[24] ),
    .B(net10347));
 sg13g2_nand2_2 _19319_ (.Y(_11706_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[24] ),
    .B(net10342));
 sg13g2_a21oi_2 _19320_ (.B1(net10361),
    .Y(_11707_),
    .A2(_11706_),
    .A1(_11705_));
 sg13g2_a21oi_2 _19321_ (.B1(_11707_),
    .Y(_11708_),
    .A2(_11602_),
    .A1(net10556));
 sg13g2_nand2_1 _19322_ (.Y(_11709_),
    .A(\u_ac_controller_soc_inst.cbus_addr[24] ),
    .B(net10208));
 sg13g2_o21ai_1 _19323_ (.B1(_11709_),
    .Y(_01805_),
    .A1(net10208),
    .A2(_11708_));
 sg13g2_nand2_1 _19324_ (.Y(_11710_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[25] ),
    .B(net10347));
 sg13g2_nand2_2 _19325_ (.Y(_11711_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[25] ),
    .B(net10343));
 sg13g2_a21oi_2 _19326_ (.B1(net10361),
    .Y(_11712_),
    .A2(_11711_),
    .A1(_11710_));
 sg13g2_a21oi_2 _19327_ (.B1(_11712_),
    .Y(_11713_),
    .A2(net10359),
    .A1(net10553));
 sg13g2_nand2_1 _19328_ (.Y(_11714_),
    .A(\u_ac_controller_soc_inst.cbus_addr[25] ),
    .B(net10208));
 sg13g2_o21ai_1 _19329_ (.B1(_11714_),
    .Y(_01806_),
    .A1(net10208),
    .A2(_11713_));
 sg13g2_nand2_1 _19330_ (.Y(_11715_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[26] ),
    .B(net10347));
 sg13g2_nand2_2 _19331_ (.Y(_11716_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[26] ),
    .B(net10343));
 sg13g2_a21oi_2 _19332_ (.B1(net10361),
    .Y(_11717_),
    .A2(_11716_),
    .A1(_11715_));
 sg13g2_a21oi_2 _19333_ (.B1(_11717_),
    .Y(_11718_),
    .A2(net10359),
    .A1(net10550));
 sg13g2_nand2_1 _19334_ (.Y(_11719_),
    .A(\u_ac_controller_soc_inst.cbus_addr[26] ),
    .B(net10208));
 sg13g2_o21ai_1 _19335_ (.B1(_11719_),
    .Y(_01807_),
    .A1(net10208),
    .A2(_11718_));
 sg13g2_nand2_1 _19336_ (.Y(_11720_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[27] ),
    .B(net10347));
 sg13g2_nand2_2 _19337_ (.Y(_11721_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[27] ),
    .B(net10343));
 sg13g2_a21oi_2 _19338_ (.B1(net10361),
    .Y(_11722_),
    .A2(_11721_),
    .A1(_11720_));
 sg13g2_a21oi_2 _19339_ (.B1(_11722_),
    .Y(_11723_),
    .A2(net10359),
    .A1(net10547));
 sg13g2_nand2_1 _19340_ (.Y(_11724_),
    .A(\u_ac_controller_soc_inst.cbus_addr[27] ),
    .B(net10208));
 sg13g2_o21ai_1 _19341_ (.B1(_11724_),
    .Y(_01808_),
    .A1(net10208),
    .A2(_11723_));
 sg13g2_nand2_1 _19342_ (.Y(_11725_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[28] ),
    .B(net10346));
 sg13g2_nand2_2 _19343_ (.Y(_11726_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[28] ),
    .B(net10343));
 sg13g2_a21oi_1 _19344_ (.A1(_11725_),
    .A2(_11726_),
    .Y(_11727_),
    .B1(net10360));
 sg13g2_a21oi_2 _19345_ (.B1(_11727_),
    .Y(_11728_),
    .A2(net10360),
    .A1(net10545));
 sg13g2_nand2_1 _19346_ (.Y(_11729_),
    .A(\u_ac_controller_soc_inst.cbus_addr[28] ),
    .B(net10209));
 sg13g2_o21ai_1 _19347_ (.B1(_11729_),
    .Y(_01809_),
    .A1(net10209),
    .A2(_11728_));
 sg13g2_nand2_1 _19348_ (.Y(_11730_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[29] ),
    .B(net10347));
 sg13g2_nand2_2 _19349_ (.Y(_11731_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[29] ),
    .B(net10342));
 sg13g2_a21oi_1 _19350_ (.A1(_11730_),
    .A2(_11731_),
    .Y(_11732_),
    .B1(net10360));
 sg13g2_a21oi_2 _19351_ (.B1(_11732_),
    .Y(_11733_),
    .A2(net10359),
    .A1(net10543));
 sg13g2_buf_2 place10737 (.A(net10735),
    .X(net10737));
 sg13g2_nand2_1 _19353_ (.Y(_11735_),
    .A(\u_ac_controller_soc_inst.cbus_addr[29] ),
    .B(net10207));
 sg13g2_o21ai_1 _19354_ (.B1(_11735_),
    .Y(_01810_),
    .A1(net10207),
    .A2(_11733_));
 sg13g2_buf_2 place10708 (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[4] ),
    .X(net10708));
 sg13g2_nand2_1 _19356_ (.Y(_11737_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[2] ),
    .B(net10352));
 sg13g2_buf_2 place10659 (.A(net10658),
    .X(net10659));
 sg13g2_nand2_1 _19358_ (.Y(_11739_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[2] ),
    .B(net10344));
 sg13g2_a21oi_1 _19359_ (.A1(_11737_),
    .A2(_11739_),
    .Y(_11740_),
    .B1(net10356));
 sg13g2_a21oi_1 _19360_ (.A1(net10540),
    .A2(net10357),
    .Y(_11741_),
    .B1(_11740_));
 sg13g2_buf_2 place10384 (.A(_09828_),
    .X(net10384));
 sg13g2_nand2_1 _19362_ (.Y(_11743_),
    .A(\u_ac_controller_soc_inst.cbus_addr[2] ),
    .B(net10213));
 sg13g2_o21ai_1 _19363_ (.B1(_11743_),
    .Y(_01811_),
    .A1(net10214),
    .A2(_11741_));
 sg13g2_nand2_1 _19364_ (.Y(_11744_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[30] ),
    .B(net10346));
 sg13g2_nand2_2 _19365_ (.Y(_11745_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[30] ),
    .B(net10343));
 sg13g2_a21oi_1 _19366_ (.A1(_11744_),
    .A2(_11745_),
    .Y(_11746_),
    .B1(net10360));
 sg13g2_a21oi_2 _19367_ (.B1(_11746_),
    .Y(_11747_),
    .A2(net10360),
    .A1(net10537));
 sg13g2_nand2_1 _19368_ (.Y(_11748_),
    .A(\u_ac_controller_soc_inst.cbus_addr[30] ),
    .B(net10209));
 sg13g2_o21ai_1 _19369_ (.B1(_11748_),
    .Y(_01812_),
    .A1(net10209),
    .A2(_11747_));
 sg13g2_nand2_1 _19370_ (.Y(_11749_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[31] ),
    .B(net10346));
 sg13g2_nand2_1 _19371_ (.Y(_11750_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[31] ),
    .B(net10341));
 sg13g2_a21oi_1 _19372_ (.A1(_11749_),
    .A2(_11750_),
    .Y(_11751_),
    .B1(net10359));
 sg13g2_a21oi_2 _19373_ (.B1(_11751_),
    .Y(_11752_),
    .A2(net10359),
    .A1(net10534));
 sg13g2_nand2_1 _19374_ (.Y(_11753_),
    .A(\u_ac_controller_soc_inst.cbus_addr[31] ),
    .B(net10209));
 sg13g2_o21ai_1 _19375_ (.B1(_11753_),
    .Y(_01813_),
    .A1(net10209),
    .A2(_11752_));
 sg13g2_nand2_1 _19376_ (.Y(_11754_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[3] ),
    .B(net10352));
 sg13g2_nand2_1 _19377_ (.Y(_11755_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[3] ),
    .B(net10344));
 sg13g2_a21oi_1 _19378_ (.A1(_11754_),
    .A2(_11755_),
    .Y(_11756_),
    .B1(net10356));
 sg13g2_a21oi_1 _19379_ (.A1(net10532),
    .A2(net10357),
    .Y(_11757_),
    .B1(_11756_));
 sg13g2_buf_2 place10382 (.A(_09847_),
    .X(net10382));
 sg13g2_nand2_1 _19381_ (.Y(_11759_),
    .A(\u_ac_controller_soc_inst.cbus_addr[3] ),
    .B(net10212));
 sg13g2_o21ai_1 _19382_ (.B1(_11759_),
    .Y(_01814_),
    .A1(net10212),
    .A2(_11757_));
 sg13g2_nand2_1 _19383_ (.Y(_11760_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[4] ),
    .B(net10352));
 sg13g2_nand2_1 _19384_ (.Y(_11761_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[4] ),
    .B(net10344));
 sg13g2_a21oi_1 _19385_ (.A1(_11760_),
    .A2(_11761_),
    .Y(_11762_),
    .B1(net10357));
 sg13g2_a21oi_1 _19386_ (.A1(net10530),
    .A2(net10357),
    .Y(_11763_),
    .B1(_11762_));
 sg13g2_nand2_1 _19387_ (.Y(_11764_),
    .A(\u_ac_controller_soc_inst.cbus_addr[4] ),
    .B(net10214));
 sg13g2_o21ai_1 _19388_ (.B1(_11764_),
    .Y(_01815_),
    .A1(net10214),
    .A2(_11763_));
 sg13g2_nand2_1 _19389_ (.Y(_11765_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[5] ),
    .B(net10352));
 sg13g2_nand2_1 _19390_ (.Y(_11766_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[5] ),
    .B(net10344));
 sg13g2_a21oi_1 _19391_ (.A1(_11765_),
    .A2(_11766_),
    .Y(_11767_),
    .B1(net10357));
 sg13g2_a21oi_2 _19392_ (.B1(_11767_),
    .Y(_11768_),
    .A2(net10357),
    .A1(net10529));
 sg13g2_nand2_1 _19393_ (.Y(_11769_),
    .A(net10615),
    .B(net10211));
 sg13g2_o21ai_1 _19394_ (.B1(_11769_),
    .Y(_01816_),
    .A1(net10211),
    .A2(_11768_));
 sg13g2_nand2_1 _19395_ (.Y(_11770_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[6] ),
    .B(net10352));
 sg13g2_nand2_1 _19396_ (.Y(_11771_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[6] ),
    .B(net10344));
 sg13g2_a21oi_1 _19397_ (.A1(_11770_),
    .A2(_11771_),
    .Y(_11772_),
    .B1(net10357));
 sg13g2_a21oi_2 _19398_ (.B1(_11772_),
    .Y(_11773_),
    .A2(net10357),
    .A1(net10527));
 sg13g2_nand2_1 _19399_ (.Y(_11774_),
    .A(net10614),
    .B(net10211));
 sg13g2_o21ai_1 _19400_ (.B1(_11774_),
    .Y(_01817_),
    .A1(net10211),
    .A2(_11773_));
 sg13g2_nand2_1 _19401_ (.Y(_11775_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[7] ),
    .B(net10352));
 sg13g2_nand2_1 _19402_ (.Y(_11776_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[7] ),
    .B(net10344));
 sg13g2_a21oi_1 _19403_ (.A1(_11775_),
    .A2(_11776_),
    .Y(_11777_),
    .B1(net10356));
 sg13g2_a21oi_2 _19404_ (.B1(_11777_),
    .Y(_11778_),
    .A2(net10356),
    .A1(net10525));
 sg13g2_nand2_1 _19405_ (.Y(_11779_),
    .A(net10613),
    .B(net10211));
 sg13g2_o21ai_1 _19406_ (.B1(_11779_),
    .Y(_01818_),
    .A1(net10210),
    .A2(_11778_));
 sg13g2_nand2_1 _19407_ (.Y(_11780_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[8] ),
    .B(net10350));
 sg13g2_nand2_1 _19408_ (.Y(_11781_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[8] ),
    .B(net10340));
 sg13g2_a21oi_1 _19409_ (.A1(_11780_),
    .A2(_11781_),
    .Y(_11782_),
    .B1(net10355));
 sg13g2_a21oi_2 _19410_ (.B1(_11782_),
    .Y(_11783_),
    .A2(net10355),
    .A1(net10523));
 sg13g2_nand2_1 _19411_ (.Y(_11784_),
    .A(\u_ac_controller_soc_inst.cbus_addr[8] ),
    .B(net10212));
 sg13g2_o21ai_1 _19412_ (.B1(_11784_),
    .Y(_01819_),
    .A1(net10212),
    .A2(_11783_));
 sg13g2_nand2_1 _19413_ (.Y(_11785_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_out[9] ),
    .B(net10352));
 sg13g2_nand2_1 _19414_ (.Y(_11786_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[9] ),
    .B(net10340));
 sg13g2_a21oi_1 _19415_ (.A1(_11785_),
    .A2(_11786_),
    .Y(_11787_),
    .B1(net10356));
 sg13g2_a21oi_2 _19416_ (.B1(_11787_),
    .Y(_11788_),
    .A2(net10356),
    .A1(net10522));
 sg13g2_nand2_1 _19417_ (.Y(_11789_),
    .A(net10611),
    .B(net10215));
 sg13g2_o21ai_1 _19418_ (.B1(_11789_),
    .Y(_01820_),
    .A1(net10215),
    .A2(_11788_));
 sg13g2_mux2_1 _19419_ (.A0(_00087_),
    .A1(net9810),
    .S(_07916_),
    .X(_11790_));
 sg13g2_nor2_1 _19420_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_state[1] ),
    .B(_07916_),
    .Y(_11791_));
 sg13g2_a221oi_1 _19421_ (.B2(net9810),
    .C1(\u_ac_controller_soc_inst.trap ),
    .B1(_11791_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_state[1] ),
    .Y(_11792_),
    .A2(_11790_));
 sg13g2_buf_2 place10389 (.A(net10387),
    .X(net10389));
 sg13g2_nand3_1 _19423_ (.B(_11623_),
    .C(_11620_),
    .A(_00112_),
    .Y(_11794_));
 sg13g2_o21ai_1 _19424_ (.B1(_11794_),
    .Y(_11795_),
    .A1(net11013),
    .A2(_11792_));
 sg13g2_buf_2 place10738 (.A(_00103_),
    .X(net10738));
 sg13g2_nand2_1 _19426_ (.Y(_11797_),
    .A(_00112_),
    .B(_11623_));
 sg13g2_nor4_1 _19427_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_state[1] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_do_rinst ),
    .C(net10610),
    .D(_11622_),
    .Y(_11798_));
 sg13g2_o21ai_1 _19428_ (.B1(\u_ac_controller_soc_inst.u_picorv32.mem_state[0] ),
    .Y(_11799_),
    .A1(_11795_),
    .A2(_11798_));
 sg13g2_o21ai_1 _19429_ (.B1(_11799_),
    .Y(_01825_),
    .A1(_11795_),
    .A2(_11797_));
 sg13g2_a221oi_1 _19430_ (.B2(\u_ac_controller_soc_inst.u_picorv32.mem_state[0] ),
    .C1(_11795_),
    .B1(_11798_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_do_wdata ),
    .Y(_11800_),
    .A2(_11623_));
 sg13g2_a21oi_1 _19431_ (.A1(_07914_),
    .A2(_11795_),
    .Y(_01826_),
    .B1(_11800_));
 sg13g2_and2_1 _19432_ (.A(net11048),
    .B(\u_ac_controller_soc_inst.trap ),
    .X(_11801_));
 sg13g2_and3_1 _19433_ (.X(_11802_),
    .A(_00112_),
    .B(_11623_),
    .C(_11620_));
 sg13g2_a21oi_1 _19434_ (.A1(_07935_),
    .A2(_11801_),
    .Y(_11803_),
    .B1(_11802_));
 sg13g2_a21oi_1 _19435_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_state[1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.mem_state[0] ),
    .Y(_11804_),
    .B1(net9810));
 sg13g2_o21ai_1 _19436_ (.B1(_11803_),
    .Y(_11805_),
    .A1(_11622_),
    .A2(_11804_));
 sg13g2_a22oi_1 _19437_ (.Y(_11806_),
    .B1(_11805_),
    .B2(\u_ac_controller_soc_inst.cbus_valid ),
    .A2(_11803_),
    .A1(_11623_));
 sg13g2_inv_1 _19438_ (.Y(_01827_),
    .A(_11806_));
 sg13g2_buf_2 place10406 (.A(_08363_),
    .X(net10406));
 sg13g2_and2_1 _19440_ (.A(net10609),
    .B(_11623_),
    .X(_11808_));
 sg13g2_buf_2 place10731 (.A(net10730),
    .X(net10731));
 sg13g2_buf_2 place10434 (.A(net10433),
    .X(net10434));
 sg13g2_buf_2 place10399 (.A(_08971_),
    .X(net10399));
 sg13g2_mux2_1 _19444_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[0] ),
    .A1(net10520),
    .S(net10198),
    .X(_01828_));
 sg13g2_buf_2 place10730 (.A(net10725),
    .X(net10730));
 sg13g2_and2_1 _19446_ (.A(net10604),
    .B(net10505),
    .X(_11813_));
 sg13g2_a21oi_2 _19447_ (.B1(_11813_),
    .Y(_11814_),
    .A2(net10394),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[10] ));
 sg13g2_buf_2 place10367 (.A(net10366),
    .X(net10367));
 sg13g2_buf_2 place10366 (.A(net10365),
    .X(net10366));
 sg13g2_nor2_1 _19450_ (.A(\u_ac_controller_soc_inst.cbus_wdata[10] ),
    .B(net10205),
    .Y(_11817_));
 sg13g2_a21oi_1 _19451_ (.A1(net10205),
    .A2(_11814_),
    .Y(_01829_),
    .B1(_11817_));
 sg13g2_buf_2 place10383 (.A(_09847_),
    .X(net10383));
 sg13g2_and2_1 _19453_ (.A(net10604),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[3] ),
    .X(_11819_));
 sg13g2_a21oi_2 _19454_ (.B1(_11819_),
    .Y(_11820_),
    .A2(net10394),
    .A1(net10519));
 sg13g2_buf_2 place10804 (.A(net10803),
    .X(net10804));
 sg13g2_nor2_1 _19456_ (.A(\u_ac_controller_soc_inst.cbus_wdata[11] ),
    .B(net10206),
    .Y(_11822_));
 sg13g2_a21oi_1 _19457_ (.A1(net10203),
    .A2(_11820_),
    .Y(_01830_),
    .B1(_11822_));
 sg13g2_and2_1 _19458_ (.A(net10604),
    .B(net10504),
    .X(_11823_));
 sg13g2_a21oi_2 _19459_ (.B1(_11823_),
    .Y(_11824_),
    .A2(net10394),
    .A1(net10518));
 sg13g2_buf_2 place10437 (.A(net10436),
    .X(net10437));
 sg13g2_nor2_1 _19461_ (.A(\u_ac_controller_soc_inst.cbus_wdata[12] ),
    .B(net10205),
    .Y(_11826_));
 sg13g2_a21oi_1 _19462_ (.A1(net10205),
    .A2(_11824_),
    .Y(_01831_),
    .B1(_11826_));
 sg13g2_and2_1 _19463_ (.A(net10604),
    .B(net10503),
    .X(_11827_));
 sg13g2_a21oi_1 _19464_ (.A1(net10517),
    .A2(net10394),
    .Y(_11828_),
    .B1(_11827_));
 sg13g2_buf_2 place10373 (.A(net10372),
    .X(net10373));
 sg13g2_nor2_1 _19466_ (.A(\u_ac_controller_soc_inst.cbus_wdata[13] ),
    .B(net10199),
    .Y(_11830_));
 sg13g2_a21oi_1 _19467_ (.A1(net10199),
    .A2(_11828_),
    .Y(_01832_),
    .B1(_11830_));
 sg13g2_and2_1 _19468_ (.A(net10604),
    .B(net10502),
    .X(_11831_));
 sg13g2_a21oi_2 _19469_ (.B1(_11831_),
    .Y(_11832_),
    .A2(net10394),
    .A1(net10516));
 sg13g2_buf_2 place10435 (.A(_08320_),
    .X(net10435));
 sg13g2_nor2_1 _19471_ (.A(\u_ac_controller_soc_inst.cbus_wdata[14] ),
    .B(net10202),
    .Y(_11834_));
 sg13g2_a21oi_1 _19472_ (.A1(net10203),
    .A2(_11832_),
    .Y(_01833_),
    .B1(_11834_));
 sg13g2_and2_1 _19473_ (.A(net10604),
    .B(net10501),
    .X(_11835_));
 sg13g2_a21oi_2 _19474_ (.B1(_11835_),
    .Y(_11836_),
    .A2(net10394),
    .A1(net10515));
 sg13g2_buf_16 clkbuf_leaf_268_clk (.X(clknet_leaf_268_clk),
    .A(clknet_8_80_0_clk));
 sg13g2_nor2_1 _19476_ (.A(\u_ac_controller_soc_inst.cbus_wdata[15] ),
    .B(net10202),
    .Y(_11838_));
 sg13g2_a21oi_1 _19477_ (.A1(net10202),
    .A2(_11836_),
    .Y(_01834_),
    .B1(_11838_));
 sg13g2_buf_16 clkbuf_leaf_267_clk (.X(clknet_leaf_267_clk),
    .A(clknet_8_77_0_clk));
 sg13g2_inv_8 _19479_ (.Y(_11840_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[16] ));
 sg13g2_nor2_1 _19480_ (.A(_11840_),
    .B(net10401),
    .Y(_11841_));
 sg13g2_a21oi_1 _19481_ (.A1(net10520),
    .A2(net10401),
    .Y(_11842_),
    .B1(_11841_));
 sg13g2_buf_2 place10371 (.A(net10370),
    .X(net10371));
 sg13g2_nor2_1 _19483_ (.A(\u_ac_controller_soc_inst.cbus_wdata[16] ),
    .B(net10203),
    .Y(_11844_));
 sg13g2_a21oi_1 _19484_ (.A1(net10203),
    .A2(_11842_),
    .Y(_01835_),
    .B1(_11844_));
 sg13g2_inv_8 _19485_ (.Y(_11845_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[17] ));
 sg13g2_nor2_1 _19486_ (.A(_11845_),
    .B(net10401),
    .Y(_11846_));
 sg13g2_a21oi_1 _19487_ (.A1(net10513),
    .A2(net10402),
    .Y(_11847_),
    .B1(_11846_));
 sg13g2_buf_2 place10362 (.A(_11501_),
    .X(net10362));
 sg13g2_nor2_1 _19489_ (.A(\u_ac_controller_soc_inst.cbus_wdata[17] ),
    .B(net10201),
    .Y(_11849_));
 sg13g2_a21oi_1 _19490_ (.A1(net10201),
    .A2(_11847_),
    .Y(_01836_),
    .B1(_11849_));
 sg13g2_nor2_1 _19491_ (.A(_08786_),
    .B(net10402),
    .Y(_11850_));
 sg13g2_a21oi_1 _19492_ (.A1(net10505),
    .A2(net10402),
    .Y(_11851_),
    .B1(_11850_));
 sg13g2_buf_2 place10451 (.A(_08292_),
    .X(net10451));
 sg13g2_buf_2 place10381 (.A(_09857_),
    .X(net10381));
 sg13g2_nor2_1 _19495_ (.A(\u_ac_controller_soc_inst.cbus_wdata[18] ),
    .B(net10201),
    .Y(_11854_));
 sg13g2_a21oi_1 _19496_ (.A1(net10201),
    .A2(_11851_),
    .Y(_01837_),
    .B1(_11854_));
 sg13g2_buf_2 place10392 (.A(_09819_),
    .X(net10392));
 sg13g2_nor2_1 _19498_ (.A(_08680_),
    .B(net10398),
    .Y(_11856_));
 sg13g2_a21oi_1 _19499_ (.A1(net10514),
    .A2(net10398),
    .Y(_11857_),
    .B1(_11856_));
 sg13g2_buf_2 place10369 (.A(net10368),
    .X(net10369));
 sg13g2_nor2_1 _19501_ (.A(\u_ac_controller_soc_inst.cbus_wdata[19] ),
    .B(net10206),
    .Y(_11859_));
 sg13g2_a21oi_1 _19502_ (.A1(net10206),
    .A2(_11857_),
    .Y(_01838_),
    .B1(_11859_));
 sg13g2_buf_2 place10363 (.A(net10362),
    .X(net10363));
 sg13g2_mux2_1 _19504_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[1] ),
    .A1(net10513),
    .S(net10198),
    .X(_01839_));
 sg13g2_buf_2 place10365 (.A(_11418_),
    .X(net10365));
 sg13g2_inv_8 _19506_ (.Y(_11862_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[20] ));
 sg13g2_nor2_1 _19507_ (.A(_11862_),
    .B(net10402),
    .Y(_11863_));
 sg13g2_a21oi_1 _19508_ (.A1(net10504),
    .A2(net10402),
    .Y(_11864_),
    .B1(_11863_));
 sg13g2_buf_2 place10370 (.A(net10369),
    .X(net10370));
 sg13g2_nor2_1 _19510_ (.A(\u_ac_controller_soc_inst.cbus_wdata[20] ),
    .B(net10206),
    .Y(_11866_));
 sg13g2_a21oi_1 _19511_ (.A1(net10206),
    .A2(_11864_),
    .Y(_01840_),
    .B1(_11866_));
 sg13g2_nor2_1 _19512_ (.A(_08801_),
    .B(net10401),
    .Y(_11867_));
 sg13g2_a21oi_1 _19513_ (.A1(net10503),
    .A2(net10402),
    .Y(_11868_),
    .B1(_11867_));
 sg13g2_buf_2 place10388 (.A(net10387),
    .X(net10388));
 sg13g2_nor2_1 _19515_ (.A(\u_ac_controller_soc_inst.cbus_wdata[21] ),
    .B(net10201),
    .Y(_11870_));
 sg13g2_a21oi_1 _19516_ (.A1(net10201),
    .A2(_11868_),
    .Y(_01841_),
    .B1(_11870_));
 sg13g2_and2_1 _19517_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[22] ),
    .B(net10398),
    .X(_11871_));
 sg13g2_a21oi_1 _19518_ (.A1(net10502),
    .A2(net10401),
    .Y(_11872_),
    .B1(_11871_));
 sg13g2_buf_2 place10368 (.A(net10367),
    .X(net10368));
 sg13g2_nor2_1 _19520_ (.A(\u_ac_controller_soc_inst.cbus_wdata[22] ),
    .B(net10200),
    .Y(_11874_));
 sg13g2_a21oi_1 _19521_ (.A1(net10200),
    .A2(_11872_),
    .Y(_01842_),
    .B1(_11874_));
 sg13g2_inv_8 _19522_ (.Y(_11875_),
    .A(net10511));
 sg13g2_nor2_1 _19523_ (.A(_11875_),
    .B(net10401),
    .Y(_11876_));
 sg13g2_a21oi_1 _19524_ (.A1(net10501),
    .A2(net10401),
    .Y(_11877_),
    .B1(_11876_));
 sg13g2_buf_2 place10386 (.A(net10385),
    .X(net10386));
 sg13g2_nor2_1 _19526_ (.A(\u_ac_controller_soc_inst.cbus_wdata[23] ),
    .B(net10199),
    .Y(_11879_));
 sg13g2_a21oi_1 _19527_ (.A1(_11808_),
    .A2(_11877_),
    .Y(_01843_),
    .B1(_11879_));
 sg13g2_and2_1 _19528_ (.A(net10604),
    .B(net10520),
    .X(_11880_));
 sg13g2_a221oi_1 _19529_ (.B2(net10398),
    .C1(_11880_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[24] ),
    .A1(net10602),
    .Y(_11881_),
    .A2(net10500));
 sg13g2_buf_2 place10358 (.A(_11602_),
    .X(net10358));
 sg13g2_nor2_1 _19531_ (.A(\u_ac_controller_soc_inst.cbus_wdata[24] ),
    .B(net10198),
    .Y(_11883_));
 sg13g2_a21oi_1 _19532_ (.A1(net10198),
    .A2(_11881_),
    .Y(_01844_),
    .B1(_11883_));
 sg13g2_and2_1 _19533_ (.A(net10604),
    .B(net10513),
    .X(_11884_));
 sg13g2_a221oi_1 _19534_ (.B2(net10398),
    .C1(_11884_),
    .B1(net10510),
    .A1(net10602),
    .Y(_11885_),
    .A2(net10499));
 sg13g2_buf_2 place10387 (.A(_09828_),
    .X(net10387));
 sg13g2_nor2_1 _19536_ (.A(\u_ac_controller_soc_inst.cbus_wdata[25] ),
    .B(_11808_),
    .Y(_11887_));
 sg13g2_a21oi_1 _19537_ (.A1(_11808_),
    .A2(_11885_),
    .Y(_01845_),
    .B1(_11887_));
 sg13g2_buf_2 place10364 (.A(_11501_),
    .X(net10364));
 sg13g2_a221oi_1 _19539_ (.B2(net10398),
    .C1(_11813_),
    .B1(net10509),
    .A1(net10602),
    .Y(_11889_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[10] ));
 sg13g2_buf_2 place10380 (.A(_11410_),
    .X(net10380));
 sg13g2_nor2_1 _19541_ (.A(\u_ac_controller_soc_inst.cbus_wdata[26] ),
    .B(net10201),
    .Y(_11891_));
 sg13g2_a21oi_1 _19542_ (.A1(net10200),
    .A2(_11889_),
    .Y(_01846_),
    .B1(_11891_));
 sg13g2_a221oi_1 _19543_ (.B2(net10398),
    .C1(_11819_),
    .B1(net10508),
    .A1(net10602),
    .Y(_11892_),
    .A2(net10519));
 sg13g2_buf_2 place10357 (.A(net10356),
    .X(net10357));
 sg13g2_nor2_1 _19545_ (.A(\u_ac_controller_soc_inst.cbus_wdata[27] ),
    .B(_11808_),
    .Y(_11894_));
 sg13g2_a21oi_1 _19546_ (.A1(_11808_),
    .A2(_11892_),
    .Y(_01847_),
    .B1(_11894_));
 sg13g2_a221oi_1 _19547_ (.B2(net10398),
    .C1(_11823_),
    .B1(net10507),
    .A1(net10602),
    .Y(_11895_),
    .A2(net10518));
 sg13g2_buf_2 place10372 (.A(_11418_),
    .X(net10372));
 sg13g2_nor2_1 _19549_ (.A(\u_ac_controller_soc_inst.cbus_wdata[28] ),
    .B(net10200),
    .Y(_11897_));
 sg13g2_a21oi_1 _19550_ (.A1(net10200),
    .A2(_11895_),
    .Y(_01848_),
    .B1(_11897_));
 sg13g2_a221oi_1 _19551_ (.B2(net10397),
    .C1(_11827_),
    .B1(net10506),
    .A1(net10602),
    .Y(_11898_),
    .A2(net10517));
 sg13g2_buf_2 place10334 (.A(net10333),
    .X(net10334));
 sg13g2_nor2_1 _19553_ (.A(\u_ac_controller_soc_inst.cbus_wdata[29] ),
    .B(net10198),
    .Y(_11900_));
 sg13g2_a21oi_1 _19554_ (.A1(net10198),
    .A2(_11898_),
    .Y(_01849_),
    .B1(_11900_));
 sg13g2_buf_2 place10345 (.A(_11605_),
    .X(net10345));
 sg13g2_mux2_1 _19556_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[2] ),
    .A1(net10505),
    .S(net10205),
    .X(_01850_));
 sg13g2_a221oi_1 _19557_ (.B2(net10397),
    .C1(_11831_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[30] ),
    .A1(net10602),
    .Y(_11902_),
    .A2(net10516));
 sg13g2_buf_2 place10348 (.A(net10345),
    .X(net10348));
 sg13g2_nor2_1 _19559_ (.A(\u_ac_controller_soc_inst.cbus_wdata[30] ),
    .B(net10200),
    .Y(_11904_));
 sg13g2_a21oi_1 _19560_ (.A1(net10200),
    .A2(_11902_),
    .Y(_01851_),
    .B1(_11904_));
 sg13g2_a221oi_1 _19561_ (.B2(net10397),
    .C1(_11835_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[31] ),
    .A1(net10602),
    .Y(_11905_),
    .A2(net10515));
 sg13g2_buf_2 place10343 (.A(net10342),
    .X(net10343));
 sg13g2_nor2_1 _19563_ (.A(\u_ac_controller_soc_inst.cbus_wdata[31] ),
    .B(net10199),
    .Y(_11907_));
 sg13g2_a21oi_1 _19564_ (.A1(net10199),
    .A2(_11905_),
    .Y(_01852_),
    .B1(_11907_));
 sg13g2_buf_2 place10350 (.A(_11605_),
    .X(net10350));
 sg13g2_mux2_1 _19566_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[3] ),
    .S(net10205),
    .X(_01853_));
 sg13g2_buf_2 place10356 (.A(net10355),
    .X(net10356));
 sg13g2_mux2_1 _19568_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[4] ),
    .A1(net10504),
    .S(net10205),
    .X(_01854_));
 sg13g2_buf_2 place10354 (.A(_11602_),
    .X(net10354));
 sg13g2_mux2_1 _19570_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[5] ),
    .A1(net10503),
    .S(net10204),
    .X(_01855_));
 sg13g2_buf_2 place10374 (.A(net10373),
    .X(net10374));
 sg13g2_mux2_1 _19572_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[6] ),
    .A1(net10502),
    .S(net10202),
    .X(_01856_));
 sg13g2_buf_2 place10359 (.A(_11602_),
    .X(net10359));
 sg13g2_mux2_1 _19574_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[7] ),
    .A1(net10501),
    .S(net10199),
    .X(_01857_));
 sg13g2_a21oi_2 _19575_ (.B1(_11880_),
    .Y(_11913_),
    .A2(net10394),
    .A1(net10500));
 sg13g2_buf_2 place10355 (.A(_11602_),
    .X(net10355));
 sg13g2_nor2_1 _19577_ (.A(\u_ac_controller_soc_inst.cbus_wdata[8] ),
    .B(net10204),
    .Y(_11915_));
 sg13g2_a21oi_1 _19578_ (.A1(net10204),
    .A2(_11913_),
    .Y(_01858_),
    .B1(_11915_));
 sg13g2_a21oi_2 _19579_ (.B1(_11884_),
    .Y(_11916_),
    .A2(net10394),
    .A1(net10499));
 sg13g2_buf_2 place10335 (.A(_11938_),
    .X(net10335));
 sg13g2_nor2_1 _19581_ (.A(\u_ac_controller_soc_inst.cbus_wdata[9] ),
    .B(net10205),
    .Y(_11918_));
 sg13g2_a21oi_1 _19582_ (.A1(net10204),
    .A2(_11916_),
    .Y(_01859_),
    .B1(_11918_));
 sg13g2_nand2_2 _19583_ (.Y(_11919_),
    .A(_11620_),
    .B(net10198));
 sg13g2_nor3_1 _19584_ (.A(net10571),
    .B(net10597),
    .C(net10603),
    .Y(_11920_));
 sg13g2_nor2_1 _19585_ (.A(_09265_),
    .B(_11920_),
    .Y(_11921_));
 sg13g2_nand2_1 _19586_ (.Y(_11922_),
    .A(\u_ac_controller_soc_inst.cbus_wstrb[0] ),
    .B(net10207));
 sg13g2_o21ai_1 _19587_ (.B1(_11922_),
    .Y(_01860_),
    .A1(_11919_),
    .A2(_11921_));
 sg13g2_nor2_1 _19588_ (.A(_09048_),
    .B(_09265_),
    .Y(_11923_));
 sg13g2_nand2_1 _19589_ (.Y(_11924_),
    .A(\u_ac_controller_soc_inst.cbus_wstrb[1] ),
    .B(net10207));
 sg13g2_o21ai_1 _19590_ (.B1(_11924_),
    .Y(_01861_),
    .A1(_11919_),
    .A2(_11923_));
 sg13g2_nand2b_1 _19591_ (.Y(_11925_),
    .B(net10596),
    .A_N(net10601));
 sg13g2_a21oi_1 _19592_ (.A1(net10571),
    .A2(_11925_),
    .Y(_11926_),
    .B1(net10397));
 sg13g2_buf_2 place10361 (.A(net10360),
    .X(net10361));
 sg13g2_nand2_1 _19594_ (.Y(_11928_),
    .A(\u_ac_controller_soc_inst.cbus_wstrb[2] ),
    .B(net10207));
 sg13g2_o21ai_1 _19595_ (.B1(_11928_),
    .Y(_01862_),
    .A1(_11919_),
    .A2(_11926_));
 sg13g2_buf_2 place10338 (.A(net10337),
    .X(net10338));
 sg13g2_o21ai_1 _19597_ (.B1(net10571),
    .Y(_11930_),
    .A1(net10601),
    .A2(net10596));
 sg13g2_a21oi_1 _19598_ (.A1(_08963_),
    .A2(_11930_),
    .Y(_11931_),
    .B1(_11919_));
 sg13g2_a21o_1 _19599_ (.A2(net10207),
    .A1(\u_ac_controller_soc_inst.cbus_wstrb[3] ),
    .B1(_11931_),
    .X(_01863_));
 sg13g2_and3_2 _19600_ (.X(_11932_),
    .A(_07697_),
    .B(_07940_),
    .C(_07969_));
 sg13g2_nand2_1 _19601_ (.Y(_11933_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_do_rdata ),
    .B(net10695));
 sg13g2_o21ai_1 _19602_ (.B1(_11933_),
    .Y(_11934_),
    .A1(_07953_),
    .A2(_00112_));
 sg13g2_a21oi_2 _19603_ (.B1(_11934_),
    .Y(_11935_),
    .A2(_07940_),
    .A1(_07697_));
 sg13g2_buf_2 place10375 (.A(net10372),
    .X(net10375));
 sg13g2_nor2_1 _19605_ (.A(_00109_),
    .B(_08365_),
    .Y(_11937_));
 sg13g2_nor2_2 _19606_ (.A(net10695),
    .B(\u_ac_controller_soc_inst.u_picorv32.cpu_state[5] ),
    .Y(_11938_));
 sg13g2_buf_2 place10337 (.A(net10335),
    .X(net10337));
 sg13g2_nand2_2 _19608_ (.Y(_11940_),
    .A(_09819_),
    .B(_11938_));
 sg13g2_o21ai_1 _19609_ (.B1(net11051),
    .Y(_11941_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpu_state[2] ),
    .A2(_11940_));
 sg13g2_a221oi_1 _19610_ (.B2(_08316_),
    .C1(_11941_),
    .B1(_11937_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpu_state[4] ),
    .Y(_11942_),
    .A2(_08365_));
 sg13g2_o21ai_1 _19611_ (.B1(_11942_),
    .Y(_11943_),
    .A1(_11932_),
    .A2(_11935_));
 sg13g2_buf_2 place10336 (.A(net10335),
    .X(net10336));
 sg13g2_buf_16 clkbuf_leaf_269_clk (.X(clknet_leaf_269_clk),
    .A(clknet_8_83_0_clk));
 sg13g2_buf_2 place10325 (.A(_12041_),
    .X(net10325));
 sg13g2_buf_2 place10317 (.A(_02186_),
    .X(net10317));
 sg13g2_or2_1 _19616_ (.X(_11948_),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_srai ),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_sra ));
 sg13g2_buf_2 place10324 (.A(net10323),
    .X(net10324));
 sg13g2_buf_2 place10360 (.A(net10359),
    .X(net10360));
 sg13g2_inv_2 _19619_ (.Y(_11951_),
    .A(_00055_));
 sg13g2_a22oi_1 _19620_ (.Y(_11952_),
    .B1(net10331),
    .B2(_11951_),
    .A2(net10442),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[4] ));
 sg13g2_buf_16 clkbuf_leaf_271_clk (.X(clknet_leaf_271_clk),
    .A(clknet_8_81_0_clk));
 sg13g2_buf_16 clkbuf_leaf_270_clk (.X(clknet_leaf_270_clk),
    .A(clknet_8_80_0_clk));
 sg13g2_inv_1 _19623_ (.Y(_11955_),
    .A(_00053_));
 sg13g2_a221oi_1 _19624_ (.B2(_11955_),
    .C1(net10413),
    .B1(net10331),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[1] ),
    .Y(_11956_),
    .A2(net10442));
 sg13g2_a21oi_1 _19625_ (.A1(net10413),
    .A2(_11952_),
    .Y(_11957_),
    .B1(_11956_));
 sg13g2_buf_2 place10318 (.A(net10317),
    .X(net10318));
 sg13g2_buf_2 place10323 (.A(net10321),
    .X(net10323));
 sg13g2_buf_2 place10311 (.A(_03816_),
    .X(net10311));
 sg13g2_buf_2 place10320 (.A(_02186_),
    .X(net10320));
 sg13g2_buf_2 place10310 (.A(_04546_),
    .X(net10310));
 sg13g2_buf_2 place10314 (.A(_03816_),
    .X(net10314));
 sg13g2_buf_2 place10322 (.A(net10321),
    .X(net10322));
 sg13g2_buf_2 place10313 (.A(net10311),
    .X(net10313));
 sg13g2_mux4_1 _19634_ (.S0(net10959),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][0] ),
    .S1(net10895),
    .X(_11966_));
 sg13g2_mux4_1 _19635_ (.S0(net10959),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][0] ),
    .S1(net10896),
    .X(_11967_));
 sg13g2_mux4_1 _19636_ (.S0(net10959),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][0] ),
    .S1(net10895),
    .X(_11968_));
 sg13g2_mux4_1 _19637_ (.S0(net10965),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][0] ),
    .S1(net10893),
    .X(_11969_));
 sg13g2_buf_2 place10312 (.A(net10311),
    .X(net10312));
 sg13g2_buf_2 place10306 (.A(_07148_),
    .X(net10306));
 sg13g2_buf_2 place10321 (.A(_12041_),
    .X(net10321));
 sg13g2_buf_2 place10305 (.A(_07148_),
    .X(net10305));
 sg13g2_buf_2 place10308 (.A(net10307),
    .X(net10308));
 sg13g2_mux4_1 _19643_ (.S0(net10885),
    .A0(_11966_),
    .A1(_11967_),
    .A2(_11968_),
    .A3(_11969_),
    .S1(_00008_),
    .X(_11975_));
 sg13g2_mux4_1 _19644_ (.S0(net10959),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][0] ),
    .S1(net10895),
    .X(_11976_));
 sg13g2_mux4_1 _19645_ (.S0(net10959),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][0] ),
    .S1(net10896),
    .X(_11977_));
 sg13g2_mux4_1 _19646_ (.S0(net10964),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][0] ),
    .S1(net10895),
    .X(_11978_));
 sg13g2_mux4_1 _19647_ (.S0(net10959),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][0] ),
    .S1(net10896),
    .X(_11979_));
 sg13g2_mux4_1 _19648_ (.S0(net10885),
    .A0(_11976_),
    .A1(_11977_),
    .A2(_11978_),
    .A3(_11979_),
    .S1(net10881),
    .X(_11980_));
 sg13g2_buf_16 clkbuf_leaf_275_clk (.X(clknet_leaf_275_clk),
    .A(clknet_8_71_0_clk));
 sg13g2_buf_16 clkbuf_leaf_273_clk (.X(clknet_leaf_273_clk),
    .A(clknet_8_80_0_clk));
 sg13g2_buf_16 clkbuf_leaf_272_clk (.X(clknet_leaf_272_clk),
    .A(clknet_8_80_0_clk));
 sg13g2_mux2_1 _19652_ (.A0(_11975_),
    .A1(_11980_),
    .S(net10872),
    .X(_11984_));
 sg13g2_buf_2 place10316 (.A(_03750_),
    .X(net10316));
 sg13g2_buf_2 place10300 (.A(_07720_),
    .X(net10300));
 sg13g2_nor4_1 _19655_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[16] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18] ),
    .D(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15] ),
    .Y(_11987_));
 sg13g2_a21oi_2 _19656_ (.B1(\u_ac_controller_soc_inst.u_picorv32.is_lui_auipc_jal ),
    .Y(_11988_),
    .A2(_11987_),
    .A1(_00132_));
 sg13g2_buf_2 place10319 (.A(_02186_),
    .X(net10319));
 sg13g2_buf_2 place10298 (.A(net10297),
    .X(net10298));
 sg13g2_buf_2 place10344 (.A(net10340),
    .X(net10344));
 sg13g2_nor2b_1 _19660_ (.A(net10272),
    .B_N(net10268),
    .Y(_11992_));
 sg13g2_inv_1 _19661_ (.Y(_11993_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[0] ));
 sg13g2_buf_2 place10303 (.A(_07193_),
    .X(net10303));
 sg13g2_nor3_1 _19663_ (.A(net10595),
    .B(_11993_),
    .C(net10334),
    .Y(_11995_));
 sg13g2_a221oi_1 _19664_ (.B2(_11992_),
    .C1(_11995_),
    .B1(_11984_),
    .A1(net10701),
    .Y(_11996_),
    .A2(_11957_));
 sg13g2_buf_2 place10309 (.A(_06692_),
    .X(net10309));
 sg13g2_buf_2 place10302 (.A(net10301),
    .X(net10302));
 sg13g2_buf_16 clkbuf_leaf_276_clk (.X(clknet_leaf_276_clk),
    .A(clknet_8_71_0_clk));
 sg13g2_nor2_1 _19668_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[0] ),
    .B(net10334),
    .Y(_12000_));
 sg13g2_o21ai_1 _19669_ (.B1(net10595),
    .Y(_12001_),
    .A1(net9672),
    .A2(_12000_));
 sg13g2_o21ai_1 _19670_ (.B1(_12001_),
    .Y(_01895_),
    .A1(net9672),
    .A2(_11996_));
 sg13g2_inv_2 _19671_ (.Y(_12002_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[10] ));
 sg13g2_a22oi_1 _19672_ (.Y(_12003_),
    .B1(net10528),
    .B2(net10671),
    .A2(net10526),
    .A1(net10670));
 sg13g2_nor2_1 _19673_ (.A(net10670),
    .B(net10526),
    .Y(_12004_));
 sg13g2_nor2_1 _19674_ (.A(_12003_),
    .B(_12004_),
    .Y(_12005_));
 sg13g2_a21oi_1 _19675_ (.A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[7] ),
    .A2(net10524),
    .Y(_12006_),
    .B1(_12005_));
 sg13g2_or2_1 _19676_ (.X(_12007_),
    .B(net10524),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[7] ));
 sg13g2_o21ai_1 _19677_ (.B1(_12007_),
    .Y(_12008_),
    .A1(net10669),
    .A2(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[8] ));
 sg13g2_nor2_1 _19678_ (.A(_12006_),
    .B(_12008_),
    .Y(_12009_));
 sg13g2_a21oi_2 _19679_ (.B1(_12009_),
    .Y(_12010_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[8] ),
    .A1(net10669));
 sg13g2_buf_2 place10301 (.A(net10300),
    .X(net10301));
 sg13g2_a21o_1 _19681_ (.A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[0] ),
    .A1(net10595),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[1] ),
    .X(_12012_));
 sg13g2_a21o_1 _19682_ (.A2(net10538),
    .A1(net10675),
    .B1(net10531),
    .X(_12013_));
 sg13g2_a21o_1 _19683_ (.A2(net10538),
    .A1(net10675),
    .B1(net10673),
    .X(_12014_));
 sg13g2_and3_1 _19684_ (.X(_12015_),
    .A(net10595),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[0] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[1] ));
 sg13g2_a221oi_1 _19685_ (.B2(_12014_),
    .C1(_12015_),
    .B1(_12013_),
    .A1(net10572),
    .Y(_12016_),
    .A2(_12012_));
 sg13g2_buf_2 place10295 (.A(_07774_),
    .X(net10295));
 sg13g2_nor2_1 _19687_ (.A(net10673),
    .B(net10531),
    .Y(_12018_));
 sg13g2_nor3_1 _19688_ (.A(net10675),
    .B(net10531),
    .C(net10539),
    .Y(_12019_));
 sg13g2_nor3_1 _19689_ (.A(net10675),
    .B(net10673),
    .C(net10539),
    .Y(_12020_));
 sg13g2_or3_1 _19690_ (.A(_12018_),
    .B(_12019_),
    .C(_12020_),
    .X(_12021_));
 sg13g2_buf_2 place10297 (.A(net10296),
    .X(net10297));
 sg13g2_o21ai_1 _19692_ (.B1(_08701_),
    .Y(_12023_),
    .A1(_12016_),
    .A2(_12021_));
 sg13g2_nor3_1 _19693_ (.A(_08701_),
    .B(_12016_),
    .C(_12021_),
    .Y(_12024_));
 sg13g2_a21oi_2 _19694_ (.B1(_12024_),
    .Y(_12025_),
    .A2(_12023_),
    .A1(net10672));
 sg13g2_xor2_1 _19695_ (.B(net10526),
    .A(net10670),
    .X(_12026_));
 sg13g2_o21ai_1 _19696_ (.B1(_12026_),
    .Y(_12027_),
    .A1(net10671),
    .A2(net10528));
 sg13g2_or3_1 _19697_ (.A(_12008_),
    .B(_12025_),
    .C(_12027_),
    .X(_12028_));
 sg13g2_buf_2 place10292 (.A(_07972_),
    .X(net10292));
 sg13g2_nand3_1 _19699_ (.B(_12010_),
    .C(_12028_),
    .A(_08709_),
    .Y(_12030_));
 sg13g2_a21oi_1 _19700_ (.A1(_12010_),
    .A2(_12028_),
    .Y(_12031_),
    .B1(_08709_));
 sg13g2_a21o_2 _19701_ (.A2(_12030_),
    .A1(net10668),
    .B1(_12031_),
    .X(_12032_));
 sg13g2_buf_2 place10293 (.A(net10292),
    .X(net10293));
 sg13g2_xnor2_1 _19703_ (.Y(_12034_),
    .A(net10694),
    .B(_12032_));
 sg13g2_a21oi_1 _19704_ (.A1(net10293),
    .A2(_12034_),
    .Y(_12035_),
    .B1(net9671));
 sg13g2_nor2_1 _19705_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[10] ),
    .B(_12034_),
    .Y(_12036_));
 sg13g2_buf_2 place10299 (.A(_07720_),
    .X(net10299));
 sg13g2_inv_2 _19707_ (.Y(_12038_),
    .A(_00060_));
 sg13g2_nor2_1 _19708_ (.A(_00063_),
    .B(net10412),
    .Y(_12039_));
 sg13g2_a21oi_1 _19709_ (.A1(_12038_),
    .A2(net10411),
    .Y(_12040_),
    .B1(_12039_));
 sg13g2_nor3_1 _19710_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_sh[2] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_sh[3] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.reg_sh[4] ),
    .Y(_12041_));
 sg13g2_buf_2 place10296 (.A(net10295),
    .X(net10296));
 sg13g2_buf_2 place10291 (.A(_08031_),
    .X(net10291));
 sg13g2_nand2_1 _19713_ (.Y(_02178_),
    .A(net10584),
    .B(net10440));
 sg13g2_o21ai_1 _19714_ (.B1(_02178_),
    .Y(_02179_),
    .A1(_00068_),
    .A2(net10438));
 sg13g2_buf_2 place10290 (.A(net10289),
    .X(net10290));
 sg13g2_inv_2 _19716_ (.Y(_02181_),
    .A(_00065_));
 sg13g2_a22oi_1 _19717_ (.Y(_02182_),
    .B1(net10331),
    .B2(_02181_),
    .A2(net10441),
    .A1(net10591));
 sg13g2_nand2_1 _19718_ (.Y(_02183_),
    .A(net10321),
    .B(_02182_));
 sg13g2_o21ai_1 _19719_ (.B1(_02183_),
    .Y(_02184_),
    .A1(net10322),
    .A2(_02179_));
 sg13g2_o21ai_1 _19720_ (.B1(_02184_),
    .Y(_02185_),
    .A1(net10290),
    .A2(_12040_));
 sg13g2_nor2b_2 _19721_ (.A(\u_ac_controller_soc_inst.u_picorv32.instr_lui ),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.is_lui_auipc_jal ),
    .Y(_02186_));
 sg13g2_buf_16 clkbuf_leaf_284_clk (.X(clknet_leaf_284_clk),
    .A(clknet_8_68_0_clk));
 sg13g2_buf_2 place10326 (.A(net10325),
    .X(net10326));
 sg13g2_buf_2 place10286 (.A(_08945_),
    .X(net10286));
 sg13g2_buf_16 clkbuf_leaf_281_clk (.X(clknet_leaf_281_clk),
    .A(clknet_8_69_0_clk));
 sg13g2_mux4_1 _19726_ (.S0(net10954),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][10] ),
    .S1(net10916),
    .X(_02191_));
 sg13g2_mux4_1 _19727_ (.S0(net10954),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][10] ),
    .S1(net10916),
    .X(_02192_));
 sg13g2_buf_16 clkbuf_leaf_279_clk (.X(clknet_leaf_279_clk),
    .A(clknet_8_69_0_clk));
 sg13g2_buf_16 clkbuf_leaf_278_clk (.X(clknet_leaf_278_clk),
    .A(clknet_8_69_0_clk));
 sg13g2_mux4_1 _19730_ (.S0(net10954),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][10] ),
    .S1(net10916),
    .X(_02195_));
 sg13g2_mux4_1 _19731_ (.S0(net10954),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][10] ),
    .S1(net10916),
    .X(_02196_));
 sg13g2_mux4_1 _19732_ (.S0(net10888),
    .A0(_02191_),
    .A1(_02192_),
    .A2(_02195_),
    .A3(_02196_),
    .S1(net10872),
    .X(_02197_));
 sg13g2_mux4_1 _19733_ (.S0(net10962),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][10] ),
    .S1(net10897),
    .X(_02198_));
 sg13g2_mux4_1 _19734_ (.S0(net10962),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][10] ),
    .S1(net10897),
    .X(_02199_));
 sg13g2_buf_16 clkbuf_leaf_285_clk (.X(clknet_leaf_285_clk),
    .A(clknet_8_80_0_clk));
 sg13g2_buf_2 place10294 (.A(_07972_),
    .X(net10294));
 sg13g2_mux4_1 _19737_ (.S0(net10961),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][10] ),
    .S1(net10898),
    .X(_02202_));
 sg13g2_mux4_1 _19738_ (.S0(net10961),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][10] ),
    .S1(net10898),
    .X(_02203_));
 sg13g2_mux4_1 _19739_ (.S0(net10889),
    .A0(_02198_),
    .A1(_02199_),
    .A2(_02202_),
    .A3(_02203_),
    .S1(net10873),
    .X(_02204_));
 sg13g2_buf_2 place10289 (.A(_08314_),
    .X(net10289));
 sg13g2_mux2_1 _19741_ (.A0(_02197_),
    .A1(_02204_),
    .S(net10882),
    .X(_02206_));
 sg13g2_a22oi_1 _19742_ (.Y(_02207_),
    .B1(_02206_),
    .B2(net10266),
    .A2(net10319),
    .A1(net10498));
 sg13g2_nor2_1 _19743_ (.A(net10271),
    .B(_02207_),
    .Y(_02208_));
 sg13g2_a221oi_1 _19744_ (.B2(net10704),
    .C1(_02208_),
    .B1(_02185_),
    .A1(net10292),
    .Y(_02209_),
    .A2(_12036_));
 sg13g2_or2_1 _19745_ (.X(_02210_),
    .B(_02209_),
    .A(net9671));
 sg13g2_o21ai_1 _19746_ (.B1(_02210_),
    .Y(_01896_),
    .A1(_12002_),
    .A2(_12035_));
 sg13g2_nand2_1 _19747_ (.Y(_02211_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[10] ),
    .B(_12032_));
 sg13g2_o21ai_1 _19748_ (.B1(net10694),
    .Y(_02212_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[10] ),
    .A2(_12032_));
 sg13g2_nand2_1 _19749_ (.Y(_02213_),
    .A(_02211_),
    .B(_02212_));
 sg13g2_xor2_1 _19750_ (.B(_02213_),
    .A(net10693),
    .X(_02214_));
 sg13g2_nor2_1 _19751_ (.A(net10591),
    .B(net10335),
    .Y(_02215_));
 sg13g2_buf_2 place10285 (.A(_08945_),
    .X(net10285));
 sg13g2_buf_2 place10284 (.A(net10283),
    .X(net10284));
 sg13g2_mux2_1 _19754_ (.A0(_00061_),
    .A1(_00064_),
    .S(net10322),
    .X(_02218_));
 sg13g2_buf_2 place10282 (.A(_08997_),
    .X(net10282));
 sg13g2_nand2_1 _19756_ (.Y(_02220_),
    .A(net10582),
    .B(net10440));
 sg13g2_o21ai_1 _19757_ (.B1(_02220_),
    .Y(_02221_),
    .A1(_00069_),
    .A2(net10438));
 sg13g2_buf_2 place10276 (.A(_09836_),
    .X(net10276));
 sg13g2_inv_2 _19759_ (.Y(_02223_),
    .A(_00066_));
 sg13g2_a22oi_1 _19760_ (.Y(_02224_),
    .B1(_11948_),
    .B2(_02223_),
    .A2(net10440),
    .A1(net10588));
 sg13g2_nand2_1 _19761_ (.Y(_02225_),
    .A(net10321),
    .B(_02224_));
 sg13g2_o21ai_1 _19762_ (.B1(_02225_),
    .Y(_02226_),
    .A1(net10321),
    .A2(_02221_));
 sg13g2_o21ai_1 _19763_ (.B1(_02226_),
    .Y(_02227_),
    .A1(net10290),
    .A2(_02218_));
 sg13g2_buf_16 clkbuf_leaf_288_clk (.X(clknet_leaf_288_clk),
    .A(clknet_8_85_0_clk));
 sg13g2_buf_2 place10288 (.A(net10287),
    .X(net10288));
 sg13g2_buf_2 place10287 (.A(net10286),
    .X(net10287));
 sg13g2_buf_2 place10315 (.A(net10314),
    .X(net10315));
 sg13g2_mux4_1 _19768_ (.S0(net10935),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][11] ),
    .S1(net10932),
    .X(_02232_));
 sg13g2_buf_2 place10281 (.A(_08997_),
    .X(net10281));
 sg13g2_buf_2 place10275 (.A(_09848_),
    .X(net10275));
 sg13g2_mux4_1 _19771_ (.S0(net10947),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][11] ),
    .S1(net10933),
    .X(_02235_));
 sg13g2_buf_2 place10273 (.A(_11411_),
    .X(net10273));
 sg13g2_buf_2 place10272 (.A(net10271),
    .X(net10272));
 sg13g2_buf_2 place10267 (.A(net10266),
    .X(net10267));
 sg13g2_buf_2 place10261 (.A(_03309_),
    .X(net10261));
 sg13g2_mux4_1 _19776_ (.S0(net10947),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][11] ),
    .S1(net10923),
    .X(_02240_));
 sg13g2_buf_16 clkbuf_leaf_293_clk (.X(clknet_leaf_293_clk),
    .A(clknet_8_94_0_clk));
 sg13g2_buf_2 place10274 (.A(_11411_),
    .X(net10274));
 sg13g2_mux4_1 _19779_ (.S0(net10949),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][11] ),
    .S1(net10933),
    .X(_02243_));
 sg13g2_buf_2 place10260 (.A(_03933_),
    .X(net10260));
 sg13g2_mux4_1 _19781_ (.S0(net10892),
    .A0(_02232_),
    .A1(_02235_),
    .A2(_02240_),
    .A3(_02243_),
    .S1(net10871),
    .X(_02245_));
 sg13g2_buf_16 clkbuf_leaf_292_clk (.X(clknet_leaf_292_clk),
    .A(clknet_8_87_0_clk));
 sg13g2_buf_16 clkbuf_leaf_289_clk (.X(clknet_leaf_289_clk),
    .A(clknet_8_87_0_clk));
 sg13g2_mux4_1 _19784_ (.S0(net10947),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][11] ),
    .S1(net10932),
    .X(_02248_));
 sg13g2_buf_2 place10283 (.A(net10282),
    .X(net10283));
 sg13g2_buf_16 clkbuf_leaf_299_clk (.X(clknet_leaf_299_clk),
    .A(clknet_8_87_0_clk));
 sg13g2_mux4_1 _19787_ (.S0(net10947),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][11] ),
    .S1(net10932),
    .X(_02251_));
 sg13g2_buf_16 clkbuf_leaf_295_clk (.X(clknet_leaf_295_clk),
    .A(clknet_8_86_0_clk));
 sg13g2_buf_2 place10259 (.A(_06402_),
    .X(net10259));
 sg13g2_buf_2 place10271 (.A(_11940_),
    .X(net10271));
 sg13g2_buf_2 place10270 (.A(net10269),
    .X(net10270));
 sg13g2_mux4_1 _19792_ (.S0(net10935),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][11] ),
    .S1(net10932),
    .X(_02256_));
 sg13g2_buf_2 place10277 (.A(net10276),
    .X(net10277));
 sg13g2_buf_16 clkbuf_leaf_315_clk (.X(clknet_leaf_315_clk),
    .A(clknet_8_92_0_clk));
 sg13g2_mux4_1 _19795_ (.S0(net10948),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][11] ),
    .S1(net10934),
    .X(_02259_));
 sg13g2_buf_16 clkbuf_leaf_304_clk (.X(clknet_leaf_304_clk),
    .A(clknet_8_84_0_clk));
 sg13g2_buf_2 place10279 (.A(net10276),
    .X(net10279));
 sg13g2_buf_2 place10351 (.A(net10350),
    .X(net10351));
 sg13g2_mux4_1 _19799_ (.S0(net10884),
    .A0(_02248_),
    .A1(_02251_),
    .A2(_02256_),
    .A3(_02259_),
    .S1(net10871),
    .X(_02263_));
 sg13g2_mux2_1 _19800_ (.A0(_02245_),
    .A1(_02263_),
    .S(net10879),
    .X(_02264_));
 sg13g2_a22oi_1 _19801_ (.Y(_02265_),
    .B1(_02264_),
    .B2(net10267),
    .A2(net10319),
    .A1(net10497));
 sg13g2_nor2_1 _19802_ (.A(net10271),
    .B(_02265_),
    .Y(_02266_));
 sg13g2_a221oi_1 _19803_ (.B2(net10703),
    .C1(_02266_),
    .B1(_02227_),
    .A1(_02214_),
    .Y(_02267_),
    .A2(_02215_));
 sg13g2_nor2_1 _19804_ (.A(net10335),
    .B(_02214_),
    .Y(_02268_));
 sg13g2_o21ai_1 _19805_ (.B1(net10591),
    .Y(_02269_),
    .A1(net9665),
    .A2(_02268_));
 sg13g2_o21ai_1 _19806_ (.B1(_02269_),
    .Y(_01897_),
    .A1(net9665),
    .A2(_02267_));
 sg13g2_nand3_1 _19807_ (.B(_02211_),
    .C(_02212_),
    .A(_08754_),
    .Y(_02270_));
 sg13g2_a21oi_1 _19808_ (.A1(_02211_),
    .A2(_02212_),
    .Y(_02271_),
    .B1(_08754_));
 sg13g2_a21o_2 _19809_ (.A2(_02270_),
    .A1(net10693),
    .B1(_02271_),
    .X(_02272_));
 sg13g2_buf_2 place10349 (.A(net10345),
    .X(net10349));
 sg13g2_xnor2_1 _19811_ (.Y(_02274_),
    .A(net10692),
    .B(_02272_));
 sg13g2_nor2_1 _19812_ (.A(net10588),
    .B(_02274_),
    .Y(_02275_));
 sg13g2_nor2_1 _19813_ (.A(_00062_),
    .B(net10322),
    .Y(_02276_));
 sg13g2_a21oi_1 _19814_ (.A1(_02181_),
    .A2(net10321),
    .Y(_02277_),
    .B1(_02276_));
 sg13g2_buf_16 clkbuf_leaf_301_clk (.X(clknet_leaf_301_clk),
    .A(clknet_8_85_0_clk));
 sg13g2_nand2_1 _19816_ (.Y(_02279_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[13] ),
    .B(net10440));
 sg13g2_o21ai_1 _19817_ (.B1(_02279_),
    .Y(_02280_),
    .A1(_00067_),
    .A2(net10438));
 sg13g2_buf_2 place10258 (.A(_06419_),
    .X(net10258));
 sg13g2_inv_1 _19819_ (.Y(_02282_),
    .A(_00070_));
 sg13g2_a22oi_1 _19820_ (.Y(_02283_),
    .B1(net10332),
    .B2(_02282_),
    .A2(net10440),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[16] ));
 sg13g2_nand2_1 _19821_ (.Y(_02284_),
    .A(net10406),
    .B(_02283_));
 sg13g2_o21ai_1 _19822_ (.B1(_02284_),
    .Y(_02285_),
    .A1(net10411),
    .A2(_02280_));
 sg13g2_o21ai_1 _19823_ (.B1(_02285_),
    .Y(_02286_),
    .A1(net10290),
    .A2(_02277_));
 sg13g2_mux4_1 _19824_ (.S0(net10971),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][12] ),
    .S1(net10907),
    .X(_02287_));
 sg13g2_mux4_1 _19825_ (.S0(net10971),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][12] ),
    .S1(net10906),
    .X(_02288_));
 sg13g2_mux4_1 _19826_ (.S0(net10971),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][12] ),
    .S1(net10907),
    .X(_02289_));
 sg13g2_mux4_1 _19827_ (.S0(net10974),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][12] ),
    .S1(net10910),
    .X(_02290_));
 sg13g2_buf_2 place10269 (.A(_11940_),
    .X(net10269));
 sg13g2_mux4_1 _19829_ (.S0(net10891),
    .A0(_02287_),
    .A1(_02288_),
    .A2(_02289_),
    .A3(_02290_),
    .S1(net10875),
    .X(_02292_));
 sg13g2_mux4_1 _19830_ (.S0(net10974),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][12] ),
    .S1(net10905),
    .X(_02293_));
 sg13g2_mux4_1 _19831_ (.S0(net10975),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][12] ),
    .S1(net10909),
    .X(_02294_));
 sg13g2_buf_2 place10265 (.A(_11988_),
    .X(net10265));
 sg13g2_buf_16 clkbuf_leaf_314_clk (.X(clknet_leaf_314_clk),
    .A(clknet_8_92_0_clk));
 sg13g2_mux4_1 _19834_ (.S0(net10973),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][12] ),
    .S1(net10910),
    .X(_02297_));
 sg13g2_mux4_1 _19835_ (.S0(net10973),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][12] ),
    .S1(net10910),
    .X(_02298_));
 sg13g2_mux4_1 _19836_ (.S0(net10891),
    .A0(_02293_),
    .A1(_02294_),
    .A2(_02297_),
    .A3(_02298_),
    .S1(net10874),
    .X(_02299_));
 sg13g2_mux2_1 _19837_ (.A0(_02292_),
    .A1(_02299_),
    .S(net10881),
    .X(_02300_));
 sg13g2_a22oi_1 _19838_ (.Y(_02301_),
    .B1(_02300_),
    .B2(net10266),
    .A2(net10319),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[12] ));
 sg13g2_nor2_1 _19839_ (.A(net10271),
    .B(_02301_),
    .Y(_02302_));
 sg13g2_a221oi_1 _19840_ (.B2(net10704),
    .C1(_02302_),
    .B1(_02286_),
    .A1(net10292),
    .Y(_02303_),
    .A2(_02275_));
 sg13g2_a21oi_1 _19841_ (.A1(net10292),
    .A2(_02274_),
    .Y(_02304_),
    .B1(net9671));
 sg13g2_nand2b_1 _19842_ (.Y(_02305_),
    .B(net10588),
    .A_N(_02304_));
 sg13g2_o21ai_1 _19843_ (.B1(_02305_),
    .Y(_01898_),
    .A1(net9671),
    .A2(_02303_));
 sg13g2_inv_2 _19844_ (.Y(_02306_),
    .A(net10691));
 sg13g2_or4_1 _19845_ (.A(_02306_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[13] ),
    .C(net10333),
    .D(_11943_),
    .X(_02307_));
 sg13g2_nand3_1 _19846_ (.B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[13] ),
    .C(net10292),
    .A(_02306_),
    .Y(_02308_));
 sg13g2_a21oi_1 _19847_ (.A1(net10693),
    .A2(_02270_),
    .Y(_02309_),
    .B1(_02271_));
 sg13g2_a21oi_1 _19848_ (.A1(net10588),
    .A2(_02272_),
    .Y(_02310_),
    .B1(net10692));
 sg13g2_a21oi_1 _19849_ (.A1(_08758_),
    .A2(_02309_),
    .Y(_02311_),
    .B1(_02310_));
 sg13g2_a21oi_1 _19850_ (.A1(_02307_),
    .A2(_02308_),
    .Y(_02312_),
    .B1(_02311_));
 sg13g2_nor2_2 _19851_ (.A(net10691),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[13] ),
    .Y(_02313_));
 sg13g2_nand3b_1 _19852_ (.B(_02313_),
    .C(net10292),
    .Y(_02314_),
    .A_N(_11943_));
 sg13g2_nor2_1 _19853_ (.A(_02306_),
    .B(_08761_),
    .Y(_02315_));
 sg13g2_nand2_1 _19854_ (.Y(_02316_),
    .A(net10292),
    .B(_02315_));
 sg13g2_a221oi_1 _19855_ (.B2(_02316_),
    .C1(_02310_),
    .B1(_02314_),
    .A1(_08758_),
    .Y(_02317_),
    .A2(_02309_));
 sg13g2_buf_16 clkbuf_leaf_313_clk (.X(clknet_leaf_313_clk),
    .A(clknet_8_92_0_clk));
 sg13g2_buf_16 clkbuf_leaf_311_clk (.X(clknet_leaf_311_clk),
    .A(clknet_8_86_0_clk));
 sg13g2_mux4_1 _19858_ (.S0(net10966),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][13] ),
    .S1(net10893),
    .X(_02320_));
 sg13g2_mux4_1 _19859_ (.S0(net10966),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][13] ),
    .S1(net10893),
    .X(_02321_));
 sg13g2_mux4_1 _19860_ (.S0(net10965),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][13] ),
    .S1(net10893),
    .X(_02322_));
 sg13g2_mux4_1 _19861_ (.S0(net10965),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][13] ),
    .S1(net10900),
    .X(_02323_));
 sg13g2_buf_16 clkbuf_leaf_308_clk (.X(clknet_leaf_308_clk),
    .A(clknet_8_83_0_clk));
 sg13g2_mux4_1 _19863_ (.S0(net10890),
    .A0(_02320_),
    .A1(_02321_),
    .A2(_02322_),
    .A3(_02323_),
    .S1(net10874),
    .X(_02325_));
 sg13g2_mux4_1 _19864_ (.S0(net10966),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][13] ),
    .S1(net10904),
    .X(_02326_));
 sg13g2_mux4_1 _19865_ (.S0(net10966),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][13] ),
    .S1(net10904),
    .X(_02327_));
 sg13g2_mux4_1 _19866_ (.S0(net10966),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][13] ),
    .S1(net10904),
    .X(_02328_));
 sg13g2_mux4_1 _19867_ (.S0(net10964),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][13] ),
    .S1(net10895),
    .X(_02329_));
 sg13g2_mux4_1 _19868_ (.S0(net10890),
    .A0(_02326_),
    .A1(_02327_),
    .A2(_02328_),
    .A3(_02329_),
    .S1(net10874),
    .X(_02330_));
 sg13g2_mux2_1 _19869_ (.A0(_02325_),
    .A1(_02330_),
    .S(net10881),
    .X(_02331_));
 sg13g2_a22oi_1 _19870_ (.Y(_02332_),
    .B1(_02331_),
    .B2(net10267),
    .A2(net10319),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[13] ));
 sg13g2_inv_2 _19871_ (.Y(_02333_),
    .A(_00063_));
 sg13g2_nand2_1 _19872_ (.Y(_02334_),
    .A(_02333_),
    .B(net10411));
 sg13g2_o21ai_1 _19873_ (.B1(_02334_),
    .Y(_02335_),
    .A1(_00066_),
    .A2(net10411));
 sg13g2_nor2_2 _19874_ (.A(net10441),
    .B(_11948_),
    .Y(_02336_));
 sg13g2_inv_1 _19875_ (.Y(_02337_),
    .A(_00071_));
 sg13g2_a22oi_1 _19876_ (.Y(_02338_),
    .B1(net10332),
    .B2(_02337_),
    .A2(net10440),
    .A1(net10577));
 sg13g2_nor2_1 _19877_ (.A(net10325),
    .B(_02338_),
    .Y(_02339_));
 sg13g2_a221oi_1 _19878_ (.B2(_02336_),
    .C1(_02339_),
    .B1(_02335_),
    .A1(net10321),
    .Y(_02340_),
    .A2(_02179_));
 sg13g2_nand2b_1 _19879_ (.Y(_02341_),
    .B(net10704),
    .A_N(_02340_));
 sg13g2_o21ai_1 _19880_ (.B1(_02341_),
    .Y(_02342_),
    .A1(net10271),
    .A2(_02332_));
 sg13g2_mux2_1 _19881_ (.A0(_02342_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[13] ),
    .S(_11943_),
    .X(_02343_));
 sg13g2_or3_1 _19882_ (.A(_02312_),
    .B(_02317_),
    .C(_02343_),
    .X(_01899_));
 sg13g2_inv_2 _19883_ (.Y(_02344_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[14] ));
 sg13g2_or4_1 _19884_ (.A(_02344_),
    .B(net10584),
    .C(_11938_),
    .D(_11943_),
    .X(_02345_));
 sg13g2_buf_16 clkbuf_leaf_306_clk (.X(clknet_leaf_306_clk),
    .A(clknet_8_81_0_clk));
 sg13g2_nand3_1 _19886_ (.B(net10584),
    .C(net10292),
    .A(_02344_),
    .Y(_02347_));
 sg13g2_a221oi_1 _19887_ (.B2(net10692),
    .C1(_02272_),
    .B1(net10588),
    .A1(net10691),
    .Y(_02348_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[13] ));
 sg13g2_nor3_1 _19888_ (.A(net10692),
    .B(net10588),
    .C(_02315_),
    .Y(_02349_));
 sg13g2_nor3_1 _19889_ (.A(_02313_),
    .B(_02348_),
    .C(_02349_),
    .Y(_02350_));
 sg13g2_a21oi_1 _19890_ (.A1(_02345_),
    .A2(_02347_),
    .Y(_02351_),
    .B1(_02350_));
 sg13g2_buf_2 place10266 (.A(_11988_),
    .X(net10266));
 sg13g2_nor4_1 _19892_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[14] ),
    .B(net10584),
    .C(_11938_),
    .D(_11943_),
    .Y(_02353_));
 sg13g2_inv_2 _19893_ (.Y(_02354_),
    .A(net10585));
 sg13g2_nor3_1 _19894_ (.A(_02344_),
    .B(_02354_),
    .C(_11938_),
    .Y(_02355_));
 sg13g2_o21ai_1 _19895_ (.B1(_02350_),
    .Y(_02356_),
    .A1(_02353_),
    .A2(_02355_));
 sg13g2_buf_2 place10332 (.A(_11948_),
    .X(net10332));
 sg13g2_mux2_1 _19897_ (.A0(_00064_),
    .A1(_00067_),
    .S(net10321),
    .X(_02358_));
 sg13g2_inv_2 _19898_ (.Y(_02359_),
    .A(_00072_));
 sg13g2_a22oi_1 _19899_ (.Y(_02360_),
    .B1(net10332),
    .B2(_02359_),
    .A2(net10440),
    .A1(net10575));
 sg13g2_nand2_1 _19900_ (.Y(_02361_),
    .A(net10407),
    .B(_02360_));
 sg13g2_o21ai_1 _19901_ (.B1(_02361_),
    .Y(_02362_),
    .A1(net10406),
    .A2(_02221_));
 sg13g2_o21ai_1 _19902_ (.B1(_02362_),
    .Y(_02363_),
    .A1(net10290),
    .A2(_02358_));
 sg13g2_mux4_1 _19903_ (.S0(net10937),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][14] ),
    .S1(net10920),
    .X(_02364_));
 sg13g2_mux4_1 _19904_ (.S0(net10937),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][14] ),
    .S1(net10920),
    .X(_02365_));
 sg13g2_buf_2 place10346 (.A(net10345),
    .X(net10346));
 sg13g2_buf_2 place10762 (.A(_00004_),
    .X(net10762));
 sg13g2_mux4_1 _19907_ (.S0(net10936),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][14] ),
    .S1(net10920),
    .X(_02368_));
 sg13g2_mux4_1 _19908_ (.S0(net10936),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][14] ),
    .S1(net10920),
    .X(_02369_));
 sg13g2_mux4_1 _19909_ (.S0(net10886),
    .A0(_02364_),
    .A1(_02365_),
    .A2(_02368_),
    .A3(_02369_),
    .S1(net10877),
    .X(_02370_));
 sg13g2_mux4_1 _19910_ (.S0(net10936),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][14] ),
    .S1(net10919),
    .X(_02371_));
 sg13g2_mux4_1 _19911_ (.S0(net10936),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][14] ),
    .S1(net10919),
    .X(_02372_));
 sg13g2_buf_2 place10257 (.A(_06549_),
    .X(net10257));
 sg13g2_mux4_1 _19913_ (.S0(net10936),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][14] ),
    .S1(net10919),
    .X(_02374_));
 sg13g2_mux4_1 _19914_ (.S0(net10936),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][14] ),
    .S1(net10919),
    .X(_02375_));
 sg13g2_mux4_1 _19915_ (.S0(net10886),
    .A0(_02371_),
    .A1(_02372_),
    .A2(_02374_),
    .A3(_02375_),
    .S1(net10869),
    .X(_02376_));
 sg13g2_mux2_1 _19916_ (.A0(_02370_),
    .A1(_02376_),
    .S(net10879),
    .X(_02377_));
 sg13g2_a22oi_1 _19917_ (.Y(_02378_),
    .B1(_02377_),
    .B2(net10267),
    .A2(net10319),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[14] ));
 sg13g2_nor2_1 _19918_ (.A(net10271),
    .B(_02378_),
    .Y(_02379_));
 sg13g2_a21oi_1 _19919_ (.A1(net10703),
    .A2(_02363_),
    .Y(_02380_),
    .B1(_02379_));
 sg13g2_nor2_1 _19920_ (.A(net9666),
    .B(_02380_),
    .Y(_02381_));
 sg13g2_a21oi_1 _19921_ (.A1(net10584),
    .A2(net9665),
    .Y(_02382_),
    .B1(_02381_));
 sg13g2_nand3b_1 _19922_ (.B(_02356_),
    .C(_02382_),
    .Y(_01900_),
    .A_N(_02351_));
 sg13g2_xor2_1 _19923_ (.B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[9] ),
    .A(net10668),
    .X(_02383_));
 sg13g2_xor2_1 _19924_ (.B(net10589),
    .A(net10692),
    .X(_02384_));
 sg13g2_and2_1 _19925_ (.A(net10694),
    .B(net10593),
    .X(_02385_));
 sg13g2_nor2_1 _19926_ (.A(net10694),
    .B(net10593),
    .Y(_02386_));
 sg13g2_xnor2_1 _19927_ (.Y(_02387_),
    .A(net10693),
    .B(net10591));
 sg13g2_nor3_1 _19928_ (.A(_02385_),
    .B(_02386_),
    .C(_02387_),
    .Y(_02388_));
 sg13g2_nor2_1 _19929_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[14] ),
    .B(net10584),
    .Y(_02389_));
 sg13g2_nor2_2 _19930_ (.A(_02344_),
    .B(_02354_),
    .Y(_02390_));
 sg13g2_nor4_1 _19931_ (.A(_02313_),
    .B(_02315_),
    .C(_02389_),
    .D(_02390_),
    .Y(_02391_));
 sg13g2_nand4_1 _19932_ (.B(_02384_),
    .C(_02388_),
    .A(_02383_),
    .Y(_02392_),
    .D(_02391_));
 sg13g2_buf_2 place10347 (.A(net10346),
    .X(net10347));
 sg13g2_a21oi_1 _19934_ (.A1(_12010_),
    .A2(_12028_),
    .Y(_02394_),
    .B1(_02392_));
 sg13g2_inv_1 _19935_ (.Y(_02395_),
    .A(net10692));
 sg13g2_nor2_1 _19936_ (.A(_02395_),
    .B(_08758_),
    .Y(_02396_));
 sg13g2_a22oi_1 _19937_ (.Y(_02397_),
    .B1(net10521),
    .B2(net10668),
    .A2(net10593),
    .A1(net10694));
 sg13g2_o21ai_1 _19938_ (.B1(net10589),
    .Y(_02398_),
    .A1(net10693),
    .A2(net10591));
 sg13g2_nor3_1 _19939_ (.A(_02386_),
    .B(_02397_),
    .C(_02398_),
    .Y(_02399_));
 sg13g2_o21ai_1 _19940_ (.B1(net10692),
    .Y(_02400_),
    .A1(net10693),
    .A2(net10591));
 sg13g2_nor3_1 _19941_ (.A(_02386_),
    .B(_02397_),
    .C(_02400_),
    .Y(_02401_));
 sg13g2_nand2_1 _19942_ (.Y(_02402_),
    .A(net10693),
    .B(net10591));
 sg13g2_a21oi_1 _19943_ (.A1(_02395_),
    .A2(_08758_),
    .Y(_02403_),
    .B1(_02402_));
 sg13g2_nor4_1 _19944_ (.A(_02396_),
    .B(_02399_),
    .C(_02401_),
    .D(_02403_),
    .Y(_02404_));
 sg13g2_o21ai_1 _19945_ (.B1(_02404_),
    .Y(_02405_),
    .A1(_02306_),
    .A2(_08761_));
 sg13g2_nor2_1 _19946_ (.A(_02313_),
    .B(_02389_),
    .Y(_02406_));
 sg13g2_a21o_2 _19947_ (.A2(_02406_),
    .A1(_02405_),
    .B1(_02390_),
    .X(_02407_));
 sg13g2_buf_2 place10340 (.A(_11612_),
    .X(net10340));
 sg13g2_nor2_1 _19949_ (.A(_02394_),
    .B(_02407_),
    .Y(_02409_));
 sg13g2_xnor2_1 _19950_ (.Y(_02410_),
    .A(net10690),
    .B(_02409_));
 sg13g2_nor2_1 _19951_ (.A(net10582),
    .B(net10335),
    .Y(_02411_));
 sg13g2_buf_2 place10268 (.A(net10266),
    .X(net10268));
 sg13g2_nor2_1 _19953_ (.A(_00068_),
    .B(net10406),
    .Y(_02413_));
 sg13g2_a21oi_1 _19954_ (.A1(_02181_),
    .A2(net10406),
    .Y(_02414_),
    .B1(_02413_));
 sg13g2_nand2_1 _19955_ (.Y(_02415_),
    .A(net10573),
    .B(_08310_));
 sg13g2_o21ai_1 _19956_ (.B1(_02415_),
    .Y(_02416_),
    .A1(_00073_),
    .A2(net10438));
 sg13g2_nand2_1 _19957_ (.Y(_02417_),
    .A(net10325),
    .B(_02283_));
 sg13g2_o21ai_1 _19958_ (.B1(_02417_),
    .Y(_02418_),
    .A1(net10325),
    .A2(_02416_));
 sg13g2_o21ai_1 _19959_ (.B1(_02418_),
    .Y(_02419_),
    .A1(net10290),
    .A2(_02414_));
 sg13g2_mux4_1 _19960_ (.S0(net10963),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][15] ),
    .S1(net10899),
    .X(_02420_));
 sg13g2_mux4_1 _19961_ (.S0(net10963),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][15] ),
    .S1(net10899),
    .X(_02421_));
 sg13g2_mux4_1 _19962_ (.S0(net10963),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][15] ),
    .S1(net10899),
    .X(_02422_));
 sg13g2_buf_2 place10256 (.A(_06604_),
    .X(net10256));
 sg13g2_buf_2 place10263 (.A(net10261),
    .X(net10263));
 sg13g2_mux4_1 _19965_ (.S0(net10963),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][15] ),
    .S1(net10899),
    .X(_02425_));
 sg13g2_mux4_1 _19966_ (.S0(net10889),
    .A0(_02420_),
    .A1(_02421_),
    .A2(_02422_),
    .A3(_02425_),
    .S1(net10873),
    .X(_02426_));
 sg13g2_mux4_1 _19967_ (.S0(net10962),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][15] ),
    .S1(net10897),
    .X(_02427_));
 sg13g2_mux4_1 _19968_ (.S0(net10968),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][15] ),
    .S1(net10901),
    .X(_02428_));
 sg13g2_mux4_1 _19969_ (.S0(net10969),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][15] ),
    .S1(net10903),
    .X(_02429_));
 sg13g2_mux4_1 _19970_ (.S0(net10961),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][15] ),
    .S1(net10894),
    .X(_02430_));
 sg13g2_mux4_1 _19971_ (.S0(net10889),
    .A0(_02427_),
    .A1(_02428_),
    .A2(_02429_),
    .A3(_02430_),
    .S1(net10873),
    .X(_02431_));
 sg13g2_mux2_1 _19972_ (.A0(_02426_),
    .A1(_02431_),
    .S(net10882),
    .X(_02432_));
 sg13g2_a22oi_1 _19973_ (.Y(_02433_),
    .B1(_02432_),
    .B2(net10267),
    .A2(net10319),
    .A1(net10496));
 sg13g2_nor2_1 _19974_ (.A(net10271),
    .B(_02433_),
    .Y(_02434_));
 sg13g2_a221oi_1 _19975_ (.B2(net10703),
    .C1(_02434_),
    .B1(_02419_),
    .A1(_02410_),
    .Y(_02435_),
    .A2(_02411_));
 sg13g2_buf_2 place10262 (.A(net10261),
    .X(net10262));
 sg13g2_nor2_1 _19977_ (.A(net10335),
    .B(_02410_),
    .Y(_02437_));
 sg13g2_o21ai_1 _19978_ (.B1(net10582),
    .Y(_02438_),
    .A1(net9666),
    .A2(_02437_));
 sg13g2_o21ai_1 _19979_ (.B1(_02438_),
    .Y(_01901_),
    .A1(net9666),
    .A2(_02435_));
 sg13g2_inv_1 _19980_ (.Y(_02439_),
    .A(net10690));
 sg13g2_nor3_1 _19981_ (.A(net10582),
    .B(_02394_),
    .C(_02407_),
    .Y(_02440_));
 sg13g2_o21ai_1 _19982_ (.B1(net10582),
    .Y(_02441_),
    .A1(_02394_),
    .A2(_02407_));
 sg13g2_o21ai_1 _19983_ (.B1(_02441_),
    .Y(_02442_),
    .A1(_02439_),
    .A2(_02440_));
 sg13g2_xnor2_1 _19984_ (.Y(_02443_),
    .A(net10689),
    .B(_02442_));
 sg13g2_nor2_1 _19985_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[16] ),
    .B(_02443_),
    .Y(_02444_));
 sg13g2_nor2_1 _19986_ (.A(_00069_),
    .B(net10407),
    .Y(_02445_));
 sg13g2_a21oi_1 _19987_ (.A1(_02223_),
    .A2(net10407),
    .Y(_02446_),
    .B1(_02445_));
 sg13g2_nand2_1 _19988_ (.Y(_02447_),
    .A(net10566),
    .B(_08310_));
 sg13g2_o21ai_1 _19989_ (.B1(_02447_),
    .Y(_02448_),
    .A1(_00074_),
    .A2(net10438));
 sg13g2_nand2_1 _19990_ (.Y(_02449_),
    .A(net10327),
    .B(_02338_));
 sg13g2_o21ai_1 _19991_ (.B1(_02449_),
    .Y(_02450_),
    .A1(net10327),
    .A2(_02448_));
 sg13g2_o21ai_1 _19992_ (.B1(_02450_),
    .Y(_02451_),
    .A1(net10290),
    .A2(_02446_));
 sg13g2_buf_2 place10264 (.A(_02336_),
    .X(net10264));
 sg13g2_buf_2 place10327 (.A(net10326),
    .X(net10327));
 sg13g2_mux4_1 _19995_ (.S0(net10961),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][16] ),
    .S1(net10894),
    .X(_02454_));
 sg13g2_mux4_1 _19996_ (.S0(net10960),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][16] ),
    .S1(net10896),
    .X(_02455_));
 sg13g2_mux4_1 _19997_ (.S0(net10960),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][16] ),
    .S1(net10896),
    .X(_02456_));
 sg13g2_mux4_1 _19998_ (.S0(net10960),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][16] ),
    .S1(net10896),
    .X(_02457_));
 sg13g2_mux4_1 _19999_ (.S0(net10888),
    .A0(_02454_),
    .A1(_02455_),
    .A2(_02456_),
    .A3(_02457_),
    .S1(net10872),
    .X(_02458_));
 sg13g2_mux4_1 _20000_ (.S0(net10961),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][16] ),
    .S1(net10894),
    .X(_02459_));
 sg13g2_mux4_1 _20001_ (.S0(net10961),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][16] ),
    .S1(net10894),
    .X(_02460_));
 sg13g2_mux4_1 _20002_ (.S0(net10959),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][16] ),
    .S1(net10896),
    .X(_02461_));
 sg13g2_mux4_1 _20003_ (.S0(net10959),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][16] ),
    .S1(net10896),
    .X(_02462_));
 sg13g2_buf_2 place10429 (.A(net10428),
    .X(net10429));
 sg13g2_mux4_1 _20005_ (.S0(net10888),
    .A0(_02459_),
    .A1(_02460_),
    .A2(_02461_),
    .A3(_02462_),
    .S1(net10872),
    .X(_02464_));
 sg13g2_mux2_1 _20006_ (.A0(_02458_),
    .A1(_02464_),
    .S(net10882),
    .X(_02465_));
 sg13g2_a22oi_1 _20007_ (.Y(_02466_),
    .B1(_02465_),
    .B2(net10267),
    .A2(net10319),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[16] ));
 sg13g2_nor2_1 _20008_ (.A(net10269),
    .B(_02466_),
    .Y(_02467_));
 sg13g2_a221oi_1 _20009_ (.B2(net10703),
    .C1(_02467_),
    .B1(_02451_),
    .A1(_07972_),
    .Y(_02468_),
    .A2(_02444_));
 sg13g2_and2_1 _20010_ (.A(_07972_),
    .B(_02443_),
    .X(_02469_));
 sg13g2_o21ai_1 _20011_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[16] ),
    .Y(_02470_),
    .A1(net9666),
    .A2(_02469_));
 sg13g2_o21ai_1 _20012_ (.B1(_02470_),
    .Y(_01902_),
    .A1(net9666),
    .A2(_02468_));
 sg13g2_a21o_1 _20013_ (.A2(_02442_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[16] ),
    .B1(net10689),
    .X(_02471_));
 sg13g2_or2_1 _20014_ (.X(_02472_),
    .B(_02442_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[16] ));
 sg13g2_nand2_1 _20015_ (.Y(_02473_),
    .A(_02471_),
    .B(_02472_));
 sg13g2_xnor2_1 _20016_ (.Y(_02474_),
    .A(net10688),
    .B(_02473_));
 sg13g2_nor2_1 _20017_ (.A(net10577),
    .B(net10336),
    .Y(_02475_));
 sg13g2_nor2_1 _20018_ (.A(_00067_),
    .B(net10327),
    .Y(_02476_));
 sg13g2_a21oi_1 _20019_ (.A1(_02282_),
    .A2(net10327),
    .Y(_02477_),
    .B1(_02476_));
 sg13g2_nand2_1 _20020_ (.Y(_02478_),
    .A(net10563),
    .B(_08310_));
 sg13g2_o21ai_1 _20021_ (.B1(_02478_),
    .Y(_02479_),
    .A1(_00075_),
    .A2(_08312_));
 sg13g2_nand2_1 _20022_ (.Y(_02480_),
    .A(net10327),
    .B(_02360_));
 sg13g2_o21ai_1 _20023_ (.B1(_02480_),
    .Y(_02481_),
    .A1(net10327),
    .A2(_02479_));
 sg13g2_o21ai_1 _20024_ (.B1(_02481_),
    .Y(_02482_),
    .A1(net10289),
    .A2(_02477_));
 sg13g2_mux4_1 _20025_ (.S0(net10965),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][17] ),
    .S1(net10900),
    .X(_02483_));
 sg13g2_mux4_1 _20026_ (.S0(net10968),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][17] ),
    .S1(net10900),
    .X(_02484_));
 sg13g2_mux4_1 _20027_ (.S0(net10968),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][17] ),
    .S1(net10900),
    .X(_02485_));
 sg13g2_mux4_1 _20028_ (.S0(net10965),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][17] ),
    .S1(net10900),
    .X(_02486_));
 sg13g2_mux4_1 _20029_ (.S0(net10890),
    .A0(_02483_),
    .A1(_02484_),
    .A2(_02485_),
    .A3(_02486_),
    .S1(net10874),
    .X(_02487_));
 sg13g2_mux4_1 _20030_ (.S0(net10968),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][17] ),
    .S1(net10901),
    .X(_02488_));
 sg13g2_mux4_1 _20031_ (.S0(net10968),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][17] ),
    .S1(net10901),
    .X(_02489_));
 sg13g2_mux4_1 _20032_ (.S0(net10966),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][17] ),
    .S1(net10904),
    .X(_02490_));
 sg13g2_mux4_1 _20033_ (.S0(net10970),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][17] ),
    .S1(net10907),
    .X(_02491_));
 sg13g2_buf_2 place10253 (.A(_07207_),
    .X(net10253));
 sg13g2_mux4_1 _20035_ (.S0(net10890),
    .A0(_02488_),
    .A1(_02489_),
    .A2(_02490_),
    .A3(_02491_),
    .S1(net10874),
    .X(_02493_));
 sg13g2_buf_2 place10391 (.A(net10390),
    .X(net10391));
 sg13g2_mux2_1 _20037_ (.A0(_02487_),
    .A1(_02493_),
    .S(net10881),
    .X(_02495_));
 sg13g2_a22oi_1 _20038_ (.Y(_02496_),
    .B1(_02495_),
    .B2(net10267),
    .A2(net10319),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[17] ));
 sg13g2_nor2_1 _20039_ (.A(net10269),
    .B(_02496_),
    .Y(_02497_));
 sg13g2_a221oi_1 _20040_ (.B2(net10706),
    .C1(_02497_),
    .B1(_02482_),
    .A1(_02474_),
    .Y(_02498_),
    .A2(_02475_));
 sg13g2_nor2_1 _20041_ (.A(net10335),
    .B(_02474_),
    .Y(_02499_));
 sg13g2_o21ai_1 _20042_ (.B1(net10577),
    .Y(_02500_),
    .A1(net9667),
    .A2(_02499_));
 sg13g2_o21ai_1 _20043_ (.B1(_02500_),
    .Y(_01903_),
    .A1(net9667),
    .A2(_02498_));
 sg13g2_a22oi_1 _20044_ (.Y(_02501_),
    .B1(_02471_),
    .B2(_02472_),
    .A2(net10577),
    .A1(net10688));
 sg13g2_nor2_1 _20045_ (.A(net10688),
    .B(net10577),
    .Y(_02502_));
 sg13g2_o21ai_1 _20046_ (.B1(net10687),
    .Y(_02503_),
    .A1(_02501_),
    .A2(_02502_));
 sg13g2_or3_1 _20047_ (.A(net10687),
    .B(_02501_),
    .C(_02502_),
    .X(_02504_));
 sg13g2_a21oi_1 _20048_ (.A1(_02503_),
    .A2(_02504_),
    .Y(_02505_),
    .B1(net10575));
 sg13g2_buf_2 place10278 (.A(net10277),
    .X(net10278));
 sg13g2_buf_2 place10328 (.A(net10326),
    .X(net10328));
 sg13g2_mux4_1 _20051_ (.S0(net10953),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][18] ),
    .S1(net10915),
    .X(_02508_));
 sg13g2_mux4_1 _20052_ (.S0(net10957),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][18] ),
    .S1(net10918),
    .X(_02509_));
 sg13g2_buf_2 place10251 (.A(net10248),
    .X(net10251));
 sg13g2_buf_2 place10378 (.A(net10376),
    .X(net10378));
 sg13g2_mux4_1 _20055_ (.S0(net10955),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][18] ),
    .S1(net10914),
    .X(_02512_));
 sg13g2_mux4_1 _20056_ (.S0(net10950),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][18] ),
    .S1(net10911),
    .X(_02513_));
 sg13g2_buf_2 place10246 (.A(_07924_),
    .X(net10246));
 sg13g2_mux4_1 _20058_ (.S0(net10887),
    .A0(_02508_),
    .A1(_02509_),
    .A2(_02512_),
    .A3(_02513_),
    .S1(net10876),
    .X(_02515_));
 sg13g2_mux4_1 _20059_ (.S0(net10955),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][18] ),
    .S1(net10914),
    .X(_02516_));
 sg13g2_mux4_1 _20060_ (.S0(net10953),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][18] ),
    .S1(_00006_),
    .X(_02517_));
 sg13g2_mux4_1 _20061_ (.S0(net10953),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][18] ),
    .S1(net10915),
    .X(_02518_));
 sg13g2_mux4_1 _20062_ (.S0(net10953),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][18] ),
    .S1(net10915),
    .X(_02519_));
 sg13g2_mux4_1 _20063_ (.S0(net10887),
    .A0(_02516_),
    .A1(_02517_),
    .A2(_02518_),
    .A3(_02519_),
    .S1(net10876),
    .X(_02520_));
 sg13g2_mux2_1 _20064_ (.A0(_02515_),
    .A1(_02520_),
    .S(net10880),
    .X(_02521_));
 sg13g2_a22oi_1 _20065_ (.Y(_02522_),
    .B1(_02521_),
    .B2(net10267),
    .A2(net10317),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[18] ));
 sg13g2_nor2_1 _20066_ (.A(net10294),
    .B(_02522_),
    .Y(_02523_));
 sg13g2_buf_2 place10236 (.A(net10235),
    .X(net10236));
 sg13g2_buf_16 clkbuf_leaf_318_clk (.X(clknet_leaf_318_clk),
    .A(clknet_8_89_0_clk));
 sg13g2_nand2_1 _20069_ (.Y(_02526_),
    .A(_02337_),
    .B(net10326));
 sg13g2_o21ai_1 _20070_ (.B1(_02526_),
    .Y(_02527_),
    .A1(_00068_),
    .A2(net10327));
 sg13g2_buf_2 place10233 (.A(net10231),
    .X(net10233));
 sg13g2_nand2_1 _20072_ (.Y(_02529_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[22] ),
    .B(_08310_));
 sg13g2_o21ai_1 _20073_ (.B1(_02529_),
    .Y(_02530_),
    .A1(_00076_),
    .A2(net10439));
 sg13g2_and2_1 _20074_ (.A(net10408),
    .B(_02530_),
    .X(_02531_));
 sg13g2_a221oi_1 _20075_ (.B2(_02336_),
    .C1(_02531_),
    .B1(_02527_),
    .A1(net10328),
    .Y(_02532_),
    .A2(_02416_));
 sg13g2_nor2_1 _20076_ (.A(net10392),
    .B(_02532_),
    .Y(_02533_));
 sg13g2_a221oi_1 _20077_ (.B2(net10392),
    .C1(_02533_),
    .B1(_02523_),
    .A1(net10294),
    .Y(_02534_),
    .A2(_02505_));
 sg13g2_and3_1 _20078_ (.X(_02535_),
    .A(net10294),
    .B(_02503_),
    .C(_02504_));
 sg13g2_o21ai_1 _20079_ (.B1(net10575),
    .Y(_02536_),
    .A1(net9667),
    .A2(_02535_));
 sg13g2_o21ai_1 _20080_ (.B1(_02536_),
    .Y(_01904_),
    .A1(net9667),
    .A2(_02534_));
 sg13g2_mux4_1 _20081_ (.S0(net10942),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][19] ),
    .S1(net10927),
    .X(_02537_));
 sg13g2_mux4_1 _20082_ (.S0(net10942),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][19] ),
    .S1(net10927),
    .X(_02538_));
 sg13g2_mux4_1 _20083_ (.S0(net10943),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][19] ),
    .S1(net10928),
    .X(_02539_));
 sg13g2_mux4_1 _20084_ (.S0(net10942),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][19] ),
    .S1(net10927),
    .X(_02540_));
 sg13g2_mux4_1 _20085_ (.S0(_00007_),
    .A0(_02537_),
    .A1(_02538_),
    .A2(_02539_),
    .A3(_02540_),
    .S1(net10870),
    .X(_02541_));
 sg13g2_mux4_1 _20086_ (.S0(net10944),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][19] ),
    .S1(net10929),
    .X(_02542_));
 sg13g2_mux4_1 _20087_ (.S0(net10944),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][19] ),
    .S1(net10929),
    .X(_02543_));
 sg13g2_mux4_1 _20088_ (.S0(net10946),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][19] ),
    .S1(net10931),
    .X(_02544_));
 sg13g2_mux4_1 _20089_ (.S0(net10946),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][19] ),
    .S1(net10931),
    .X(_02545_));
 sg13g2_mux4_1 _20090_ (.S0(net10883),
    .A0(_02542_),
    .A1(_02543_),
    .A2(_02544_),
    .A3(_02545_),
    .S1(net10870),
    .X(_02546_));
 sg13g2_mux2_1 _20091_ (.A0(_02541_),
    .A1(_02546_),
    .S(net10878),
    .X(_02547_));
 sg13g2_a22oi_1 _20092_ (.Y(_02548_),
    .B1(_02547_),
    .B2(net10265),
    .A2(net10318),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[19] ));
 sg13g2_nor2_1 _20093_ (.A(net10294),
    .B(_02548_),
    .Y(_02549_));
 sg13g2_nor2_1 _20094_ (.A(net10687),
    .B(net10575),
    .Y(_02550_));
 sg13g2_nor2_1 _20095_ (.A(net10689),
    .B(net10579),
    .Y(_02551_));
 sg13g2_a22oi_1 _20096_ (.Y(_02552_),
    .B1(net10579),
    .B2(net10689),
    .A2(net10582),
    .A1(net10690));
 sg13g2_o21ai_1 _20097_ (.B1(_08653_),
    .Y(_02553_),
    .A1(_02551_),
    .A2(_02552_));
 sg13g2_nor3_1 _20098_ (.A(_08653_),
    .B(_02551_),
    .C(_02552_),
    .Y(_02554_));
 sg13g2_a221oi_1 _20099_ (.B2(net10688),
    .C1(_02554_),
    .B1(_02553_),
    .A1(net10687),
    .Y(_02555_),
    .A2(net10575));
 sg13g2_nor2_2 _20100_ (.A(_02550_),
    .B(_02555_),
    .Y(_02556_));
 sg13g2_a21oi_2 _20101_ (.B1(_02390_),
    .Y(_02557_),
    .A2(_02406_),
    .A1(_02405_));
 sg13g2_xor2_1 _20102_ (.B(net10577),
    .A(net10688),
    .X(_02558_));
 sg13g2_xor2_1 _20103_ (.B(net10582),
    .A(net10690),
    .X(_02559_));
 sg13g2_and2_1 _20104_ (.A(net10687),
    .B(net10575),
    .X(_02560_));
 sg13g2_and2_1 _20105_ (.A(net10689),
    .B(net10579),
    .X(_02561_));
 sg13g2_nor4_1 _20106_ (.A(_02550_),
    .B(_02560_),
    .C(_02551_),
    .D(_02561_),
    .Y(_02562_));
 sg13g2_nand3_1 _20107_ (.B(_02559_),
    .C(_02562_),
    .A(_02558_),
    .Y(_02563_));
 sg13g2_buf_16 clkbuf_leaf_317_clk (.X(clknet_leaf_317_clk),
    .A(clknet_8_92_0_clk));
 sg13g2_nor2_2 _20109_ (.A(_02557_),
    .B(_02563_),
    .Y(_02565_));
 sg13g2_or2_1 _20110_ (.X(_02566_),
    .B(_02563_),
    .A(_02392_));
 sg13g2_a21oi_2 _20111_ (.B1(_02566_),
    .Y(_02567_),
    .A2(_12028_),
    .A1(_12010_));
 sg13g2_nor3_2 _20112_ (.A(_02556_),
    .B(_02565_),
    .C(_02567_),
    .Y(_02568_));
 sg13g2_xnor2_1 _20113_ (.Y(_02569_),
    .A(net10686),
    .B(_02568_));
 sg13g2_nor2_1 _20114_ (.A(net10573),
    .B(net10336),
    .Y(_02570_));
 sg13g2_nand2_1 _20115_ (.Y(_02571_),
    .A(_02359_),
    .B(net10328));
 sg13g2_o21ai_1 _20116_ (.B1(_02571_),
    .Y(_02572_),
    .A1(_00069_),
    .A2(net10328));
 sg13g2_nand2_1 _20117_ (.Y(_02573_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[23] ),
    .B(net10443));
 sg13g2_o21ai_1 _20118_ (.B1(_02573_),
    .Y(_02574_),
    .A1(_00077_),
    .A2(net10439));
 sg13g2_and2_1 _20119_ (.A(net10408),
    .B(_02574_),
    .X(_02575_));
 sg13g2_a221oi_1 _20120_ (.B2(_02336_),
    .C1(_02575_),
    .B1(_02572_),
    .A1(net10328),
    .Y(_02576_),
    .A2(_02448_));
 sg13g2_nor2_1 _20121_ (.A(net10392),
    .B(_02576_),
    .Y(_02577_));
 sg13g2_a221oi_1 _20122_ (.B2(_02570_),
    .C1(_02577_),
    .B1(_02569_),
    .A1(net10392),
    .Y(_02578_),
    .A2(_02549_));
 sg13g2_nor2_1 _20123_ (.A(net10336),
    .B(_02569_),
    .Y(_02579_));
 sg13g2_o21ai_1 _20124_ (.B1(net10573),
    .Y(_02580_),
    .A1(net9667),
    .A2(_02579_));
 sg13g2_o21ai_1 _20125_ (.B1(_02580_),
    .Y(_01905_),
    .A1(net9667),
    .A2(_02578_));
 sg13g2_buf_2 place10379 (.A(_11410_),
    .X(net10379));
 sg13g2_buf_2 place10235 (.A(net10234),
    .X(net10235));
 sg13g2_mux4_1 _20128_ (.S0(net10971),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][1] ),
    .S1(net10907),
    .X(_02583_));
 sg13g2_mux4_1 _20129_ (.S0(net10971),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][1] ),
    .S1(net10907),
    .X(_02584_));
 sg13g2_buf_2 place10393 (.A(_09453_),
    .X(net10393));
 sg13g2_buf_2 place10234 (.A(_07931_),
    .X(net10234));
 sg13g2_mux4_1 _20132_ (.S0(net10971),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][1] ),
    .S1(net10907),
    .X(_02587_));
 sg13g2_mux4_1 _20133_ (.S0(net10964),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][1] ),
    .S1(net10905),
    .X(_02588_));
 sg13g2_mux4_1 _20134_ (.S0(net10890),
    .A0(_02583_),
    .A1(_02584_),
    .A2(_02587_),
    .A3(_02588_),
    .S1(net10874),
    .X(_02589_));
 sg13g2_mux4_1 _20135_ (.S0(net10971),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][1] ),
    .S1(net10907),
    .X(_02590_));
 sg13g2_mux4_1 _20136_ (.S0(net10973),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][1] ),
    .S1(net10910),
    .X(_02591_));
 sg13g2_mux4_1 _20137_ (.S0(net10973),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][1] ),
    .S1(net10910),
    .X(_02592_));
 sg13g2_mux4_1 _20138_ (.S0(net10964),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][1] ),
    .S1(net10905),
    .X(_02593_));
 sg13g2_mux4_1 _20139_ (.S0(net10890),
    .A0(_02590_),
    .A1(_02591_),
    .A2(_02592_),
    .A3(_02593_),
    .S1(net10874),
    .X(_02594_));
 sg13g2_mux2_1 _20140_ (.A0(_02589_),
    .A1(_02594_),
    .S(net10881),
    .X(_02595_));
 sg13g2_a22oi_1 _20141_ (.Y(_02596_),
    .B1(_02595_),
    .B2(net10268),
    .A2(net10320),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[1] ));
 sg13g2_inv_1 _20142_ (.Y(_02597_),
    .A(_00058_));
 sg13g2_a22oi_1 _20143_ (.Y(_02598_),
    .B1(net10331),
    .B2(_02597_),
    .A2(net10442),
    .A1(net10528));
 sg13g2_inv_2 _20144_ (.Y(_02599_),
    .A(_00057_));
 sg13g2_a22oi_1 _20145_ (.Y(_02600_),
    .B1(net10331),
    .B2(_02599_),
    .A2(net10442),
    .A1(net10538));
 sg13g2_o21ai_1 _20146_ (.B1(_02600_),
    .Y(_02601_),
    .A1(_00056_),
    .A2(net10289));
 sg13g2_nand2_1 _20147_ (.Y(_02602_),
    .A(net10323),
    .B(_02601_));
 sg13g2_o21ai_1 _20148_ (.B1(_02602_),
    .Y(_02603_),
    .A1(net10324),
    .A2(_02598_));
 sg13g2_nand2_1 _20149_ (.Y(_02604_),
    .A(net10595),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[0] ));
 sg13g2_xor2_1 _20150_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[1] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[1] ),
    .X(_02605_));
 sg13g2_xnor2_1 _20151_ (.Y(_02606_),
    .A(_02604_),
    .B(_02605_));
 sg13g2_a22oi_1 _20152_ (.Y(_02607_),
    .B1(_02606_),
    .B2(net10293),
    .A2(_02603_),
    .A1(net10702));
 sg13g2_o21ai_1 _20153_ (.B1(_02607_),
    .Y(_02608_),
    .A1(net10272),
    .A2(_02596_));
 sg13g2_nor2_1 _20154_ (.A(net9673),
    .B(_02608_),
    .Y(_02609_));
 sg13g2_a21oi_1 _20155_ (.A1(net10400),
    .A2(net9673),
    .Y(_01906_),
    .B1(_02609_));
 sg13g2_buf_2 place10237 (.A(net10236),
    .X(net10237));
 sg13g2_inv_4 _20157_ (.A(net10573),
    .Y(_02611_));
 sg13g2_or2_1 _20158_ (.X(_02612_),
    .B(_02563_),
    .A(_02611_));
 sg13g2_or2_1 _20159_ (.X(_02613_),
    .B(_02612_),
    .A(_02392_));
 sg13g2_a21oi_1 _20160_ (.A1(_12010_),
    .A2(_12028_),
    .Y(_02614_),
    .B1(_02613_));
 sg13g2_nand2_1 _20161_ (.Y(_02615_),
    .A(net10573),
    .B(_02556_));
 sg13g2_o21ai_1 _20162_ (.B1(_02615_),
    .Y(_02616_),
    .A1(_02557_),
    .A2(_02612_));
 sg13g2_nor3_2 _20163_ (.A(net10686),
    .B(_02614_),
    .C(_02616_),
    .Y(_02617_));
 sg13g2_nor4_1 _20164_ (.A(net10573),
    .B(_02556_),
    .C(_02565_),
    .D(_02567_),
    .Y(_02618_));
 sg13g2_or2_1 _20165_ (.X(_02619_),
    .B(_02618_),
    .A(_02617_));
 sg13g2_buf_16 clkbuf_leaf_316_clk (.X(clknet_leaf_316_clk),
    .A(clknet_8_89_0_clk));
 sg13g2_xnor2_1 _20167_ (.Y(_02621_),
    .A(net10685),
    .B(_02619_));
 sg13g2_nor2_1 _20168_ (.A(net10566),
    .B(net10336),
    .Y(_02622_));
 sg13g2_nand2_1 _20169_ (.Y(_02623_),
    .A(_00070_),
    .B(net10407));
 sg13g2_nand2_1 _20170_ (.Y(_02624_),
    .A(_00073_),
    .B(net10328));
 sg13g2_nand3_1 _20171_ (.B(_02623_),
    .C(_02624_),
    .A(_02336_),
    .Y(_02625_));
 sg13g2_nand2_1 _20172_ (.Y(_02626_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[24] ),
    .B(net10443));
 sg13g2_o21ai_1 _20173_ (.B1(_02626_),
    .Y(_02627_),
    .A1(_00078_),
    .A2(net10439));
 sg13g2_nand2_1 _20174_ (.Y(_02628_),
    .A(net10409),
    .B(_02627_));
 sg13g2_nand2_1 _20175_ (.Y(_02629_),
    .A(net10328),
    .B(_02479_));
 sg13g2_nand3_1 _20176_ (.B(_02628_),
    .C(_02629_),
    .A(_02625_),
    .Y(_02630_));
 sg13g2_mux4_1 _20177_ (.S0(net10953),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][20] ),
    .S1(net10915),
    .X(_02631_));
 sg13g2_mux4_1 _20178_ (.S0(net10957),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][20] ),
    .S1(net10918),
    .X(_02632_));
 sg13g2_buf_2 place10415 (.A(net10414),
    .X(net10415));
 sg13g2_buf_2 place10398 (.A(net10397),
    .X(net10398));
 sg13g2_mux4_1 _20181_ (.S0(net10955),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][20] ),
    .S1(net10914),
    .X(_02635_));
 sg13g2_mux4_1 _20182_ (.S0(net10950),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][20] ),
    .S1(net10911),
    .X(_02636_));
 sg13g2_mux4_1 _20183_ (.S0(net10887),
    .A0(_02631_),
    .A1(_02632_),
    .A2(_02635_),
    .A3(_02636_),
    .S1(net10876),
    .X(_02637_));
 sg13g2_mux4_1 _20184_ (.S0(net10952),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][20] ),
    .S1(net10914),
    .X(_02638_));
 sg13g2_mux4_1 _20185_ (.S0(net10952),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][20] ),
    .S1(net10914),
    .X(_02639_));
 sg13g2_mux4_1 _20186_ (.S0(net10952),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][20] ),
    .S1(net10914),
    .X(_02640_));
 sg13g2_mux4_1 _20187_ (.S0(net10952),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][20] ),
    .S1(net10914),
    .X(_02641_));
 sg13g2_mux4_1 _20188_ (.S0(net10887),
    .A0(_02638_),
    .A1(_02639_),
    .A2(_02640_),
    .A3(_02641_),
    .S1(net10876),
    .X(_02642_));
 sg13g2_mux2_1 _20189_ (.A0(_02637_),
    .A1(_02642_),
    .S(net10880),
    .X(_02643_));
 sg13g2_buf_2 place10231 (.A(_07979_),
    .X(net10231));
 sg13g2_a22oi_1 _20191_ (.Y(_02645_),
    .B1(_02643_),
    .B2(net10267),
    .A2(net10317),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[20] ));
 sg13g2_nor2_1 _20192_ (.A(net10269),
    .B(_02645_),
    .Y(_02646_));
 sg13g2_a221oi_1 _20193_ (.B2(net10706),
    .C1(_02646_),
    .B1(_02630_),
    .A1(_02621_),
    .Y(_02647_),
    .A2(_02622_));
 sg13g2_nor2_1 _20194_ (.A(net10336),
    .B(_02621_),
    .Y(_02648_));
 sg13g2_o21ai_1 _20195_ (.B1(net10566),
    .Y(_02649_),
    .A1(net9668),
    .A2(_02648_));
 sg13g2_o21ai_1 _20196_ (.B1(_02649_),
    .Y(_01907_),
    .A1(net9668),
    .A2(_02647_));
 sg13g2_inv_4 _20197_ (.A(net10566),
    .Y(_02650_));
 sg13g2_o21ai_1 _20198_ (.B1(_02650_),
    .Y(_02651_),
    .A1(_02617_),
    .A2(_02618_));
 sg13g2_or4_1 _20199_ (.A(net10686),
    .B(net10685),
    .C(_02614_),
    .D(_02616_),
    .X(_02652_));
 sg13g2_inv_1 _20200_ (.Y(_02653_),
    .A(net10685));
 sg13g2_nand2_1 _20201_ (.Y(_02654_),
    .A(_02653_),
    .B(_02611_));
 sg13g2_or4_1 _20202_ (.A(_02556_),
    .B(_02565_),
    .C(_02567_),
    .D(_02654_),
    .X(_02655_));
 sg13g2_nand2_1 _20203_ (.Y(_02656_),
    .A(_02653_),
    .B(_02650_));
 sg13g2_and3_1 _20204_ (.X(_02657_),
    .A(_02652_),
    .B(_02655_),
    .C(_02656_));
 sg13g2_nand2_1 _20205_ (.Y(_02658_),
    .A(_02651_),
    .B(_02657_));
 sg13g2_xnor2_1 _20206_ (.Y(_02659_),
    .A(net10684),
    .B(_02658_));
 sg13g2_nor2_1 _20207_ (.A(net10563),
    .B(net10336),
    .Y(_02660_));
 sg13g2_nand2_1 _20208_ (.Y(_02661_),
    .A(_00071_),
    .B(net10408));
 sg13g2_nand2_1 _20209_ (.Y(_02662_),
    .A(_00074_),
    .B(net10328));
 sg13g2_nand3_1 _20210_ (.B(_02661_),
    .C(_02662_),
    .A(_02336_),
    .Y(_02663_));
 sg13g2_nand2_1 _20211_ (.Y(_02664_),
    .A(net10551),
    .B(net10443));
 sg13g2_o21ai_1 _20212_ (.B1(_02664_),
    .Y(_02665_),
    .A1(_00079_),
    .A2(net10439));
 sg13g2_nand2_1 _20213_ (.Y(_02666_),
    .A(net10409),
    .B(_02665_));
 sg13g2_nand2_1 _20214_ (.Y(_02667_),
    .A(net10328),
    .B(_02530_));
 sg13g2_nand3_1 _20215_ (.B(_02666_),
    .C(_02667_),
    .A(_02663_),
    .Y(_02668_));
 sg13g2_buf_2 place10331 (.A(_11948_),
    .X(net10331));
 sg13g2_buf_2 place10341 (.A(net10340),
    .X(net10341));
 sg13g2_mux4_1 _20218_ (.S0(net10953),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][21] ),
    .S1(net10915),
    .X(_02671_));
 sg13g2_mux4_1 _20219_ (.S0(net10957),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][21] ),
    .S1(net10918),
    .X(_02672_));
 sg13g2_mux4_1 _20220_ (.S0(net10955),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][21] ),
    .S1(net10914),
    .X(_02673_));
 sg13g2_mux4_1 _20221_ (.S0(net10950),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][21] ),
    .S1(net10911),
    .X(_02674_));
 sg13g2_mux4_1 _20222_ (.S0(net10887),
    .A0(_02671_),
    .A1(_02672_),
    .A2(_02673_),
    .A3(_02674_),
    .S1(net10876),
    .X(_02675_));
 sg13g2_mux4_1 _20223_ (.S0(net10957),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][21] ),
    .S1(net10918),
    .X(_02676_));
 sg13g2_buf_2 place10353 (.A(_11605_),
    .X(net10353));
 sg13g2_buf_2 place10227 (.A(net10226),
    .X(net10227));
 sg13g2_mux4_1 _20226_ (.S0(net10957),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][21] ),
    .S1(net10918),
    .X(_02679_));
 sg13g2_mux4_1 _20227_ (.S0(net10957),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][21] ),
    .S1(net10918),
    .X(_02680_));
 sg13g2_mux4_1 _20228_ (.S0(net10957),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][21] ),
    .S1(net10918),
    .X(_02681_));
 sg13g2_mux4_1 _20229_ (.S0(net10887),
    .A0(_02676_),
    .A1(_02679_),
    .A2(_02680_),
    .A3(_02681_),
    .S1(net10876),
    .X(_02682_));
 sg13g2_mux2_1 _20230_ (.A0(_02675_),
    .A1(_02682_),
    .S(net10880),
    .X(_02683_));
 sg13g2_a22oi_1 _20231_ (.Y(_02684_),
    .B1(_02683_),
    .B2(net10266),
    .A2(net10317),
    .A1(net10495));
 sg13g2_nor2_1 _20232_ (.A(net10269),
    .B(_02684_),
    .Y(_02685_));
 sg13g2_a221oi_1 _20233_ (.B2(net10706),
    .C1(_02685_),
    .B1(_02668_),
    .A1(_02659_),
    .Y(_02686_),
    .A2(_02660_));
 sg13g2_nor2_1 _20234_ (.A(net10336),
    .B(_02659_),
    .Y(_02687_));
 sg13g2_o21ai_1 _20235_ (.B1(net10563),
    .Y(_02688_),
    .A1(net9668),
    .A2(_02687_));
 sg13g2_o21ai_1 _20236_ (.B1(_02688_),
    .Y(_01908_),
    .A1(net9668),
    .A2(_02686_));
 sg13g2_or2_1 _20237_ (.X(_02689_),
    .B(net10562),
    .A(net10684));
 sg13g2_and2_1 _20238_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[20] ),
    .B(net10566),
    .X(_02690_));
 sg13g2_buf_2 place10232 (.A(net10231),
    .X(net10232));
 sg13g2_and2_1 _20240_ (.A(net10684),
    .B(net10562),
    .X(_02692_));
 sg13g2_buf_2 place10307 (.A(net10306),
    .X(net10307));
 sg13g2_a21o_1 _20242_ (.A2(_02690_),
    .A1(_02689_),
    .B1(_02692_),
    .X(_02694_));
 sg13g2_nand2_1 _20243_ (.Y(_02695_),
    .A(net10563),
    .B(net10566));
 sg13g2_nand2_1 _20244_ (.Y(_02696_),
    .A(net10685),
    .B(net10563));
 sg13g2_a221oi_1 _20245_ (.B2(_02696_),
    .C1(_02617_),
    .B1(_02695_),
    .A1(_02611_),
    .Y(_02697_),
    .A2(_02568_));
 sg13g2_nand2_1 _20246_ (.Y(_02698_),
    .A(net10684),
    .B(net10566));
 sg13g2_nand2_1 _20247_ (.Y(_02699_),
    .A(net10685),
    .B(net10684));
 sg13g2_a221oi_1 _20248_ (.B2(_02699_),
    .C1(_02617_),
    .B1(_02698_),
    .A1(_02611_),
    .Y(_02700_),
    .A2(_02568_));
 sg13g2_nor3_2 _20249_ (.A(_02694_),
    .B(_02697_),
    .C(_02700_),
    .Y(_02701_));
 sg13g2_xnor2_1 _20250_ (.Y(_02702_),
    .A(net10682),
    .B(_02701_));
 sg13g2_nor2_1 _20251_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[22] ),
    .B(net10338),
    .Y(_02703_));
 sg13g2_nor2_1 _20252_ (.A(_00075_),
    .B(net10408),
    .Y(_02704_));
 sg13g2_a21oi_1 _20253_ (.A1(_02359_),
    .A2(net10408),
    .Y(_02705_),
    .B1(_02704_));
 sg13g2_inv_1 _20254_ (.Y(_02706_),
    .A(_00080_));
 sg13g2_a22oi_1 _20255_ (.Y(_02707_),
    .B1(net10332),
    .B2(_02706_),
    .A2(net10443),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[26] ));
 sg13g2_nand2_1 _20256_ (.Y(_02708_),
    .A(net10408),
    .B(_02707_));
 sg13g2_o21ai_1 _20257_ (.B1(_02708_),
    .Y(_02709_),
    .A1(net10408),
    .A2(_02574_));
 sg13g2_o21ai_1 _20258_ (.B1(_02709_),
    .Y(_02710_),
    .A1(_08314_),
    .A2(_02705_));
 sg13g2_mux4_1 _20259_ (.S0(net10938),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][22] ),
    .S1(net10922),
    .X(_02711_));
 sg13g2_mux4_1 _20260_ (.S0(net10938),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][22] ),
    .S1(net10922),
    .X(_02712_));
 sg13g2_mux4_1 _20261_ (.S0(net10938),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][22] ),
    .S1(net10922),
    .X(_02713_));
 sg13g2_mux4_1 _20262_ (.S0(net10938),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][22] ),
    .S1(net10922),
    .X(_02714_));
 sg13g2_mux4_1 _20263_ (.S0(net10892),
    .A0(_02711_),
    .A1(_02712_),
    .A2(_02713_),
    .A3(_02714_),
    .S1(net10877),
    .X(_02715_));
 sg13g2_mux4_1 _20264_ (.S0(net10951),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][22] ),
    .S1(net10913),
    .X(_02716_));
 sg13g2_mux4_1 _20265_ (.S0(net10951),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][22] ),
    .S1(net10913),
    .X(_02717_));
 sg13g2_mux4_1 _20266_ (.S0(net10951),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][22] ),
    .S1(net10913),
    .X(_02718_));
 sg13g2_mux4_1 _20267_ (.S0(net10951),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][22] ),
    .S1(net10913),
    .X(_02719_));
 sg13g2_mux4_1 _20268_ (.S0(net10892),
    .A0(_02716_),
    .A1(_02717_),
    .A2(_02718_),
    .A3(_02719_),
    .S1(net10877),
    .X(_02720_));
 sg13g2_mux2_1 _20269_ (.A0(_02715_),
    .A1(_02720_),
    .S(net10880),
    .X(_02721_));
 sg13g2_a22oi_1 _20270_ (.Y(_02722_),
    .B1(_02721_),
    .B2(_11988_),
    .A2(net10317),
    .A1(net10494));
 sg13g2_nor2_1 _20271_ (.A(net10269),
    .B(_02722_),
    .Y(_02723_));
 sg13g2_a221oi_1 _20272_ (.B2(net10706),
    .C1(_02723_),
    .B1(_02710_),
    .A1(_02702_),
    .Y(_02724_),
    .A2(_02703_));
 sg13g2_buf_2 place10333 (.A(_11938_),
    .X(net10333));
 sg13g2_nor2_1 _20274_ (.A(net10336),
    .B(_02702_),
    .Y(_02726_));
 sg13g2_o21ai_1 _20275_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[22] ),
    .Y(_02727_),
    .A1(net9668),
    .A2(_02726_));
 sg13g2_o21ai_1 _20276_ (.B1(_02727_),
    .Y(_01909_),
    .A1(net9668),
    .A2(_02724_));
 sg13g2_nand2b_1 _20277_ (.Y(_02728_),
    .B(_02701_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[22] ));
 sg13g2_nor2b_1 _20278_ (.A(_02701_),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[22] ),
    .Y(_02729_));
 sg13g2_a21oi_1 _20279_ (.A1(net10682),
    .A2(_02728_),
    .Y(_02730_),
    .B1(_02729_));
 sg13g2_xnor2_1 _20280_ (.Y(_02731_),
    .A(_09675_),
    .B(_02730_));
 sg13g2_nand3_1 _20281_ (.B(net10294),
    .C(_02731_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[23] ),
    .Y(_02732_));
 sg13g2_or4_1 _20282_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[23] ),
    .B(net10338),
    .C(net9669),
    .D(_02731_),
    .X(_02733_));
 sg13g2_inv_1 _20283_ (.Y(_02734_),
    .A(_00076_));
 sg13g2_nor2_1 _20284_ (.A(_00073_),
    .B(net10329),
    .Y(_02735_));
 sg13g2_a21oi_1 _20285_ (.A1(_02734_),
    .A2(net10329),
    .Y(_02736_),
    .B1(_02735_));
 sg13g2_nand2_1 _20286_ (.Y(_02737_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[27] ),
    .B(net10443));
 sg13g2_o21ai_1 _20287_ (.B1(_02737_),
    .Y(_02738_),
    .A1(_00081_),
    .A2(net10439));
 sg13g2_nor2_1 _20288_ (.A(net10264),
    .B(net10329),
    .Y(_02739_));
 sg13g2_a22oi_1 _20289_ (.Y(_02740_),
    .B1(_02738_),
    .B2(_02739_),
    .A2(_02627_),
    .A1(net10329));
 sg13g2_o21ai_1 _20290_ (.B1(_02740_),
    .Y(_02741_),
    .A1(_08314_),
    .A2(_02736_));
 sg13g2_mux4_1 _20291_ (.S0(net10937),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][23] ),
    .S1(net10921),
    .X(_02742_));
 sg13g2_mux4_1 _20292_ (.S0(net10937),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][23] ),
    .S1(net10921),
    .X(_02743_));
 sg13g2_mux4_1 _20293_ (.S0(net10937),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][23] ),
    .S1(net10921),
    .X(_02744_));
 sg13g2_mux4_1 _20294_ (.S0(net10937),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][23] ),
    .S1(net10921),
    .X(_02745_));
 sg13g2_mux4_1 _20295_ (.S0(net10886),
    .A0(_02742_),
    .A1(_02743_),
    .A2(_02744_),
    .A3(_02745_),
    .S1(net10877),
    .X(_02746_));
 sg13g2_mux4_1 _20296_ (.S0(net10950),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][23] ),
    .S1(net10912),
    .X(_02747_));
 sg13g2_mux4_1 _20297_ (.S0(net10952),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][23] ),
    .S1(net10912),
    .X(_02748_));
 sg13g2_mux4_1 _20298_ (.S0(net10952),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][23] ),
    .S1(net10912),
    .X(_02749_));
 sg13g2_mux4_1 _20299_ (.S0(net10952),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][23] ),
    .S1(net10912),
    .X(_02750_));
 sg13g2_mux4_1 _20300_ (.S0(net10892),
    .A0(_02747_),
    .A1(_02748_),
    .A2(_02749_),
    .A3(_02750_),
    .S1(net10877),
    .X(_02751_));
 sg13g2_mux2_1 _20301_ (.A0(_02746_),
    .A1(_02751_),
    .S(net10880),
    .X(_02752_));
 sg13g2_a22oi_1 _20302_ (.Y(_02753_),
    .B1(_02752_),
    .B2(_11988_),
    .A2(net10317),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[23] ));
 sg13g2_nor2_1 _20303_ (.A(net10269),
    .B(_02753_),
    .Y(_02754_));
 sg13g2_a21oi_1 _20304_ (.A1(net10707),
    .A2(_02741_),
    .Y(_02755_),
    .B1(_02754_));
 sg13g2_nor2_1 _20305_ (.A(net9668),
    .B(_02755_),
    .Y(_02756_));
 sg13g2_a21oi_1 _20306_ (.A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[23] ),
    .A2(net9669),
    .Y(_02757_),
    .B1(_02756_));
 sg13g2_nand3_1 _20307_ (.B(_02733_),
    .C(_02757_),
    .A(_02732_),
    .Y(_01910_));
 sg13g2_inv_2 _20308_ (.Y(_02758_),
    .A(_00077_));
 sg13g2_nor2_1 _20309_ (.A(_00074_),
    .B(net10329),
    .Y(_02759_));
 sg13g2_a21oi_1 _20310_ (.A1(_02758_),
    .A2(net10329),
    .Y(_02760_),
    .B1(_02759_));
 sg13g2_nand2_1 _20311_ (.Y(_02761_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[28] ),
    .B(net10443));
 sg13g2_o21ai_1 _20312_ (.B1(_02761_),
    .Y(_02762_),
    .A1(_00082_),
    .A2(net10439));
 sg13g2_a22oi_1 _20313_ (.Y(_02763_),
    .B1(_02739_),
    .B2(_02762_),
    .A2(_02665_),
    .A1(net10329));
 sg13g2_o21ai_1 _20314_ (.B1(_02763_),
    .Y(_02764_),
    .A1(_08314_),
    .A2(_02760_));
 sg13g2_nor2_1 _20315_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[23] ),
    .B(net10557),
    .Y(_02765_));
 sg13g2_and2_1 _20316_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[23] ),
    .B(net10557),
    .X(_02766_));
 sg13g2_buf_2 place10342 (.A(net10341),
    .X(net10342));
 sg13g2_nor2_1 _20318_ (.A(net10682),
    .B(net10560),
    .Y(_02768_));
 sg13g2_and2_1 _20319_ (.A(net10682),
    .B(net10560),
    .X(_02769_));
 sg13g2_nor4_1 _20320_ (.A(_02765_),
    .B(_02766_),
    .C(_02768_),
    .D(_02769_),
    .Y(_02770_));
 sg13g2_nor2_1 _20321_ (.A(net10685),
    .B(net10566),
    .Y(_02771_));
 sg13g2_nor2_1 _20322_ (.A(net10684),
    .B(net10562),
    .Y(_02772_));
 sg13g2_nor4_1 _20323_ (.A(_02771_),
    .B(_02692_),
    .C(_02772_),
    .D(_02690_),
    .Y(_02773_));
 sg13g2_nand2_1 _20324_ (.Y(_02774_),
    .A(_02770_),
    .B(_02773_));
 sg13g2_a221oi_1 _20325_ (.B2(_02690_),
    .C1(_02692_),
    .B1(_02689_),
    .A1(net10682),
    .Y(_02775_),
    .A2(net10560));
 sg13g2_buf_2 place10304 (.A(_07193_),
    .X(net10304));
 sg13g2_or2_1 _20327_ (.X(_02777_),
    .B(_02768_),
    .A(_02765_));
 sg13g2_buf_2 place10390 (.A(net10389),
    .X(net10390));
 sg13g2_nor2_1 _20329_ (.A(_02775_),
    .B(_02777_),
    .Y(_02779_));
 sg13g2_nor2_1 _20330_ (.A(_02766_),
    .B(_02779_),
    .Y(_02780_));
 sg13g2_o21ai_1 _20331_ (.B1(_02780_),
    .Y(_02781_),
    .A1(_02619_),
    .A2(_02774_));
 sg13g2_xor2_1 _20332_ (.B(_02781_),
    .A(net10681),
    .X(_02782_));
 sg13g2_nor2_1 _20333_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[24] ),
    .B(net10338),
    .Y(_02783_));
 sg13g2_mux4_1 _20334_ (.S0(net10938),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][24] ),
    .S1(net10922),
    .X(_02784_));
 sg13g2_mux4_1 _20335_ (.S0(net10938),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][24] ),
    .S1(net10922),
    .X(_02785_));
 sg13g2_mux4_1 _20336_ (.S0(net10938),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][24] ),
    .S1(net10922),
    .X(_02786_));
 sg13g2_mux4_1 _20337_ (.S0(net10938),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][24] ),
    .S1(net10922),
    .X(_02787_));
 sg13g2_mux4_1 _20338_ (.S0(net10892),
    .A0(_02784_),
    .A1(_02785_),
    .A2(_02786_),
    .A3(_02787_),
    .S1(net10877),
    .X(_02788_));
 sg13g2_mux4_1 _20339_ (.S0(net10951),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][24] ),
    .S1(net10913),
    .X(_02789_));
 sg13g2_mux4_1 _20340_ (.S0(net10951),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][24] ),
    .S1(net10913),
    .X(_02790_));
 sg13g2_mux4_1 _20341_ (.S0(net10951),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][24] ),
    .S1(net10913),
    .X(_02791_));
 sg13g2_mux4_1 _20342_ (.S0(net10951),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][24] ),
    .S1(net10913),
    .X(_02792_));
 sg13g2_mux4_1 _20343_ (.S0(net10892),
    .A0(_02789_),
    .A1(_02790_),
    .A2(_02791_),
    .A3(_02792_),
    .S1(net10877),
    .X(_02793_));
 sg13g2_mux2_1 _20344_ (.A0(_02788_),
    .A1(_02793_),
    .S(net10880),
    .X(_02794_));
 sg13g2_a22oi_1 _20345_ (.Y(_02795_),
    .B1(_02794_),
    .B2(_11988_),
    .A2(net10317),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[24] ));
 sg13g2_nor2_1 _20346_ (.A(net10269),
    .B(_02795_),
    .Y(_02796_));
 sg13g2_a221oi_1 _20347_ (.B2(_02783_),
    .C1(_02796_),
    .B1(_02782_),
    .A1(net10707),
    .Y(_02797_),
    .A2(_02764_));
 sg13g2_nor2_1 _20348_ (.A(net10338),
    .B(_02782_),
    .Y(_02798_));
 sg13g2_o21ai_1 _20349_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[24] ),
    .Y(_02799_),
    .A1(net9669),
    .A2(_02798_));
 sg13g2_o21ai_1 _20350_ (.B1(_02799_),
    .Y(_01911_),
    .A1(net9669),
    .A2(_02797_));
 sg13g2_nand2_1 _20351_ (.Y(_02800_),
    .A(net10680),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[25] ));
 sg13g2_nor2_1 _20352_ (.A(net10338),
    .B(_02800_),
    .Y(_02801_));
 sg13g2_o21ai_1 _20353_ (.B1(_02781_),
    .Y(_02802_),
    .A1(net10681),
    .A2(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[24] ));
 sg13g2_nor4_1 _20354_ (.A(net10680),
    .B(net10551),
    .C(net10338),
    .D(net9669),
    .Y(_02803_));
 sg13g2_nor3_1 _20355_ (.A(_02801_),
    .B(_02802_),
    .C(_02803_),
    .Y(_02804_));
 sg13g2_and2_1 _20356_ (.A(net10681),
    .B(net10554),
    .X(_02805_));
 sg13g2_buf_2 place10255 (.A(net10254),
    .X(net10255));
 sg13g2_or4_1 _20358_ (.A(net10680),
    .B(_08610_),
    .C(net10338),
    .D(_02805_),
    .X(_02807_));
 sg13g2_nand2_2 _20359_ (.Y(_02808_),
    .A(net10681),
    .B(net10554));
 sg13g2_nand3_1 _20360_ (.B(net10294),
    .C(_02808_),
    .A(net10680),
    .Y(_02809_));
 sg13g2_or3_1 _20361_ (.A(net10551),
    .B(net9669),
    .C(_02809_),
    .X(_02810_));
 sg13g2_and3_1 _20362_ (.X(_02811_),
    .A(_02802_),
    .B(_02807_),
    .C(_02810_));
 sg13g2_nor4_1 _20363_ (.A(net10680),
    .B(net10551),
    .C(net10338),
    .D(_02808_),
    .Y(_02812_));
 sg13g2_inv_1 _20364_ (.Y(_02813_),
    .A(_00083_));
 sg13g2_a22oi_1 _20365_ (.Y(_02814_),
    .B1(net10332),
    .B2(_02813_),
    .A2(net10443),
    .A1(net10541));
 sg13g2_o21ai_1 _20366_ (.B1(_02814_),
    .Y(_02815_),
    .A1(_00075_),
    .A2(_08314_));
 sg13g2_nand2b_1 _20367_ (.Y(_02816_),
    .B(net10264),
    .A_N(_00078_));
 sg13g2_nand3_1 _20368_ (.B(_02707_),
    .C(_02816_),
    .A(net10326),
    .Y(_02817_));
 sg13g2_o21ai_1 _20369_ (.B1(_02817_),
    .Y(_02818_),
    .A1(net10329),
    .A2(_02815_));
 sg13g2_nor2_1 _20370_ (.A(net10392),
    .B(_02818_),
    .Y(_02819_));
 sg13g2_mux4_1 _20371_ (.S0(net10949),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][25] ),
    .S1(net10933),
    .X(_02820_));
 sg13g2_mux4_1 _20372_ (.S0(net10948),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][25] ),
    .S1(net10934),
    .X(_02821_));
 sg13g2_mux4_1 _20373_ (.S0(net10948),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][25] ),
    .S1(net10934),
    .X(_02822_));
 sg13g2_mux4_1 _20374_ (.S0(net10949),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][25] ),
    .S1(net10933),
    .X(_02823_));
 sg13g2_mux4_1 _20375_ (.S0(net10884),
    .A0(_02820_),
    .A1(_02821_),
    .A2(_02822_),
    .A3(_02823_),
    .S1(net10871),
    .X(_02824_));
 sg13g2_mux4_1 _20376_ (.S0(net10939),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][25] ),
    .S1(net10924),
    .X(_02825_));
 sg13g2_mux4_1 _20377_ (.S0(net10939),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][25] ),
    .S1(net10924),
    .X(_02826_));
 sg13g2_mux4_1 _20378_ (.S0(net10944),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][25] ),
    .S1(net10929),
    .X(_02827_));
 sg13g2_mux4_1 _20379_ (.S0(net10939),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][25] ),
    .S1(net10924),
    .X(_02828_));
 sg13g2_mux4_1 _20380_ (.S0(net10883),
    .A0(_02825_),
    .A1(_02826_),
    .A2(_02827_),
    .A3(_02828_),
    .S1(net10871),
    .X(_02829_));
 sg13g2_mux2_1 _20381_ (.A0(_02824_),
    .A1(_02829_),
    .S(net10879),
    .X(_02830_));
 sg13g2_a22oi_1 _20382_ (.Y(_02831_),
    .B1(_02830_),
    .B2(net10265),
    .A2(net10318),
    .A1(net10493));
 sg13g2_nor2_1 _20383_ (.A(net10270),
    .B(_02831_),
    .Y(_02832_));
 sg13g2_nor3_1 _20384_ (.A(_02812_),
    .B(_02819_),
    .C(_02832_),
    .Y(_02833_));
 sg13g2_nor2_1 _20385_ (.A(net9669),
    .B(_02833_),
    .Y(_02834_));
 sg13g2_a221oi_1 _20386_ (.B2(_02801_),
    .C1(_02834_),
    .B1(_02805_),
    .A1(net10551),
    .Y(_02835_),
    .A2(net9669));
 sg13g2_o21ai_1 _20387_ (.B1(_02835_),
    .Y(_01912_),
    .A1(_02804_),
    .A2(_02811_));
 sg13g2_inv_1 _20388_ (.Y(_02836_),
    .A(_00079_));
 sg13g2_mux4_1 _20389_ (.S0(net10264),
    .A0(net10536),
    .A1(_02734_),
    .A2(_02738_),
    .A3(_02836_),
    .S1(net10330),
    .X(_02837_));
 sg13g2_inv_1 _20390_ (.Y(_02838_),
    .A(net10679));
 sg13g2_and2_1 _20391_ (.A(net10680),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[25] ),
    .X(_02839_));
 sg13g2_buf_2 place10218 (.A(_10072_),
    .X(net10218));
 sg13g2_nor2_1 _20393_ (.A(net10681),
    .B(net10554),
    .Y(_02841_));
 sg13g2_nor2_1 _20394_ (.A(net10680),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[25] ),
    .Y(_02842_));
 sg13g2_nor4_1 _20395_ (.A(_02805_),
    .B(_02839_),
    .C(_02841_),
    .D(_02842_),
    .Y(_02843_));
 sg13g2_and2_1 _20396_ (.A(_02770_),
    .B(_02843_),
    .X(_02844_));
 sg13g2_buf_2 place10226 (.A(_09954_),
    .X(net10226));
 sg13g2_inv_1 _20398_ (.Y(_02846_),
    .A(_02844_));
 sg13g2_a21oi_1 _20399_ (.A1(net10682),
    .A2(net10560),
    .Y(_02847_),
    .B1(_02766_));
 sg13g2_nor3_1 _20400_ (.A(_02765_),
    .B(_02841_),
    .C(_02847_),
    .Y(_02848_));
 sg13g2_nand2b_1 _20401_ (.Y(_02849_),
    .B(_02808_),
    .A_N(_02848_));
 sg13g2_a21oi_1 _20402_ (.A1(net10552),
    .A2(_02849_),
    .Y(_02850_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[25] ));
 sg13g2_nor2_1 _20403_ (.A(net10552),
    .B(_02849_),
    .Y(_02851_));
 sg13g2_nor2_2 _20404_ (.A(_02850_),
    .B(_02851_),
    .Y(_02852_));
 sg13g2_inv_1 _20405_ (.Y(_02853_),
    .A(_02852_));
 sg13g2_o21ai_1 _20406_ (.B1(_02853_),
    .Y(_02854_),
    .A1(_02701_),
    .A2(_02846_));
 sg13g2_xnor2_1 _20407_ (.Y(_02855_),
    .A(_02838_),
    .B(_02854_));
 sg13g2_nor2_1 _20408_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[26] ),
    .B(net10337),
    .Y(_02856_));
 sg13g2_mux4_1 _20409_ (.S0(net10942),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][26] ),
    .S1(net10927),
    .X(_02857_));
 sg13g2_mux4_1 _20410_ (.S0(net10944),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][26] ),
    .S1(net10929),
    .X(_02858_));
 sg13g2_mux4_1 _20411_ (.S0(net10944),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][26] ),
    .S1(net10929),
    .X(_02859_));
 sg13g2_mux4_1 _20412_ (.S0(net10942),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][26] ),
    .S1(net10927),
    .X(_02860_));
 sg13g2_mux4_1 _20413_ (.S0(net10883),
    .A0(_02857_),
    .A1(_02858_),
    .A2(_02859_),
    .A3(_02860_),
    .S1(net10870),
    .X(_02861_));
 sg13g2_mux4_1 _20414_ (.S0(net10944),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][26] ),
    .S1(net10929),
    .X(_02862_));
 sg13g2_mux4_1 _20415_ (.S0(net10943),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][26] ),
    .S1(net10928),
    .X(_02863_));
 sg13g2_mux4_1 _20416_ (.S0(net10946),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][26] ),
    .S1(net10931),
    .X(_02864_));
 sg13g2_mux4_1 _20417_ (.S0(net10946),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][26] ),
    .S1(net10931),
    .X(_02865_));
 sg13g2_mux4_1 _20418_ (.S0(net10883),
    .A0(_02862_),
    .A1(_02863_),
    .A2(_02864_),
    .A3(_02865_),
    .S1(net10870),
    .X(_02866_));
 sg13g2_mux2_1 _20419_ (.A0(_02861_),
    .A1(_02866_),
    .S(net10878),
    .X(_02867_));
 sg13g2_a22oi_1 _20420_ (.Y(_02868_),
    .B1(_02867_),
    .B2(net10265),
    .A2(net10318),
    .A1(net10492));
 sg13g2_nor2_1 _20421_ (.A(net10270),
    .B(_02868_),
    .Y(_02869_));
 sg13g2_a221oi_1 _20422_ (.B2(_02856_),
    .C1(_02869_),
    .B1(_02855_),
    .A1(net10707),
    .Y(_02870_),
    .A2(_02837_));
 sg13g2_nor2_1 _20423_ (.A(net10337),
    .B(_02855_),
    .Y(_02871_));
 sg13g2_o21ai_1 _20424_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[26] ),
    .Y(_02872_),
    .A1(net9665),
    .A2(_02871_));
 sg13g2_o21ai_1 _20425_ (.B1(_02872_),
    .Y(_01913_),
    .A1(net9665),
    .A2(_02870_));
 sg13g2_nand3_1 _20426_ (.B(net10562),
    .C(_02844_),
    .A(net10548),
    .Y(_02873_));
 sg13g2_nand3_1 _20427_ (.B(net10548),
    .C(_02844_),
    .A(net10683),
    .Y(_02874_));
 sg13g2_nand3_1 _20428_ (.B(_02655_),
    .C(_02656_),
    .A(_02652_),
    .Y(_02875_));
 sg13g2_a221oi_1 _20429_ (.B2(_02874_),
    .C1(_02875_),
    .B1(_02873_),
    .A1(_02650_),
    .Y(_02876_),
    .A2(_02619_));
 sg13g2_nand4_1 _20430_ (.B(net10548),
    .C(net10562),
    .A(net10683),
    .Y(_02877_),
    .D(_02844_));
 sg13g2_o21ai_1 _20431_ (.B1(_02877_),
    .Y(_02878_),
    .A1(_08605_),
    .A2(_02853_));
 sg13g2_or2_1 _20432_ (.X(_02879_),
    .B(_02878_),
    .A(_02876_));
 sg13g2_or2_1 _20433_ (.X(_02880_),
    .B(net10563),
    .A(net10548));
 sg13g2_or2_1 _20434_ (.X(_02881_),
    .B(net10548),
    .A(net10683));
 sg13g2_a221oi_1 _20435_ (.B2(_02881_),
    .C1(_02852_),
    .B1(_02880_),
    .A1(_02651_),
    .Y(_02882_),
    .A2(_02657_));
 sg13g2_nand2_1 _20436_ (.Y(_02883_),
    .A(_08605_),
    .B(_02846_));
 sg13g2_or2_1 _20437_ (.X(_02884_),
    .B(_02881_),
    .A(net10562));
 sg13g2_a21oi_1 _20438_ (.A1(_02883_),
    .A2(_02884_),
    .Y(_02885_),
    .B1(_02852_));
 sg13g2_or3_1 _20439_ (.A(_02838_),
    .B(_02882_),
    .C(_02885_),
    .X(_02886_));
 sg13g2_nor2b_1 _20440_ (.A(_02879_),
    .B_N(_02886_),
    .Y(_02887_));
 sg13g2_xor2_1 _20441_ (.B(_02887_),
    .A(net10678),
    .X(_02888_));
 sg13g2_nor4_1 _20442_ (.A(net10546),
    .B(net10339),
    .C(net9670),
    .D(_02888_),
    .Y(_02889_));
 sg13g2_nand3_1 _20443_ (.B(net10294),
    .C(_02888_),
    .A(net10546),
    .Y(_02890_));
 sg13g2_mux4_1 _20444_ (.S0(net10264),
    .A0(net10533),
    .A1(_02758_),
    .A2(_02762_),
    .A3(_02706_),
    .S1(net10330),
    .X(_02891_));
 sg13g2_mux4_1 _20445_ (.S0(net10945),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][27] ),
    .S1(net10930),
    .X(_02892_));
 sg13g2_mux4_1 _20446_ (.S0(net10945),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][27] ),
    .S1(net10930),
    .X(_02893_));
 sg13g2_mux4_1 _20447_ (.S0(net10945),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][27] ),
    .S1(net10930),
    .X(_02894_));
 sg13g2_mux4_1 _20448_ (.S0(net10945),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][27] ),
    .S1(net10930),
    .X(_02895_));
 sg13g2_mux4_1 _20449_ (.S0(net10883),
    .A0(_02892_),
    .A1(_02893_),
    .A2(_02894_),
    .A3(_02895_),
    .S1(net10871),
    .X(_02896_));
 sg13g2_mux4_1 _20450_ (.S0(net10945),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][27] ),
    .S1(net10930),
    .X(_02897_));
 sg13g2_mux4_1 _20451_ (.S0(net10944),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][27] ),
    .S1(net10929),
    .X(_02898_));
 sg13g2_mux4_1 _20452_ (.S0(net10946),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][27] ),
    .S1(net10930),
    .X(_02899_));
 sg13g2_mux4_1 _20453_ (.S0(net10946),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][27] ),
    .S1(net10931),
    .X(_02900_));
 sg13g2_mux4_1 _20454_ (.S0(net10883),
    .A0(_02897_),
    .A1(_02898_),
    .A2(_02899_),
    .A3(_02900_),
    .S1(net10871),
    .X(_02901_));
 sg13g2_mux2_1 _20455_ (.A0(_02896_),
    .A1(_02901_),
    .S(net10879),
    .X(_02902_));
 sg13g2_a22oi_1 _20456_ (.Y(_02903_),
    .B1(_02902_),
    .B2(_11988_),
    .A2(net10318),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[27] ));
 sg13g2_nor2_1 _20457_ (.A(net10270),
    .B(_02903_),
    .Y(_02904_));
 sg13g2_a21oi_1 _20458_ (.A1(net10707),
    .A2(_02891_),
    .Y(_02905_),
    .B1(_02904_));
 sg13g2_mux2_1 _20459_ (.A0(_02905_),
    .A1(_08798_),
    .S(net9670),
    .X(_02906_));
 sg13g2_nand3b_1 _20460_ (.B(_02890_),
    .C(_02906_),
    .Y(_01914_),
    .A_N(_02889_));
 sg13g2_nor2_1 _20461_ (.A(_08586_),
    .B(net10439),
    .Y(_02907_));
 sg13g2_nor2_1 _20462_ (.A(net10330),
    .B(_02907_),
    .Y(_02908_));
 sg13g2_nor2_1 _20463_ (.A(_00081_),
    .B(_08314_),
    .Y(_02909_));
 sg13g2_nor2b_1 _20464_ (.A(_02909_),
    .B_N(_02814_),
    .Y(_02910_));
 sg13g2_a22oi_1 _20465_ (.Y(_02911_),
    .B1(_02910_),
    .B2(net10330),
    .A2(_02908_),
    .A1(_02816_));
 sg13g2_xnor2_1 _20466_ (.Y(_02912_),
    .A(net10679),
    .B(net10548));
 sg13g2_xnor2_1 _20467_ (.Y(_02913_),
    .A(net10678),
    .B(net10546));
 sg13g2_nor2_1 _20468_ (.A(net10686),
    .B(net10573),
    .Y(_02914_));
 sg13g2_nor3_1 _20469_ (.A(_02912_),
    .B(_02913_),
    .C(_02914_),
    .Y(_02915_));
 sg13g2_and3_2 _20470_ (.X(_02916_),
    .A(_02773_),
    .B(_02844_),
    .C(_02915_));
 sg13g2_o21ai_1 _20471_ (.B1(_02916_),
    .Y(_02917_),
    .A1(_02565_),
    .A2(_02567_));
 sg13g2_buf_2 place10239 (.A(net10235),
    .X(net10239));
 sg13g2_nor3_1 _20473_ (.A(net10554),
    .B(_02766_),
    .C(_02839_),
    .Y(_02919_));
 sg13g2_o21ai_1 _20474_ (.B1(_02919_),
    .Y(_02920_),
    .A1(_02775_),
    .A2(_02777_));
 sg13g2_nor3_1 _20475_ (.A(net10681),
    .B(_02766_),
    .C(_02839_),
    .Y(_02921_));
 sg13g2_o21ai_1 _20476_ (.B1(_02921_),
    .Y(_02922_),
    .A1(_02775_),
    .A2(_02777_));
 sg13g2_a21oi_1 _20477_ (.A1(_02800_),
    .A2(_02841_),
    .Y(_02923_),
    .B1(_02842_));
 sg13g2_and3_1 _20478_ (.X(_02924_),
    .A(_02920_),
    .B(_02922_),
    .C(_02923_));
 sg13g2_a21oi_1 _20479_ (.A1(net10549),
    .A2(_02924_),
    .Y(_02925_),
    .B1(net10679));
 sg13g2_nor2_1 _20480_ (.A(net10549),
    .B(_02924_),
    .Y(_02926_));
 sg13g2_nand2_1 _20481_ (.Y(_02927_),
    .A(net10678),
    .B(net10546));
 sg13g2_o21ai_1 _20482_ (.B1(_02927_),
    .Y(_02928_),
    .A1(_02925_),
    .A2(_02926_));
 sg13g2_or2_1 _20483_ (.X(_02929_),
    .B(net10546),
    .A(net10678));
 sg13g2_a21o_2 _20484_ (.A2(net10573),
    .A1(net10686),
    .B1(_02556_),
    .X(_02930_));
 sg13g2_a22oi_1 _20485_ (.Y(_02931_),
    .B1(_02916_),
    .B2(_02930_),
    .A2(_02929_),
    .A1(_02928_));
 sg13g2_buf_2 place10215 (.A(_11625_),
    .X(net10215));
 sg13g2_nand2_1 _20487_ (.Y(_02933_),
    .A(_02917_),
    .B(_02931_));
 sg13g2_xor2_1 _20488_ (.B(_02933_),
    .A(net10677),
    .X(_02934_));
 sg13g2_nor2_1 _20489_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[28] ),
    .B(net10339),
    .Y(_02935_));
 sg13g2_mux4_1 _20490_ (.S0(net10943),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][28] ),
    .S1(net10928),
    .X(_02936_));
 sg13g2_mux4_1 _20491_ (.S0(net10943),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][28] ),
    .S1(net10928),
    .X(_02937_));
 sg13g2_mux4_1 _20492_ (.S0(net10943),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][28] ),
    .S1(net10928),
    .X(_02938_));
 sg13g2_mux4_1 _20493_ (.S0(net10942),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][28] ),
    .S1(net10927),
    .X(_02939_));
 sg13g2_mux4_1 _20494_ (.S0(net10883),
    .A0(_02936_),
    .A1(_02937_),
    .A2(_02938_),
    .A3(_02939_),
    .S1(net10870),
    .X(_02940_));
 sg13g2_mux4_1 _20495_ (.S0(net10943),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][28] ),
    .S1(net10928),
    .X(_02941_));
 sg13g2_mux4_1 _20496_ (.S0(net10943),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][28] ),
    .S1(net10928),
    .X(_02942_));
 sg13g2_mux4_1 _20497_ (.S0(net10943),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][28] ),
    .S1(net10928),
    .X(_02943_));
 sg13g2_mux4_1 _20498_ (.S0(net10946),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][28] ),
    .S1(net10931),
    .X(_02944_));
 sg13g2_mux4_1 _20499_ (.S0(net10883),
    .A0(_02941_),
    .A1(_02942_),
    .A2(_02943_),
    .A3(_02944_),
    .S1(net10870),
    .X(_02945_));
 sg13g2_mux2_1 _20500_ (.A0(_02940_),
    .A1(_02945_),
    .S(net10878),
    .X(_02946_));
 sg13g2_a22oi_1 _20501_ (.Y(_02947_),
    .B1(_02946_),
    .B2(net10265),
    .A2(net10318),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[28] ));
 sg13g2_nor2_1 _20502_ (.A(net10270),
    .B(_02947_),
    .Y(_02948_));
 sg13g2_a221oi_1 _20503_ (.B2(_02935_),
    .C1(_02948_),
    .B1(_02934_),
    .A1(net10707),
    .Y(_02949_),
    .A2(_02911_));
 sg13g2_nor2_1 _20504_ (.A(net10339),
    .B(_02934_),
    .Y(_02950_));
 sg13g2_o21ai_1 _20505_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[28] ),
    .Y(_02951_),
    .A1(net9670),
    .A2(_02950_));
 sg13g2_o21ai_1 _20506_ (.B1(_02951_),
    .Y(_01915_),
    .A1(net9670),
    .A2(_02949_));
 sg13g2_inv_2 _20507_ (.Y(_02952_),
    .A(net10544));
 sg13g2_nand3_1 _20508_ (.B(_02917_),
    .C(_02931_),
    .A(_02952_),
    .Y(_02953_));
 sg13g2_a21oi_1 _20509_ (.A1(_02917_),
    .A2(_02931_),
    .Y(_02954_),
    .B1(_02952_));
 sg13g2_a21o_1 _20510_ (.A2(_02953_),
    .A1(net10677),
    .B1(_02954_),
    .X(_02955_));
 sg13g2_xor2_1 _20511_ (.B(_02955_),
    .A(net10676),
    .X(_02956_));
 sg13g2_nor2_1 _20512_ (.A(net10541),
    .B(net10339),
    .Y(_02957_));
 sg13g2_nor2_1 _20513_ (.A(_00082_),
    .B(net10409),
    .Y(_02958_));
 sg13g2_a21oi_1 _20514_ (.A1(_02836_),
    .A2(net10409),
    .Y(_02959_),
    .B1(_02958_));
 sg13g2_nor2_2 _20515_ (.A(_02336_),
    .B(net10406),
    .Y(_02960_));
 sg13g2_a22oi_1 _20516_ (.Y(_02961_),
    .B1(_02960_),
    .B2(net10536),
    .A2(_02907_),
    .A1(net10409));
 sg13g2_o21ai_1 _20517_ (.B1(_02961_),
    .Y(_02962_),
    .A1(_08314_),
    .A2(_02959_));
 sg13g2_mux4_1 _20518_ (.S0(net10949),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][29] ),
    .S1(net10933),
    .X(_02963_));
 sg13g2_mux4_1 _20519_ (.S0(net10948),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][29] ),
    .S1(net10934),
    .X(_02964_));
 sg13g2_mux4_1 _20520_ (.S0(net10948),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][29] ),
    .S1(net10934),
    .X(_02965_));
 sg13g2_mux4_1 _20521_ (.S0(net10949),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][29] ),
    .S1(net10933),
    .X(_02966_));
 sg13g2_mux4_1 _20522_ (.S0(net10884),
    .A0(_02963_),
    .A1(_02964_),
    .A2(_02965_),
    .A3(_02966_),
    .S1(net10871),
    .X(_02967_));
 sg13g2_mux4_1 _20523_ (.S0(net10948),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][29] ),
    .S1(net10934),
    .X(_02968_));
 sg13g2_mux4_1 _20524_ (.S0(net10948),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][29] ),
    .S1(net10934),
    .X(_02969_));
 sg13g2_mux4_1 _20525_ (.S0(net10948),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][29] ),
    .S1(net10934),
    .X(_02970_));
 sg13g2_mux4_1 _20526_ (.S0(net10949),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][29] ),
    .S1(net10933),
    .X(_02971_));
 sg13g2_mux4_1 _20527_ (.S0(net10884),
    .A0(_02968_),
    .A1(_02969_),
    .A2(_02970_),
    .A3(_02971_),
    .S1(net10871),
    .X(_02972_));
 sg13g2_mux2_1 _20528_ (.A0(_02967_),
    .A1(_02972_),
    .S(net10879),
    .X(_02973_));
 sg13g2_a22oi_1 _20529_ (.Y(_02974_),
    .B1(_02973_),
    .B2(net10265),
    .A2(net10318),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[29] ));
 sg13g2_nor2_1 _20530_ (.A(net10270),
    .B(_02974_),
    .Y(_02975_));
 sg13g2_a221oi_1 _20531_ (.B2(net10707),
    .C1(_02975_),
    .B1(_02962_),
    .A1(_02956_),
    .Y(_02976_),
    .A2(_02957_));
 sg13g2_nor2_1 _20532_ (.A(net10339),
    .B(_02956_),
    .Y(_02977_));
 sg13g2_o21ai_1 _20533_ (.B1(net10541),
    .Y(_02978_),
    .A1(net9670),
    .A2(_02977_));
 sg13g2_o21ai_1 _20534_ (.B1(_02978_),
    .Y(_01916_),
    .A1(net9670),
    .A2(_02976_));
 sg13g2_buf_2 place10198 (.A(_11808_),
    .X(net10198));
 sg13g2_buf_2 place10197 (.A(_03826_),
    .X(net10197));
 sg13g2_mux4_1 _20537_ (.S0(net10968),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][2] ),
    .S1(net10901),
    .X(_02981_));
 sg13g2_mux4_1 _20538_ (.S0(net10968),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][2] ),
    .S1(net10901),
    .X(_02982_));
 sg13g2_mux4_1 _20539_ (.S0(net10968),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][2] ),
    .S1(net10901),
    .X(_02983_));
 sg13g2_mux4_1 _20540_ (.S0(net10969),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][2] ),
    .S1(net10903),
    .X(_02984_));
 sg13g2_mux4_1 _20541_ (.S0(net10889),
    .A0(_02981_),
    .A1(_02982_),
    .A2(_02983_),
    .A3(_02984_),
    .S1(net10873),
    .X(_02985_));
 sg13g2_mux4_1 _20542_ (.S0(net10969),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][2] ),
    .S1(net10901),
    .X(_02986_));
 sg13g2_mux4_1 _20543_ (.S0(net10967),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][2] ),
    .S1(net10902),
    .X(_02987_));
 sg13g2_mux4_1 _20544_ (.S0(net10969),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][2] ),
    .S1(net10903),
    .X(_02988_));
 sg13g2_mux4_1 _20545_ (.S0(net10969),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][2] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][2] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][2] ),
    .S1(net10903),
    .X(_02989_));
 sg13g2_mux4_1 _20546_ (.S0(net10889),
    .A0(_02986_),
    .A1(_02987_),
    .A2(_02988_),
    .A3(_02989_),
    .S1(net10873),
    .X(_02990_));
 sg13g2_mux2_1 _20547_ (.A0(_02985_),
    .A1(_02990_),
    .S(net10882),
    .X(_02991_));
 sg13g2_a22oi_1 _20548_ (.Y(_02992_),
    .B1(_02991_),
    .B2(net10268),
    .A2(net10320),
    .A1(net10491));
 sg13g2_a22oi_1 _20549_ (.Y(_02993_),
    .B1(net10331),
    .B2(_12038_),
    .A2(net10442),
    .A1(net10526));
 sg13g2_inv_2 _20550_ (.Y(_02994_),
    .A(_00059_));
 sg13g2_a22oi_1 _20551_ (.Y(_02995_),
    .B1(net10331),
    .B2(_02994_),
    .A2(net10442),
    .A1(net10531));
 sg13g2_o21ai_1 _20552_ (.B1(_02995_),
    .Y(_02996_),
    .A1(_00053_),
    .A2(net10289));
 sg13g2_nand2_1 _20553_ (.Y(_02997_),
    .A(net10324),
    .B(_02996_));
 sg13g2_o21ai_1 _20554_ (.B1(_02997_),
    .Y(_02998_),
    .A1(net10324),
    .A2(_02993_));
 sg13g2_a21o_2 _20555_ (.A2(_12012_),
    .A1(net10572),
    .B1(_12015_),
    .X(_02999_));
 sg13g2_xnor2_1 _20556_ (.Y(_03000_),
    .A(net10675),
    .B(net10538));
 sg13g2_xnor2_1 _20557_ (.Y(_03001_),
    .A(_02999_),
    .B(_03000_));
 sg13g2_a22oi_1 _20558_ (.Y(_03002_),
    .B1(_03001_),
    .B2(net10293),
    .A2(_02998_),
    .A1(net10702));
 sg13g2_o21ai_1 _20559_ (.B1(_03002_),
    .Y(_03003_),
    .A1(net10272),
    .A2(_02992_));
 sg13g2_mux2_1 _20560_ (.A0(_03003_),
    .A1(net10538),
    .S(net9673),
    .X(_01917_));
 sg13g2_a21oi_1 _20561_ (.A1(net10443),
    .A2(net10330),
    .Y(_03004_),
    .B1(net10332));
 sg13g2_nand2_1 _20562_ (.Y(_03005_),
    .A(_00080_),
    .B(net10409));
 sg13g2_nand2_1 _20563_ (.Y(_03006_),
    .A(_00083_),
    .B(net10330));
 sg13g2_nand3_1 _20564_ (.B(_03005_),
    .C(_03006_),
    .A(net10264),
    .Y(_03007_));
 sg13g2_o21ai_1 _20565_ (.B1(_03007_),
    .Y(_03008_),
    .A1(_08586_),
    .A2(_03004_));
 sg13g2_or2_1 _20566_ (.X(_03009_),
    .B(net10541),
    .A(net10676));
 sg13g2_and2_1 _20567_ (.A(net10676),
    .B(net10541),
    .X(_03010_));
 sg13g2_buf_2 place10254 (.A(net10253),
    .X(net10254));
 sg13g2_a21oi_1 _20569_ (.A1(_02955_),
    .A2(_03009_),
    .Y(_03012_),
    .B1(_03010_));
 sg13g2_xnor2_1 _20570_ (.Y(_03013_),
    .A(net10674),
    .B(_03012_));
 sg13g2_nor2_1 _20571_ (.A(net10536),
    .B(net10339),
    .Y(_03014_));
 sg13g2_mux4_1 _20572_ (.S0(net10941),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][30] ),
    .S1(net10926),
    .X(_03015_));
 sg13g2_mux4_1 _20573_ (.S0(net10941),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][30] ),
    .S1(net10926),
    .X(_03016_));
 sg13g2_mux4_1 _20574_ (.S0(net10941),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][30] ),
    .S1(net10926),
    .X(_03017_));
 sg13g2_mux4_1 _20575_ (.S0(net10941),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][30] ),
    .S1(net10926),
    .X(_03018_));
 sg13g2_mux4_1 _20576_ (.S0(_00007_),
    .A0(_03015_),
    .A1(_03016_),
    .A2(_03017_),
    .A3(_03018_),
    .S1(net10869),
    .X(_03019_));
 sg13g2_mux4_1 _20577_ (.S0(net10939),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][30] ),
    .S1(net10924),
    .X(_03020_));
 sg13g2_mux4_1 _20578_ (.S0(net10941),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][30] ),
    .S1(net10926),
    .X(_03021_));
 sg13g2_mux4_1 _20579_ (.S0(net10941),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][30] ),
    .S1(net10926),
    .X(_03022_));
 sg13g2_mux4_1 _20580_ (.S0(net10941),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][30] ),
    .S1(net10926),
    .X(_03023_));
 sg13g2_mux4_1 _20581_ (.S0(_00007_),
    .A0(_03020_),
    .A1(_03021_),
    .A2(_03022_),
    .A3(_03023_),
    .S1(net10869),
    .X(_03024_));
 sg13g2_mux2_1 _20582_ (.A0(_03019_),
    .A1(_03024_),
    .S(net10878),
    .X(_03025_));
 sg13g2_a22oi_1 _20583_ (.Y(_03026_),
    .B1(_03025_),
    .B2(net10265),
    .A2(net10318),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[30] ));
 sg13g2_nor2_1 _20584_ (.A(net10270),
    .B(_03026_),
    .Y(_03027_));
 sg13g2_a221oi_1 _20585_ (.B2(_03014_),
    .C1(_03027_),
    .B1(_03013_),
    .A1(net10707),
    .Y(_03028_),
    .A2(_03008_));
 sg13g2_nor2_1 _20586_ (.A(net10339),
    .B(_03013_),
    .Y(_03029_));
 sg13g2_o21ai_1 _20587_ (.B1(net10536),
    .Y(_03030_),
    .A1(net9670),
    .A2(_03029_));
 sg13g2_o21ai_1 _20588_ (.B1(_03030_),
    .Y(_01918_),
    .A1(net9670),
    .A2(_03028_));
 sg13g2_nand2_1 _20589_ (.Y(_03031_),
    .A(_11948_),
    .B(_11937_));
 sg13g2_and2_1 _20590_ (.A(_11942_),
    .B(_03031_),
    .X(_03032_));
 sg13g2_o21ai_1 _20591_ (.B1(_03032_),
    .Y(_03033_),
    .A1(_11932_),
    .A2(_11935_));
 sg13g2_buf_2 place10196 (.A(_06688_),
    .X(net10196));
 sg13g2_nor2_1 _20593_ (.A(net10677),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[28] ),
    .Y(_03035_));
 sg13g2_nand2_1 _20594_ (.Y(_03036_),
    .A(net10677),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[28] ));
 sg13g2_o21ai_1 _20595_ (.B1(_03036_),
    .Y(_03037_),
    .A1(_02927_),
    .A2(_03035_));
 sg13g2_o21ai_1 _20596_ (.B1(_03009_),
    .Y(_03038_),
    .A1(_03010_),
    .A2(_03037_));
 sg13g2_nand2b_2 _20597_ (.Y(_03039_),
    .B(_03038_),
    .A_N(net10536));
 sg13g2_nor3_1 _20598_ (.A(_02876_),
    .B(_02878_),
    .C(_03039_),
    .Y(_03040_));
 sg13g2_nand3_1 _20599_ (.B(net10542),
    .C(net10544),
    .A(net10535),
    .Y(_03041_));
 sg13g2_nand3_1 _20600_ (.B(net10535),
    .C(net10544),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[29] ),
    .Y(_03042_));
 sg13g2_a22oi_1 _20601_ (.Y(_03043_),
    .B1(_03041_),
    .B2(_03042_),
    .A2(_02931_),
    .A1(_02917_));
 sg13g2_nand3_1 _20602_ (.B(net10535),
    .C(net10542),
    .A(net10677),
    .Y(_03044_));
 sg13g2_nand3_1 _20603_ (.B(net10676),
    .C(net10535),
    .A(net10677),
    .Y(_03045_));
 sg13g2_a22oi_1 _20604_ (.Y(_03046_),
    .B1(_03044_),
    .B2(_03045_),
    .A2(_02931_),
    .A1(_02917_));
 sg13g2_nand4_1 _20605_ (.B(net10535),
    .C(net10542),
    .A(net10677),
    .Y(_03047_),
    .D(net10544));
 sg13g2_nand4_1 _20606_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[29] ),
    .C(net10535),
    .A(net10677),
    .Y(_03048_),
    .D(net10544));
 sg13g2_nand3_1 _20607_ (.B(net10535),
    .C(net10542),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[29] ),
    .Y(_03049_));
 sg13g2_nand3_1 _20608_ (.B(_03048_),
    .C(_03049_),
    .A(_03047_),
    .Y(_03050_));
 sg13g2_nor4_1 _20609_ (.A(net10674),
    .B(_03043_),
    .C(_03046_),
    .D(_03050_),
    .Y(_03051_));
 sg13g2_nor2_1 _20610_ (.A(net10676),
    .B(net10541),
    .Y(_03052_));
 sg13g2_nand2b_1 _20611_ (.Y(_03053_),
    .B(_03036_),
    .A_N(_03035_));
 sg13g2_nor4_2 _20612_ (.A(_02913_),
    .B(_03010_),
    .C(_03052_),
    .Y(_03054_),
    .D(_03053_));
 sg13g2_nor2_1 _20613_ (.A(_03054_),
    .B(_03039_),
    .Y(_03055_));
 sg13g2_or2_1 _20614_ (.X(_03056_),
    .B(_03055_),
    .A(_03051_));
 sg13g2_a21oi_1 _20615_ (.A1(_02886_),
    .A2(_03040_),
    .Y(_03057_),
    .B1(_03056_));
 sg13g2_nor3_1 _20616_ (.A(net10533),
    .B(_03033_),
    .C(_03057_),
    .Y(_03058_));
 sg13g2_and2_1 _20617_ (.A(net10679),
    .B(_03054_),
    .X(_03059_));
 sg13g2_nor2_1 _20618_ (.A(_02882_),
    .B(_02885_),
    .Y(_03060_));
 sg13g2_a221oi_1 _20619_ (.B2(_03060_),
    .C1(_03039_),
    .B1(_03059_),
    .A1(_02879_),
    .Y(_03061_),
    .A2(_03054_));
 sg13g2_xnor2_1 _20620_ (.Y(_03062_),
    .A(_11497_),
    .B(_03061_));
 sg13g2_and2_1 _20621_ (.A(net10674),
    .B(net10533),
    .X(_03063_));
 sg13g2_or3_1 _20622_ (.A(_03043_),
    .B(_03046_),
    .C(_03050_),
    .X(_03064_));
 sg13g2_nor4_1 _20623_ (.A(net10674),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[31] ),
    .C(_08586_),
    .D(_03064_),
    .Y(_03065_));
 sg13g2_nand3_1 _20624_ (.B(net10533),
    .C(_03064_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[31] ),
    .Y(_03066_));
 sg13g2_nand2b_1 _20625_ (.Y(_03067_),
    .B(_03066_),
    .A_N(_03065_));
 sg13g2_a221oi_1 _20626_ (.B2(_03063_),
    .C1(_03067_),
    .B1(_03062_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[31] ),
    .Y(_03068_),
    .A2(_03058_));
 sg13g2_nand3_1 _20627_ (.B(_08586_),
    .C(net10294),
    .A(_11497_),
    .Y(_03069_));
 sg13g2_nor4_1 _20628_ (.A(_03033_),
    .B(_03069_),
    .C(_03061_),
    .D(_03051_),
    .Y(_03070_));
 sg13g2_mux4_1 _20629_ (.S0(net10940),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][31] ),
    .S1(net10925),
    .X(_03071_));
 sg13g2_mux4_1 _20630_ (.S0(net10940),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][31] ),
    .S1(net10925),
    .X(_03072_));
 sg13g2_mux4_1 _20631_ (.S0(net10940),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][31] ),
    .S1(net10925),
    .X(_03073_));
 sg13g2_mux4_1 _20632_ (.S0(net10940),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][31] ),
    .S1(net10925),
    .X(_03074_));
 sg13g2_mux4_1 _20633_ (.S0(_00007_),
    .A0(_03071_),
    .A1(_03072_),
    .A2(_03073_),
    .A3(_03074_),
    .S1(net10870),
    .X(_03075_));
 sg13g2_mux4_1 _20634_ (.S0(net10947),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][31] ),
    .S1(net10923),
    .X(_03076_));
 sg13g2_mux4_1 _20635_ (.S0(net10947),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][31] ),
    .S1(net10923),
    .X(_03077_));
 sg13g2_mux4_1 _20636_ (.S0(net10939),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][31] ),
    .S1(net10924),
    .X(_03078_));
 sg13g2_mux4_1 _20637_ (.S0(net10939),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][31] ),
    .S1(net10924),
    .X(_03079_));
 sg13g2_mux4_1 _20638_ (.S0(net10886),
    .A0(_03076_),
    .A1(_03077_),
    .A2(_03078_),
    .A3(_03079_),
    .S1(net10869),
    .X(_03080_));
 sg13g2_mux2_1 _20639_ (.A0(_03075_),
    .A1(_03080_),
    .S(net10878),
    .X(_03081_));
 sg13g2_a22oi_1 _20640_ (.Y(_03082_),
    .B1(_03081_),
    .B2(net10265),
    .A2(net10318),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[31] ));
 sg13g2_nand2_1 _20641_ (.Y(_03083_),
    .A(net10536),
    .B(net10330));
 sg13g2_o21ai_1 _20642_ (.B1(_03083_),
    .Y(_03084_),
    .A1(_08798_),
    .A2(net10330));
 sg13g2_nand3_1 _20643_ (.B(net10264),
    .C(_03084_),
    .A(net10707),
    .Y(_03085_));
 sg13g2_o21ai_1 _20644_ (.B1(_03085_),
    .Y(_03086_),
    .A1(net10270),
    .A2(_03082_));
 sg13g2_mux2_1 _20645_ (.A0(_03086_),
    .A1(net10533),
    .S(_03033_),
    .X(_03087_));
 sg13g2_nor2_1 _20646_ (.A(_03070_),
    .B(_03087_),
    .Y(_03088_));
 sg13g2_o21ai_1 _20647_ (.B1(_03088_),
    .Y(_01919_),
    .A1(net10339),
    .A2(_03068_));
 sg13g2_mux4_1 _20648_ (.S0(net10962),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][3] ),
    .S1(net10898),
    .X(_03089_));
 sg13g2_mux4_1 _20649_ (.S0(net10962),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][3] ),
    .S1(net10898),
    .X(_03090_));
 sg13g2_mux4_1 _20650_ (.S0(net10954),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][3] ),
    .S1(net10916),
    .X(_03091_));
 sg13g2_mux4_1 _20651_ (.S0(net10956),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][3] ),
    .S1(net10916),
    .X(_03092_));
 sg13g2_mux4_1 _20652_ (.S0(net10888),
    .A0(_03089_),
    .A1(_03090_),
    .A2(_03091_),
    .A3(_03092_),
    .S1(net10872),
    .X(_03093_));
 sg13g2_mux4_1 _20653_ (.S0(net10962),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][3] ),
    .S1(net10897),
    .X(_03094_));
 sg13g2_mux4_1 _20654_ (.S0(net10962),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][3] ),
    .S1(net10898),
    .X(_03095_));
 sg13g2_mux4_1 _20655_ (.S0(net10956),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][3] ),
    .S1(net10916),
    .X(_03096_));
 sg13g2_mux4_1 _20656_ (.S0(net10961),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][3] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][3] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][3] ),
    .S1(net10898),
    .X(_03097_));
 sg13g2_mux4_1 _20657_ (.S0(net10888),
    .A0(_03094_),
    .A1(_03095_),
    .A2(_03096_),
    .A3(_03097_),
    .S1(net10872),
    .X(_03098_));
 sg13g2_mux2_1 _20658_ (.A0(_03093_),
    .A1(_03098_),
    .S(net10882),
    .X(_03099_));
 sg13g2_a22oi_1 _20659_ (.Y(_03100_),
    .B1(_03099_),
    .B2(net10268),
    .A2(net10320),
    .A1(net10490));
 sg13g2_nand2_1 _20660_ (.Y(_03101_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[7] ),
    .B(net10442));
 sg13g2_o21ai_1 _20661_ (.B1(_03101_),
    .Y(_03102_),
    .A1(_00061_),
    .A2(net10438));
 sg13g2_o21ai_1 _20662_ (.B1(_11952_),
    .Y(_03103_),
    .A1(_00057_),
    .A2(net10289));
 sg13g2_mux2_1 _20663_ (.A0(_03102_),
    .A1(_03103_),
    .S(net10324),
    .X(_03104_));
 sg13g2_o21ai_1 _20664_ (.B1(_02999_),
    .Y(_03105_),
    .A1(net10675),
    .A2(net10538));
 sg13g2_nand2_1 _20665_ (.Y(_03106_),
    .A(net10675),
    .B(net10538));
 sg13g2_nand2_1 _20666_ (.Y(_03107_),
    .A(_03105_),
    .B(_03106_));
 sg13g2_xnor2_1 _20667_ (.Y(_03108_),
    .A(net10673),
    .B(net10531));
 sg13g2_xnor2_1 _20668_ (.Y(_03109_),
    .A(_03107_),
    .B(_03108_));
 sg13g2_a22oi_1 _20669_ (.Y(_03110_),
    .B1(_03109_),
    .B2(net10293),
    .A2(_03104_),
    .A1(net10702));
 sg13g2_o21ai_1 _20670_ (.B1(_03110_),
    .Y(_03111_),
    .A1(net10272),
    .A2(_03100_));
 sg13g2_mux2_1 _20671_ (.A0(_03111_),
    .A1(net10531),
    .S(net9673),
    .X(_01920_));
 sg13g2_mux4_1 _20672_ (.S0(net10956),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][4] ),
    .S1(net10917),
    .X(_03112_));
 sg13g2_mux4_1 _20673_ (.S0(net10956),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][4] ),
    .S1(net10917),
    .X(_03113_));
 sg13g2_mux4_1 _20674_ (.S0(net10956),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][4] ),
    .S1(net10917),
    .X(_03114_));
 sg13g2_mux4_1 _20675_ (.S0(net10956),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][4] ),
    .S1(net10917),
    .X(_03115_));
 sg13g2_mux4_1 _20676_ (.S0(net10887),
    .A0(_03112_),
    .A1(_03113_),
    .A2(_03114_),
    .A3(_03115_),
    .S1(net10876),
    .X(_03116_));
 sg13g2_mux4_1 _20677_ (.S0(net10955),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][4] ),
    .S1(net10917),
    .X(_03117_));
 sg13g2_mux4_1 _20678_ (.S0(net10955),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][4] ),
    .S1(net10917),
    .X(_03118_));
 sg13g2_mux4_1 _20679_ (.S0(net10955),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][4] ),
    .S1(net10917),
    .X(_03119_));
 sg13g2_mux4_1 _20680_ (.S0(net10955),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][4] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][4] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][4] ),
    .S1(net10917),
    .X(_03120_));
 sg13g2_mux4_1 _20681_ (.S0(net10887),
    .A0(_03117_),
    .A1(_03118_),
    .A2(_03119_),
    .A3(_03120_),
    .S1(net10876),
    .X(_03121_));
 sg13g2_mux2_1 _20682_ (.A0(_03116_),
    .A1(_03121_),
    .S(net10882),
    .X(_03122_));
 sg13g2_a22oi_1 _20683_ (.Y(_03123_),
    .B1(_03122_),
    .B2(net10268),
    .A2(net10320),
    .A1(net10489));
 sg13g2_nor2_1 _20684_ (.A(_00056_),
    .B(net10324),
    .Y(_03124_));
 sg13g2_a21oi_1 _20685_ (.A1(_02994_),
    .A2(net10324),
    .Y(_03125_),
    .B1(_03124_));
 sg13g2_nand2_1 _20686_ (.Y(_03126_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[8] ),
    .B(net10442));
 sg13g2_o21ai_1 _20687_ (.B1(_03126_),
    .Y(_03127_),
    .A1(_00062_),
    .A2(net10438));
 sg13g2_nand2_1 _20688_ (.Y(_03128_),
    .A(net10324),
    .B(_02598_));
 sg13g2_o21ai_1 _20689_ (.B1(_03128_),
    .Y(_03129_),
    .A1(net10323),
    .A2(_03127_));
 sg13g2_o21ai_1 _20690_ (.B1(_03129_),
    .Y(_03130_),
    .A1(net10289),
    .A2(_03125_));
 sg13g2_nor2_1 _20691_ (.A(_12016_),
    .B(_12021_),
    .Y(_03131_));
 sg13g2_xnor2_1 _20692_ (.Y(_03132_),
    .A(net10672),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[4] ));
 sg13g2_xnor2_1 _20693_ (.Y(_03133_),
    .A(_03131_),
    .B(_03132_));
 sg13g2_a22oi_1 _20694_ (.Y(_03134_),
    .B1(_03133_),
    .B2(net10293),
    .A2(_03130_),
    .A1(net10702));
 sg13g2_o21ai_1 _20695_ (.B1(_03134_),
    .Y(_03135_),
    .A1(net10272),
    .A2(_03123_));
 sg13g2_nor2_1 _20696_ (.A(net9673),
    .B(_03135_),
    .Y(_03136_));
 sg13g2_a21oi_1 _20697_ (.A1(_08701_),
    .A2(net9673),
    .Y(_01921_),
    .B1(_03136_));
 sg13g2_xnor2_1 _20698_ (.Y(_03137_),
    .A(net10671),
    .B(_12025_));
 sg13g2_nor2_1 _20699_ (.A(net10528),
    .B(net10334),
    .Y(_03138_));
 sg13g2_nor2_1 _20700_ (.A(_00055_),
    .B(net10413),
    .Y(_03139_));
 sg13g2_a21oi_1 _20701_ (.A1(_11955_),
    .A2(net10413),
    .Y(_03140_),
    .B1(_03139_));
 sg13g2_a22oi_1 _20702_ (.Y(_03141_),
    .B1(net10331),
    .B2(_02333_),
    .A2(net10441),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[9] ));
 sg13g2_mux2_1 _20703_ (.A0(_02993_),
    .A1(_03141_),
    .S(net10413),
    .X(_03142_));
 sg13g2_o21ai_1 _20704_ (.B1(_03142_),
    .Y(_03143_),
    .A1(net10289),
    .A2(_03140_));
 sg13g2_mux4_1 _20705_ (.S0(net10963),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][5] ),
    .S1(net10899),
    .X(_03144_));
 sg13g2_mux4_1 _20706_ (.S0(net10963),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][5] ),
    .S1(net10899),
    .X(_03145_));
 sg13g2_mux4_1 _20707_ (.S0(net10963),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][5] ),
    .S1(net10899),
    .X(_03146_));
 sg13g2_mux4_1 _20708_ (.S0(net10963),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][5] ),
    .S1(net10899),
    .X(_03147_));
 sg13g2_mux4_1 _20709_ (.S0(net10889),
    .A0(_03144_),
    .A1(_03145_),
    .A2(_03146_),
    .A3(_03147_),
    .S1(net10873),
    .X(_03148_));
 sg13g2_mux4_1 _20710_ (.S0(net10969),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][5] ),
    .S1(net10903),
    .X(_03149_));
 sg13g2_mux4_1 _20711_ (.S0(net10967),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][5] ),
    .S1(net10902),
    .X(_03150_));
 sg13g2_mux4_1 _20712_ (.S0(net10969),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][5] ),
    .S1(net10903),
    .X(_03151_));
 sg13g2_mux4_1 _20713_ (.S0(net10969),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][5] ),
    .S1(net10903),
    .X(_03152_));
 sg13g2_mux4_1 _20714_ (.S0(net10889),
    .A0(_03149_),
    .A1(_03150_),
    .A2(_03151_),
    .A3(_03152_),
    .S1(net10873),
    .X(_03153_));
 sg13g2_mux2_1 _20715_ (.A0(_03148_),
    .A1(_03153_),
    .S(net10882),
    .X(_03154_));
 sg13g2_a22oi_1 _20716_ (.Y(_03155_),
    .B1(_03154_),
    .B2(net10268),
    .A2(net10320),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[5] ));
 sg13g2_nor2_1 _20717_ (.A(net10272),
    .B(_03155_),
    .Y(_03156_));
 sg13g2_a221oi_1 _20718_ (.B2(net10701),
    .C1(_03156_),
    .B1(_03143_),
    .A1(_03137_),
    .Y(_03157_),
    .A2(_03138_));
 sg13g2_nor2_1 _20719_ (.A(net10334),
    .B(_03137_),
    .Y(_03158_));
 sg13g2_o21ai_1 _20720_ (.B1(net10528),
    .Y(_03159_),
    .A1(net9672),
    .A2(_03158_));
 sg13g2_o21ai_1 _20721_ (.B1(_03159_),
    .Y(_01922_),
    .A1(net9672),
    .A2(_03157_));
 sg13g2_nand2b_1 _20722_ (.Y(_03160_),
    .B(_12025_),
    .A_N(net10528));
 sg13g2_nor2b_1 _20723_ (.A(_12025_),
    .B_N(net10528),
    .Y(_03161_));
 sg13g2_a21o_2 _20724_ (.A2(_03160_),
    .A1(net10671),
    .B1(_03161_),
    .X(_03162_));
 sg13g2_buf_2 place10230 (.A(_07979_),
    .X(net10230));
 sg13g2_xnor2_1 _20726_ (.Y(_03164_),
    .A(net10670),
    .B(_03162_));
 sg13g2_nor2_1 _20727_ (.A(net10526),
    .B(_03164_),
    .Y(_03165_));
 sg13g2_nor2_1 _20728_ (.A(_00058_),
    .B(net10412),
    .Y(_03166_));
 sg13g2_a21oi_1 _20729_ (.A1(_02599_),
    .A2(net10410),
    .Y(_03167_),
    .B1(_03166_));
 sg13g2_nand2_1 _20730_ (.Y(_03168_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[10] ),
    .B(net10441));
 sg13g2_o21ai_1 _20731_ (.B1(_03168_),
    .Y(_03169_),
    .A1(_00064_),
    .A2(net10438));
 sg13g2_a22oi_1 _20732_ (.Y(_03170_),
    .B1(_03169_),
    .B2(net10411),
    .A2(_03102_),
    .A1(_02960_));
 sg13g2_o21ai_1 _20733_ (.B1(_03170_),
    .Y(_03171_),
    .A1(net10290),
    .A2(_03167_));
 sg13g2_mux4_1 _20734_ (.S0(net10970),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][6] ),
    .S1(net10908),
    .X(_03172_));
 sg13g2_mux4_1 _20735_ (.S0(net10970),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][6] ),
    .S1(net10908),
    .X(_03173_));
 sg13g2_mux4_1 _20736_ (.S0(net10972),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][6] ),
    .S1(net10906),
    .X(_03174_));
 sg13g2_mux4_1 _20737_ (.S0(net10972),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][6] ),
    .S1(net10906),
    .X(_03175_));
 sg13g2_mux4_1 _20738_ (.S0(net10891),
    .A0(_03172_),
    .A1(_03173_),
    .A2(_03174_),
    .A3(_03175_),
    .S1(net10875),
    .X(_03176_));
 sg13g2_mux4_1 _20739_ (.S0(net10972),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][6] ),
    .S1(net10908),
    .X(_03177_));
 sg13g2_mux4_1 _20740_ (.S0(net10972),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][6] ),
    .S1(net10908),
    .X(_03178_));
 sg13g2_mux4_1 _20741_ (.S0(net10972),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][6] ),
    .S1(net10908),
    .X(_03179_));
 sg13g2_mux4_1 _20742_ (.S0(net10974),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][6] ),
    .S1(net10905),
    .X(_03180_));
 sg13g2_mux4_1 _20743_ (.S0(net10891),
    .A0(_03177_),
    .A1(_03178_),
    .A2(_03179_),
    .A3(_03180_),
    .S1(net10875),
    .X(_03181_));
 sg13g2_mux2_1 _20744_ (.A0(_03176_),
    .A1(_03181_),
    .S(net10881),
    .X(_03182_));
 sg13g2_a22oi_1 _20745_ (.Y(_03183_),
    .B1(_03182_),
    .B2(net10268),
    .A2(net10320),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[6] ));
 sg13g2_nor2_1 _20746_ (.A(net10272),
    .B(_03183_),
    .Y(_03184_));
 sg13g2_a221oi_1 _20747_ (.B2(net10702),
    .C1(_03184_),
    .B1(_03171_),
    .A1(net10293),
    .Y(_03185_),
    .A2(_03165_));
 sg13g2_and2_1 _20748_ (.A(net10293),
    .B(_03164_),
    .X(_03186_));
 sg13g2_o21ai_1 _20749_ (.B1(net10526),
    .Y(_03187_),
    .A1(net9673),
    .A2(_03186_));
 sg13g2_o21ai_1 _20750_ (.B1(_03187_),
    .Y(_01923_),
    .A1(net9673),
    .A2(_03185_));
 sg13g2_a21o_1 _20751_ (.A2(_03162_),
    .A1(net10526),
    .B1(net10670),
    .X(_03188_));
 sg13g2_o21ai_1 _20752_ (.B1(_03188_),
    .Y(_03189_),
    .A1(net10526),
    .A2(_03162_));
 sg13g2_xnor2_1 _20753_ (.Y(_03190_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[7] ),
    .B(_03189_));
 sg13g2_nor2_1 _20754_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[7] ),
    .B(net10334),
    .Y(_03191_));
 sg13g2_nor2_1 _20755_ (.A(_00060_),
    .B(net10413),
    .Y(_03192_));
 sg13g2_a21oi_1 _20756_ (.A1(_02994_),
    .A2(net10410),
    .Y(_03193_),
    .B1(_03192_));
 sg13g2_nand2_1 _20757_ (.Y(_03194_),
    .A(net10412),
    .B(_02182_));
 sg13g2_o21ai_1 _20758_ (.B1(_03194_),
    .Y(_03195_),
    .A1(net10410),
    .A2(_03127_));
 sg13g2_o21ai_1 _20759_ (.B1(_03195_),
    .Y(_03196_),
    .A1(net10289),
    .A2(_03193_));
 sg13g2_mux4_1 _20760_ (.S0(net10967),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][7] ),
    .S1(net10902),
    .X(_03197_));
 sg13g2_mux4_1 _20761_ (.S0(net10970),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][7] ),
    .S1(net10908),
    .X(_03198_));
 sg13g2_mux4_1 _20762_ (.S0(net10972),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][7] ),
    .S1(net10906),
    .X(_03199_));
 sg13g2_mux4_1 _20763_ (.S0(net10967),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][7] ),
    .S1(net10902),
    .X(_03200_));
 sg13g2_mux4_1 _20764_ (.S0(net10891),
    .A0(_03197_),
    .A1(_03198_),
    .A2(_03199_),
    .A3(_03200_),
    .S1(net10875),
    .X(_03201_));
 sg13g2_mux4_1 _20765_ (.S0(net10975),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][7] ),
    .S1(net10909),
    .X(_03202_));
 sg13g2_mux4_1 _20766_ (.S0(net10975),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][7] ),
    .S1(net10909),
    .X(_03203_));
 sg13g2_mux4_1 _20767_ (.S0(net10975),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][7] ),
    .S1(net10909),
    .X(_03204_));
 sg13g2_mux4_1 _20768_ (.S0(net10973),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][7] ),
    .S1(net10910),
    .X(_03205_));
 sg13g2_mux4_1 _20769_ (.S0(net10891),
    .A0(_03202_),
    .A1(_03203_),
    .A2(_03204_),
    .A3(_03205_),
    .S1(net10875),
    .X(_03206_));
 sg13g2_mux2_1 _20770_ (.A0(_03201_),
    .A1(_03206_),
    .S(net10881),
    .X(_03207_));
 sg13g2_a22oi_1 _20771_ (.Y(_03208_),
    .B1(_03207_),
    .B2(net10268),
    .A2(net10320),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[7] ));
 sg13g2_nor2_1 _20772_ (.A(net10272),
    .B(_03208_),
    .Y(_03209_));
 sg13g2_a221oi_1 _20773_ (.B2(net10701),
    .C1(_03209_),
    .B1(_03196_),
    .A1(_03190_),
    .Y(_03210_),
    .A2(_03191_));
 sg13g2_nor2_1 _20774_ (.A(net10334),
    .B(_03190_),
    .Y(_03211_));
 sg13g2_o21ai_1 _20775_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[7] ),
    .Y(_03212_),
    .A1(net9672),
    .A2(_03211_));
 sg13g2_o21ai_1 _20776_ (.B1(_03212_),
    .Y(_01924_),
    .A1(net9672),
    .A2(_03210_));
 sg13g2_nor2_1 _20777_ (.A(_00061_),
    .B(net10412),
    .Y(_03213_));
 sg13g2_a21oi_1 _20778_ (.A1(_11951_),
    .A2(net10412),
    .Y(_03214_),
    .B1(_03213_));
 sg13g2_mux2_1 _20779_ (.A0(_02224_),
    .A1(_03141_),
    .S(net10323),
    .X(_03215_));
 sg13g2_o21ai_1 _20780_ (.B1(_03215_),
    .Y(_03216_),
    .A1(net10290),
    .A2(_03214_));
 sg13g2_o21ai_1 _20781_ (.B1(_12006_),
    .Y(_03217_),
    .A1(_12025_),
    .A2(_12027_));
 sg13g2_nand2_1 _20782_ (.Y(_03218_),
    .A(_12007_),
    .B(_03217_));
 sg13g2_xnor2_1 _20783_ (.Y(_03219_),
    .A(net10669),
    .B(_03218_));
 sg13g2_nor2_1 _20784_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[8] ),
    .B(net10333),
    .Y(_03220_));
 sg13g2_mux4_1 _20785_ (.S0(_00005_),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][8] ),
    .S1(net10911),
    .X(_03221_));
 sg13g2_mux4_1 _20786_ (.S0(_00005_),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][8] ),
    .S1(net10911),
    .X(_03222_));
 sg13g2_mux4_1 _20787_ (.S0(net10954),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][8] ),
    .S1(net10911),
    .X(_03223_));
 sg13g2_mux4_1 _20788_ (.S0(_00005_),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][8] ),
    .S1(net10911),
    .X(_03224_));
 sg13g2_mux4_1 _20789_ (.S0(net10886),
    .A0(_03221_),
    .A1(_03222_),
    .A2(_03223_),
    .A3(_03224_),
    .S1(_00009_),
    .X(_03225_));
 sg13g2_mux4_1 _20790_ (.S0(net10958),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][8] ),
    .S1(net10895),
    .X(_03226_));
 sg13g2_mux4_1 _20791_ (.S0(net10958),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][8] ),
    .S1(net10895),
    .X(_03227_));
 sg13g2_mux4_1 _20792_ (.S0(net10958),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][8] ),
    .S1(net10895),
    .X(_03228_));
 sg13g2_mux4_1 _20793_ (.S0(net10958),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][8] ),
    .S1(_00006_),
    .X(_03229_));
 sg13g2_mux4_1 _20794_ (.S0(net10885),
    .A0(_03226_),
    .A1(_03227_),
    .A2(_03228_),
    .A3(_03229_),
    .S1(_00009_),
    .X(_03230_));
 sg13g2_mux2_1 _20795_ (.A0(_03225_),
    .A1(_03230_),
    .S(net10880),
    .X(_03231_));
 sg13g2_a22oi_1 _20796_ (.Y(_03232_),
    .B1(_03231_),
    .B2(net10266),
    .A2(_02186_),
    .A1(net10488));
 sg13g2_nor2_1 _20797_ (.A(net10271),
    .B(_03232_),
    .Y(_03233_));
 sg13g2_a221oi_1 _20798_ (.B2(_03220_),
    .C1(_03233_),
    .B1(_03219_),
    .A1(net10701),
    .Y(_03234_),
    .A2(_03216_));
 sg13g2_nor2_1 _20799_ (.A(net10333),
    .B(_03219_),
    .Y(_03235_));
 sg13g2_o21ai_1 _20800_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[8] ),
    .Y(_03236_),
    .A1(net9672),
    .A2(_03235_));
 sg13g2_o21ai_1 _20801_ (.B1(_03236_),
    .Y(_01925_),
    .A1(net9672),
    .A2(_03234_));
 sg13g2_nand2_1 _20802_ (.Y(_03237_),
    .A(_12010_),
    .B(_12028_));
 sg13g2_xor2_1 _20803_ (.B(_03237_),
    .A(net10668),
    .X(_03238_));
 sg13g2_nor2_1 _20804_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[9] ),
    .B(net10333),
    .Y(_03239_));
 sg13g2_mux4_1 _20805_ (.S0(net10967),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][9] ),
    .S1(net10902),
    .X(_03240_));
 sg13g2_mux4_1 _20806_ (.S0(net10970),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][9] ),
    .S1(net10908),
    .X(_03241_));
 sg13g2_mux4_1 _20807_ (.S0(net10972),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][9] ),
    .S1(net10906),
    .X(_03242_));
 sg13g2_mux4_1 _20808_ (.S0(net10967),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][9] ),
    .S1(net10902),
    .X(_03243_));
 sg13g2_mux4_1 _20809_ (.S0(net10891),
    .A0(_03240_),
    .A1(_03241_),
    .A2(_03242_),
    .A3(_03243_),
    .S1(net10875),
    .X(_03244_));
 sg13g2_mux4_1 _20810_ (.S0(net10975),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][9] ),
    .S1(net10909),
    .X(_03245_));
 sg13g2_mux4_1 _20811_ (.S0(net10974),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][9] ),
    .S1(net10905),
    .X(_03246_));
 sg13g2_mux4_1 _20812_ (.S0(net10975),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][9] ),
    .S1(net10909),
    .X(_03247_));
 sg13g2_mux4_1 _20813_ (.S0(net10973),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][9] ),
    .S1(net10910),
    .X(_03248_));
 sg13g2_mux4_1 _20814_ (.S0(net10891),
    .A0(_03245_),
    .A1(_03246_),
    .A2(_03247_),
    .A3(_03248_),
    .S1(net10875),
    .X(_03249_));
 sg13g2_mux2_1 _20815_ (.A0(_03244_),
    .A1(_03249_),
    .S(net10881),
    .X(_03250_));
 sg13g2_a22oi_1 _20816_ (.Y(_03251_),
    .B1(_03250_),
    .B2(net10266),
    .A2(net10320),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_pc[9] ));
 sg13g2_nor2_1 _20817_ (.A(net10293),
    .B(_03251_),
    .Y(_03252_));
 sg13g2_nand2b_1 _20818_ (.Y(_03253_),
    .B(net10322),
    .A_N(_00062_));
 sg13g2_o21ai_1 _20819_ (.B1(_03253_),
    .Y(_03254_),
    .A1(_00058_),
    .A2(net10322));
 sg13g2_and2_1 _20820_ (.A(net10411),
    .B(_02280_),
    .X(_03255_));
 sg13g2_a221oi_1 _20821_ (.B2(_02336_),
    .C1(_03255_),
    .B1(_03254_),
    .A1(net10322),
    .Y(_03256_),
    .A2(_03169_));
 sg13g2_nor2_1 _20822_ (.A(_09819_),
    .B(_03256_),
    .Y(_03257_));
 sg13g2_a221oi_1 _20823_ (.B2(_09819_),
    .C1(_03257_),
    .B1(_03252_),
    .A1(_03238_),
    .Y(_03258_),
    .A2(_03239_));
 sg13g2_nor2_1 _20824_ (.A(net10333),
    .B(_03238_),
    .Y(_03259_));
 sg13g2_o21ai_1 _20825_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[9] ),
    .Y(_03260_),
    .A1(net9671),
    .A2(_03259_));
 sg13g2_o21ai_1 _20826_ (.B1(_03260_),
    .Y(_01926_),
    .A1(net9671),
    .A2(_03258_));
 sg13g2_buf_2 place10228 (.A(net10227),
    .X(net10228));
 sg13g2_buf_2 place10195 (.A(_06720_),
    .X(net10195));
 sg13g2_mux4_1 _20829_ (.S0(net10833),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][0] ),
    .S1(net10815),
    .X(_03263_));
 sg13g2_mux4_1 _20830_ (.S0(_00000_),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][0] ),
    .S1(_00001_),
    .X(_03264_));
 sg13g2_mux4_1 _20831_ (.S0(_00000_),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][0] ),
    .S1(net10784),
    .X(_03265_));
 sg13g2_mux4_1 _20832_ (.S0(net10833),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][0] ),
    .S1(net10815),
    .X(_03266_));
 sg13g2_mux4_1 _20833_ (.S0(_00002_),
    .A0(_03263_),
    .A1(_03264_),
    .A2(_03265_),
    .A3(_03266_),
    .S1(net10771),
    .X(_03267_));
 sg13g2_mux4_1 _20834_ (.S0(net10833),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][0] ),
    .S1(net10815),
    .X(_03268_));
 sg13g2_mux4_1 _20835_ (.S0(net10827),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][0] ),
    .S1(net10808),
    .X(_03269_));
 sg13g2_mux4_1 _20836_ (.S0(net10833),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][0] ),
    .S1(net10815),
    .X(_03270_));
 sg13g2_mux4_1 _20837_ (.S0(_00000_),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][0] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][0] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][0] ),
    .S1(_00001_),
    .X(_03271_));
 sg13g2_mux4_1 _20838_ (.S0(net10778),
    .A0(_03268_),
    .A1(_03269_),
    .A2(_03270_),
    .A3(_03271_),
    .S1(net10772),
    .X(_03272_));
 sg13g2_mux2_1 _20839_ (.A0(_03267_),
    .A1(_03272_),
    .S(_00004_),
    .X(_03273_));
 sg13g2_nand2_2 _20840_ (.Y(_03274_),
    .A(_08872_),
    .B(_03273_));
 sg13g2_nor2_1 _20841_ (.A(net10418),
    .B(_03274_),
    .Y(_03275_));
 sg13g2_a21oi_2 _20842_ (.B1(_03275_),
    .Y(_03276_),
    .A2(net10418),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[0] ));
 sg13g2_buf_2 place10352 (.A(net10351),
    .X(net10352));
 sg13g2_nand2_1 _20844_ (.Y(_03278_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[0] ),
    .B(net10425));
 sg13g2_o21ai_1 _20845_ (.B1(_03278_),
    .Y(_01927_),
    .A1(net10425),
    .A2(_03276_));
 sg13g2_inv_4 _20846_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[10] ),
    .Y(_03279_));
 sg13g2_buf_2 place10428 (.A(net10427),
    .X(net10428));
 sg13g2_buf_2 place10280 (.A(net10279),
    .X(net10280));
 sg13g2_buf_2 place10377 (.A(net10376),
    .X(net10377));
 sg13g2_buf_2 place10224 (.A(net10222),
    .X(net10224));
 sg13g2_buf_2 place10250 (.A(net10248),
    .X(net10250));
 sg13g2_buf_2 place10194 (.A(_06783_),
    .X(net10194));
 sg13g2_mux4_1 _20853_ (.S0(net10832),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][10] ),
    .S1(net10809),
    .X(_03286_));
 sg13g2_mux4_1 _20854_ (.S0(net10832),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][10] ),
    .S1(net10809),
    .X(_03287_));
 sg13g2_buf_2 place10238 (.A(net10235),
    .X(net10238));
 sg13g2_buf_16 clkbuf_leaf_320_clk (.X(clknet_leaf_320_clk),
    .A(clknet_8_92_0_clk));
 sg13g2_mux4_1 _20857_ (.S0(net10832),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][10] ),
    .S1(net10809),
    .X(_03290_));
 sg13g2_buf_16 clkbuf_leaf_319_clk (.X(clknet_leaf_319_clk),
    .A(clknet_8_89_0_clk));
 sg13g2_buf_2 place10221 (.A(net10219),
    .X(net10221));
 sg13g2_mux4_1 _20860_ (.S0(net10832),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][10] ),
    .S1(net10809),
    .X(_03293_));
 sg13g2_buf_2 place10208 (.A(net10207),
    .X(net10208));
 sg13g2_buf_2 place10220 (.A(net10219),
    .X(net10220));
 sg13g2_buf_16 clkbuf_leaf_321_clk (.X(clknet_leaf_321_clk),
    .A(clknet_8_91_0_clk));
 sg13g2_mux4_1 _20864_ (.S0(net10779),
    .A0(_03286_),
    .A1(_03287_),
    .A2(_03290_),
    .A3(_03293_),
    .S1(net10768),
    .X(_03297_));
 sg13g2_mux4_1 _20865_ (.S0(net10830),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][10] ),
    .S1(net10814),
    .X(_03298_));
 sg13g2_mux4_1 _20866_ (.S0(net10829),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][10] ),
    .S1(net10813),
    .X(_03299_));
 sg13g2_buf_2 place10201 (.A(net10200),
    .X(net10201));
 sg13g2_buf_2 place10214 (.A(net10213),
    .X(net10214));
 sg13g2_mux4_1 _20869_ (.S0(net10827),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][10] ),
    .S1(net10811),
    .X(_03302_));
 sg13g2_buf_2 place10192 (.A(_06847_),
    .X(net10192));
 sg13g2_buf_2 place10213 (.A(net10212),
    .X(net10213));
 sg13g2_mux4_1 _20872_ (.S0(net10827),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][10] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][10] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][10] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][10] ),
    .S1(net10811),
    .X(_03305_));
 sg13g2_mux4_1 _20873_ (.S0(net10780),
    .A0(_03298_),
    .A1(_03299_),
    .A2(_03302_),
    .A3(_03305_),
    .S1(net10768),
    .X(_03306_));
 sg13g2_buf_2 place10219 (.A(net10218),
    .X(net10219));
 sg13g2_mux2_1 _20875_ (.A0(_03297_),
    .A1(_03306_),
    .S(net10772),
    .X(_03308_));
 sg13g2_a21oi_2 _20876_ (.B1(_08348_),
    .Y(_03309_),
    .A2(_08871_),
    .A1(_00131_));
 sg13g2_buf_2 place10187 (.A(_07153_),
    .X(net10187));
 sg13g2_buf_2 place10193 (.A(_06825_),
    .X(net10193));
 sg13g2_a221oi_1 _20879_ (.B2(_03309_),
    .C1(net10422),
    .B1(_03308_),
    .A1(net10694),
    .Y(_03312_),
    .A2(net10416));
 sg13g2_a21oi_1 _20880_ (.A1(_03279_),
    .A2(net10422),
    .Y(_01928_),
    .B1(_03312_));
 sg13g2_buf_2 place10199 (.A(_11808_),
    .X(net10199));
 sg13g2_buf_2 place10200 (.A(net10199),
    .X(net10200));
 sg13g2_buf_16 clkbuf_leaf_322_clk (.X(clknet_leaf_322_clk),
    .A(clknet_8_93_0_clk));
 sg13g2_buf_2 place10188 (.A(_07153_),
    .X(net10188));
 sg13g2_buf_2 place10191 (.A(_06866_),
    .X(net10191));
 sg13g2_mux4_1 _20886_ (.S0(net10858),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][11] ),
    .S1(net10796),
    .X(_03318_));
 sg13g2_buf_2 place10242 (.A(_07931_),
    .X(net10242));
 sg13g2_buf_2 place10189 (.A(net10188),
    .X(net10189));
 sg13g2_mux4_1 _20889_ (.S0(net10858),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][11] ),
    .S1(net10796),
    .X(_03321_));
 sg13g2_buf_2 place10190 (.A(net10189),
    .X(net10190));
 sg13g2_buf_2 place10183 (.A(_08420_),
    .X(net10183));
 sg13g2_buf_2 place10186 (.A(_08408_),
    .X(net10186));
 sg13g2_buf_2 place10181 (.A(_10080_),
    .X(net10181));
 sg13g2_mux4_1 _20894_ (.S0(net10857),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][11] ),
    .S1(net10795),
    .X(_03326_));
 sg13g2_buf_2 place10180 (.A(net10179),
    .X(net10180));
 sg13g2_buf_2 place10177 (.A(net10175),
    .X(net10177));
 sg13g2_mux4_1 _20897_ (.S0(net10859),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][11] ),
    .S1(net10797),
    .X(_03329_));
 sg13g2_buf_16 clkbuf_leaf_331_clk (.X(clknet_leaf_331_clk),
    .A(clknet_8_115_0_clk));
 sg13g2_buf_16 clkbuf_leaf_330_clk (.X(clknet_leaf_330_clk),
    .A(clknet_8_116_0_clk));
 sg13g2_mux4_1 _20900_ (.S0(net10776),
    .A0(_03318_),
    .A1(_03321_),
    .A2(_03326_),
    .A3(_03329_),
    .S1(net10766),
    .X(_03332_));
 sg13g2_buf_16 clkbuf_leaf_329_clk (.X(clknet_leaf_329_clk),
    .A(clknet_8_113_0_clk));
 sg13g2_buf_2 place10182 (.A(net10181),
    .X(net10182));
 sg13g2_mux4_1 _20903_ (.S0(net10858),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][11] ),
    .S1(net10796),
    .X(_03335_));
 sg13g2_buf_2 place10175 (.A(net10174),
    .X(net10175));
 sg13g2_buf_2 place10172 (.A(net10170),
    .X(net10172));
 sg13g2_mux4_1 _20906_ (.S0(net10858),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][11] ),
    .S1(net10796),
    .X(_03338_));
 sg13g2_buf_16 clkbuf_leaf_328_clk (.X(clknet_leaf_328_clk),
    .A(clknet_8_113_0_clk));
 sg13g2_buf_2 place10185 (.A(_08420_),
    .X(net10185));
 sg13g2_mux4_1 _20909_ (.S0(net10858),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][11] ),
    .S1(net10796),
    .X(_03341_));
 sg13g2_buf_2 place10184 (.A(net10183),
    .X(net10184));
 sg13g2_buf_16 clkbuf_leaf_325_clk (.X(clknet_leaf_325_clk),
    .A(clknet_8_113_0_clk));
 sg13g2_mux4_1 _20912_ (.S0(net10859),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][11] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][11] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][11] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][11] ),
    .S1(net10797),
    .X(_03344_));
 sg13g2_buf_16 clkbuf_leaf_323_clk (.X(clknet_leaf_323_clk),
    .A(clknet_8_93_0_clk));
 sg13g2_buf_2 place10173 (.A(net10170),
    .X(net10173));
 sg13g2_mux4_1 _20915_ (.S0(net10776),
    .A0(_03335_),
    .A1(_03338_),
    .A2(_03341_),
    .A3(_03344_),
    .S1(net10766),
    .X(_03347_));
 sg13g2_buf_2 place10168 (.A(net10166),
    .X(net10168));
 sg13g2_mux2_1 _20917_ (.A0(_03332_),
    .A1(_03347_),
    .S(net10771),
    .X(_03349_));
 sg13g2_a22oi_1 _20918_ (.Y(_03350_),
    .B1(net10261),
    .B2(_03349_),
    .A2(net10416),
    .A1(net10693));
 sg13g2_nand2_1 _20919_ (.Y(_03351_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[11] ),
    .B(net10422));
 sg13g2_o21ai_1 _20920_ (.B1(_03351_),
    .Y(_01929_),
    .A1(net10422),
    .A2(_03350_));
 sg13g2_inv_2 _20921_ (.Y(_03352_),
    .A(net10518));
 sg13g2_buf_2 place10768 (.A(_00004_),
    .X(net10768));
 sg13g2_mux4_1 _20923_ (.S0(net10836),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][12] ),
    .S1(net10818),
    .X(_03354_));
 sg13g2_mux4_1 _20924_ (.S0(net10837),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][12] ),
    .S1(net10819),
    .X(_03355_));
 sg13g2_buf_2 place10179 (.A(_10080_),
    .X(net10179));
 sg13g2_buf_2 place10225 (.A(_10047_),
    .X(net10225));
 sg13g2_mux4_1 _20927_ (.S0(net10836),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][12] ),
    .S1(net10818),
    .X(_03358_));
 sg13g2_mux4_1 _20928_ (.S0(net10839),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][12] ),
    .S1(net10821),
    .X(_03359_));
 sg13g2_buf_2 place10769 (.A(_00004_),
    .X(net10769));
 sg13g2_buf_2 place10249 (.A(net10248),
    .X(net10249));
 sg13g2_mux4_1 _20931_ (.S0(net10783),
    .A0(_03354_),
    .A1(_03355_),
    .A2(_03358_),
    .A3(_03359_),
    .S1(net10763),
    .X(_03362_));
 sg13g2_mux4_1 _20932_ (.S0(net10835),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][12] ),
    .S1(net10818),
    .X(_03363_));
 sg13g2_mux4_1 _20933_ (.S0(net10835),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][12] ),
    .S1(net10818),
    .X(_03364_));
 sg13g2_buf_2 place10339 (.A(net10337),
    .X(net10339));
 sg13g2_buf_2 place10223 (.A(net10222),
    .X(net10223));
 sg13g2_mux4_1 _20936_ (.S0(net10839),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][12] ),
    .S1(net10821),
    .X(_03367_));
 sg13g2_buf_2 place10222 (.A(_10047_),
    .X(net10222));
 sg13g2_buf_2 place10241 (.A(net10240),
    .X(net10241));
 sg13g2_mux4_1 _20939_ (.S0(net10839),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][12] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][12] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][12] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][12] ),
    .S1(net10821),
    .X(_03370_));
 sg13g2_buf_2 place10229 (.A(net10228),
    .X(net10229));
 sg13g2_buf_2 place10248 (.A(net10247),
    .X(net10248));
 sg13g2_mux4_1 _20942_ (.S0(net10783),
    .A0(_03363_),
    .A1(_03364_),
    .A2(_03367_),
    .A3(_03370_),
    .S1(net10763),
    .X(_03373_));
 sg13g2_mux2_1 _20943_ (.A0(_03362_),
    .A1(_03373_),
    .S(_00003_),
    .X(_03374_));
 sg13g2_a221oi_1 _20944_ (.B2(_03374_),
    .C1(net10423),
    .B1(_03309_),
    .A1(net10692),
    .Y(_03375_),
    .A2(net10418));
 sg13g2_a21oi_1 _20945_ (.A1(_03352_),
    .A2(net10422),
    .Y(_01930_),
    .B1(_03375_));
 sg13g2_buf_2 place10252 (.A(_07207_),
    .X(net10252));
 sg13g2_buf_2 place10247 (.A(net10246),
    .X(net10247));
 sg13g2_buf_2 place10174 (.A(_10088_),
    .X(net10174));
 sg13g2_mux4_1 _20949_ (.S0(net10841),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][13] ),
    .S1(net10822),
    .X(_03379_));
 sg13g2_mux4_1 _20950_ (.S0(net10834),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][13] ),
    .S1(net10816),
    .X(_03380_));
 sg13g2_mux4_1 _20951_ (.S0(net10834),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][13] ),
    .S1(net10815),
    .X(_03381_));
 sg13g2_mux4_1 _20952_ (.S0(net10841),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][13] ),
    .S1(net10822),
    .X(_03382_));
 sg13g2_mux4_1 _20953_ (.S0(net10782),
    .A0(_03379_),
    .A1(_03380_),
    .A2(_03381_),
    .A3(_03382_),
    .S1(net10762),
    .X(_03383_));
 sg13g2_mux4_1 _20954_ (.S0(net10834),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][13] ),
    .S1(net10816),
    .X(_03384_));
 sg13g2_mux4_1 _20955_ (.S0(net10834),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][13] ),
    .S1(net10816),
    .X(_03385_));
 sg13g2_mux4_1 _20956_ (.S0(net10834),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][13] ),
    .S1(net10816),
    .X(_03386_));
 sg13g2_mux4_1 _20957_ (.S0(net10833),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][13] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][13] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][13] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][13] ),
    .S1(net10815),
    .X(_03387_));
 sg13g2_mux4_1 _20958_ (.S0(net10782),
    .A0(_03384_),
    .A1(_03385_),
    .A2(_03386_),
    .A3(_03387_),
    .S1(net10762),
    .X(_03388_));
 sg13g2_mux2_1 _20959_ (.A0(_03383_),
    .A1(_03388_),
    .S(_00003_),
    .X(_03389_));
 sg13g2_a221oi_1 _20960_ (.B2(_03389_),
    .C1(net10421),
    .B1(net10261),
    .A1(net10691),
    .Y(_03390_),
    .A2(net10416));
 sg13g2_a21oi_1 _20961_ (.A1(_08752_),
    .A2(net10422),
    .Y(_01931_),
    .B1(_03390_));
 sg13g2_mux4_1 _20962_ (.S0(net10854),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][14] ),
    .S1(net10793),
    .X(_03391_));
 sg13g2_mux4_1 _20963_ (.S0(net10854),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][14] ),
    .S1(net10793),
    .X(_03392_));
 sg13g2_mux4_1 _20964_ (.S0(net10854),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][14] ),
    .S1(net10793),
    .X(_03393_));
 sg13g2_mux4_1 _20965_ (.S0(net10854),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][14] ),
    .S1(net10793),
    .X(_03394_));
 sg13g2_mux4_1 _20966_ (.S0(net10775),
    .A0(_03391_),
    .A1(_03392_),
    .A2(_03393_),
    .A3(_03394_),
    .S1(net10764),
    .X(_03395_));
 sg13g2_mux4_1 _20967_ (.S0(net10854),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][14] ),
    .S1(net10793),
    .X(_03396_));
 sg13g2_mux4_1 _20968_ (.S0(net10845),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][14] ),
    .S1(net10795),
    .X(_03397_));
 sg13g2_mux4_1 _20969_ (.S0(net10845),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][14] ),
    .S1(net10785),
    .X(_03398_));
 sg13g2_mux4_1 _20970_ (.S0(net10845),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][14] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][14] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][14] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][14] ),
    .S1(net10795),
    .X(_03399_));
 sg13g2_mux4_1 _20971_ (.S0(_00002_),
    .A0(_03396_),
    .A1(_03397_),
    .A2(_03398_),
    .A3(_03399_),
    .S1(net10764),
    .X(_03400_));
 sg13g2_mux2_1 _20972_ (.A0(_03395_),
    .A1(_03400_),
    .S(net10774),
    .X(_03401_));
 sg13g2_a22oi_1 _20973_ (.Y(_03402_),
    .B1(net10262),
    .B2(_03401_),
    .A2(net10416),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[14] ));
 sg13g2_nand2_1 _20974_ (.Y(_03403_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[14] ),
    .B(net10421));
 sg13g2_o21ai_1 _20975_ (.B1(_03403_),
    .Y(_01932_),
    .A1(net10421),
    .A2(_03402_));
 sg13g2_mux4_1 _20976_ (.S0(net10830),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][15] ),
    .S1(net10814),
    .X(_03404_));
 sg13g2_mux4_1 _20977_ (.S0(net10830),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][15] ),
    .S1(net10814),
    .X(_03405_));
 sg13g2_mux4_1 _20978_ (.S0(net10830),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][15] ),
    .S1(net10814),
    .X(_03406_));
 sg13g2_buf_2 place10163 (.A(_11413_),
    .X(net10163));
 sg13g2_buf_2 place10240 (.A(net10239),
    .X(net10240));
 sg13g2_mux4_1 _20981_ (.S0(net10830),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][15] ),
    .S1(net10814),
    .X(_03409_));
 sg13g2_mux4_1 _20982_ (.S0(net10780),
    .A0(_03404_),
    .A1(_03405_),
    .A2(_03406_),
    .A3(_03409_),
    .S1(net10768),
    .X(_03410_));
 sg13g2_mux4_1 _20983_ (.S0(net10830),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][15] ),
    .S1(net10814),
    .X(_03411_));
 sg13g2_mux4_1 _20984_ (.S0(net10840),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][15] ),
    .S1(net10823),
    .X(_03412_));
 sg13g2_mux4_1 _20985_ (.S0(net10844),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][15] ),
    .S1(net10826),
    .X(_03413_));
 sg13g2_mux4_1 _20986_ (.S0(net10828),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][15] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][15] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][15] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][15] ),
    .S1(net10812),
    .X(_03414_));
 sg13g2_mux4_1 _20987_ (.S0(net10780),
    .A0(_03411_),
    .A1(_03412_),
    .A2(_03413_),
    .A3(_03414_),
    .S1(net10768),
    .X(_03415_));
 sg13g2_mux2_1 _20988_ (.A0(_03410_),
    .A1(_03415_),
    .S(net10770),
    .X(_03416_));
 sg13g2_a221oi_1 _20989_ (.B2(_03416_),
    .C1(net10421),
    .B1(net10261),
    .A1(net10690),
    .Y(_03417_),
    .A2(net10416));
 sg13g2_a21oi_1 _20990_ (.A1(_08770_),
    .A2(net10421),
    .Y(_01933_),
    .B1(_03417_));
 sg13g2_mux4_1 _20991_ (.S0(net10828),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][16] ),
    .S1(net10812),
    .X(_03418_));
 sg13g2_mux4_1 _20992_ (.S0(net10828),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][16] ),
    .S1(net10808),
    .X(_03419_));
 sg13g2_mux4_1 _20993_ (.S0(net10828),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][16] ),
    .S1(net10812),
    .X(_03420_));
 sg13g2_mux4_1 _20994_ (.S0(net10827),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][16] ),
    .S1(net10811),
    .X(_03421_));
 sg13g2_mux4_1 _20995_ (.S0(net10779),
    .A0(_03418_),
    .A1(_03419_),
    .A2(_03420_),
    .A3(_03421_),
    .S1(_00004_),
    .X(_03422_));
 sg13g2_mux4_1 _20996_ (.S0(net10828),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][16] ),
    .S1(net10812),
    .X(_03423_));
 sg13g2_mux4_1 _20997_ (.S0(net10828),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][16] ),
    .S1(net10812),
    .X(_03424_));
 sg13g2_mux4_1 _20998_ (.S0(net10831),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][16] ),
    .S1(net10808),
    .X(_03425_));
 sg13g2_mux4_1 _20999_ (.S0(net10831),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][16] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][16] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][16] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][16] ),
    .S1(net10808),
    .X(_03426_));
 sg13g2_mux4_1 _21000_ (.S0(net10779),
    .A0(_03423_),
    .A1(_03424_),
    .A2(_03425_),
    .A3(_03426_),
    .S1(_00004_),
    .X(_03427_));
 sg13g2_mux2_1 _21001_ (.A0(_03422_),
    .A1(_03427_),
    .S(net10772),
    .X(_03428_));
 sg13g2_a221oi_1 _21002_ (.B2(_03428_),
    .C1(net10421),
    .B1(net10261),
    .A1(net10689),
    .Y(_03429_),
    .A2(net10416));
 sg13g2_a21oi_1 _21003_ (.A1(_11840_),
    .A2(net10420),
    .Y(_01934_),
    .B1(_03429_));
 sg13g2_mux4_1 _21004_ (.S0(net10841),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][17] ),
    .S1(net10822),
    .X(_03430_));
 sg13g2_mux4_1 _21005_ (.S0(net10841),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][17] ),
    .S1(net10822),
    .X(_03431_));
 sg13g2_mux4_1 _21006_ (.S0(net10841),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][17] ),
    .S1(net10822),
    .X(_03432_));
 sg13g2_mux4_1 _21007_ (.S0(net10834),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][17] ),
    .S1(net10816),
    .X(_03433_));
 sg13g2_mux4_1 _21008_ (.S0(net10782),
    .A0(_03430_),
    .A1(_03431_),
    .A2(_03432_),
    .A3(_03433_),
    .S1(net10762),
    .X(_03434_));
 sg13g2_mux4_1 _21009_ (.S0(net10841),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][17] ),
    .S1(net10822),
    .X(_03435_));
 sg13g2_mux4_1 _21010_ (.S0(net10841),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][17] ),
    .S1(net10822),
    .X(_03436_));
 sg13g2_mux4_1 _21011_ (.S0(net10834),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][17] ),
    .S1(net10816),
    .X(_03437_));
 sg13g2_mux4_1 _21012_ (.S0(net10836),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][17] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][17] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][17] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][17] ),
    .S1(net10817),
    .X(_03438_));
 sg13g2_mux4_1 _21013_ (.S0(net10782),
    .A0(_03435_),
    .A1(_03436_),
    .A2(_03437_),
    .A3(_03438_),
    .S1(net10762),
    .X(_03439_));
 sg13g2_mux2_1 _21014_ (.A0(_03434_),
    .A1(_03439_),
    .S(net10770),
    .X(_03440_));
 sg13g2_a221oi_1 _21015_ (.B2(_03440_),
    .C1(net10420),
    .B1(net10262),
    .A1(net10688),
    .Y(_03441_),
    .A2(_08348_));
 sg13g2_a21oi_1 _21016_ (.A1(_11845_),
    .A2(net10420),
    .Y(_01935_),
    .B1(_03441_));
 sg13g2_mux4_1 _21017_ (.S0(net10850),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][18] ),
    .S1(net10786),
    .X(_03442_));
 sg13g2_mux4_1 _21018_ (.S0(net10852),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][18] ),
    .S1(net10792),
    .X(_03443_));
 sg13g2_mux4_1 _21019_ (.S0(net10847),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][18] ),
    .S1(net10787),
    .X(_03444_));
 sg13g2_mux4_1 _21020_ (.S0(net10847),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][18] ),
    .S1(net10787),
    .X(_03445_));
 sg13g2_mux4_1 _21021_ (.S0(net10778),
    .A0(_03442_),
    .A1(_03443_),
    .A2(_03444_),
    .A3(_03445_),
    .S1(net10769),
    .X(_03446_));
 sg13g2_mux4_1 _21022_ (.S0(net10846),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][18] ),
    .S1(net10787),
    .X(_03447_));
 sg13g2_mux4_1 _21023_ (.S0(net10846),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][18] ),
    .S1(net10784),
    .X(_03448_));
 sg13g2_mux4_1 _21024_ (.S0(net10850),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][18] ),
    .S1(net10786),
    .X(_03449_));
 sg13g2_mux4_1 _21025_ (.S0(net10850),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][18] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][18] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][18] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][18] ),
    .S1(net10786),
    .X(_03450_));
 sg13g2_mux4_1 _21026_ (.S0(net10778),
    .A0(_03447_),
    .A1(_03448_),
    .A2(_03449_),
    .A3(_03450_),
    .S1(_00004_),
    .X(_03451_));
 sg13g2_mux2_1 _21027_ (.A0(_03446_),
    .A1(_03451_),
    .S(net10773),
    .X(_03452_));
 sg13g2_a221oi_1 _21028_ (.B2(_03452_),
    .C1(net10420),
    .B1(net10262),
    .A1(net10687),
    .Y(_03453_),
    .A2(net10414));
 sg13g2_a21oi_1 _21029_ (.A1(_08786_),
    .A2(net10420),
    .Y(_01936_),
    .B1(_03453_));
 sg13g2_mux4_1 _21030_ (.S0(net10863),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][19] ),
    .S1(net10801),
    .X(_03454_));
 sg13g2_mux4_1 _21031_ (.S0(net10863),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][19] ),
    .S1(net10801),
    .X(_03455_));
 sg13g2_mux4_1 _21032_ (.S0(net10863),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][19] ),
    .S1(net10801),
    .X(_03456_));
 sg13g2_mux4_1 _21033_ (.S0(net10863),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][19] ),
    .S1(net10801),
    .X(_03457_));
 sg13g2_mux4_1 _21034_ (.S0(net10777),
    .A0(_03454_),
    .A1(_03455_),
    .A2(_03456_),
    .A3(_03457_),
    .S1(net10767),
    .X(_03458_));
 sg13g2_mux4_1 _21035_ (.S0(net10867),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][19] ),
    .S1(net10805),
    .X(_03459_));
 sg13g2_buf_2 place10207 (.A(_11625_),
    .X(net10207));
 sg13g2_buf_2 place10209 (.A(net10207),
    .X(net10209));
 sg13g2_mux4_1 _21038_ (.S0(net10868),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][19] ),
    .S1(net10807),
    .X(_03462_));
 sg13g2_buf_2 place10212 (.A(_11625_),
    .X(net10212));
 sg13g2_buf_2 place10211 (.A(net10210),
    .X(net10211));
 sg13g2_mux4_1 _21041_ (.S0(net10868),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][19] ),
    .S1(net10807),
    .X(_03465_));
 sg13g2_mux4_1 _21042_ (.S0(net10868),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][19] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][19] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][19] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][19] ),
    .S1(net10807),
    .X(_03466_));
 sg13g2_mux4_1 _21043_ (.S0(net10777),
    .A0(_03459_),
    .A1(_03462_),
    .A2(_03465_),
    .A3(_03466_),
    .S1(net10767),
    .X(_03467_));
 sg13g2_mux2_1 _21044_ (.A0(_03458_),
    .A1(_03467_),
    .S(net10774),
    .X(_03468_));
 sg13g2_a22oi_1 _21045_ (.Y(_03469_),
    .B1(net10263),
    .B2(_03468_),
    .A2(net10415),
    .A1(net10686));
 sg13g2_nand2_1 _21046_ (.Y(_03470_),
    .A(net10514),
    .B(net10426));
 sg13g2_o21ai_1 _21047_ (.B1(_03470_),
    .Y(_01937_),
    .A1(net10426),
    .A2(_03469_));
 sg13g2_buf_2 place10167 (.A(net10166),
    .X(net10167));
 sg13g2_mux4_1 _21049_ (.S0(net10836),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][1] ),
    .S1(net10817),
    .X(_03472_));
 sg13g2_mux4_1 _21050_ (.S0(net10836),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][1] ),
    .S1(net10817),
    .X(_03473_));
 sg13g2_mux4_1 _21051_ (.S0(net10836),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][1] ),
    .S1(net10818),
    .X(_03474_));
 sg13g2_mux4_1 _21052_ (.S0(net10839),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][1] ),
    .S1(net10821),
    .X(_03475_));
 sg13g2_mux4_1 _21053_ (.S0(net10782),
    .A0(_03472_),
    .A1(_03473_),
    .A2(_03474_),
    .A3(_03475_),
    .S1(net10770),
    .X(_03476_));
 sg13g2_mux4_1 _21054_ (.S0(net10836),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][1] ),
    .S1(net10817),
    .X(_03477_));
 sg13g2_mux4_1 _21055_ (.S0(net10835),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][1] ),
    .S1(net10817),
    .X(_03478_));
 sg13g2_mux4_1 _21056_ (.S0(net10839),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][1] ),
    .S1(net10821),
    .X(_03479_));
 sg13g2_mux4_1 _21057_ (.S0(net10835),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][1] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][1] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][1] ),
    .S1(net10817),
    .X(_03480_));
 sg13g2_mux4_1 _21058_ (.S0(net10782),
    .A0(_03477_),
    .A1(_03478_),
    .A2(_03479_),
    .A3(_03480_),
    .S1(net10770),
    .X(_03481_));
 sg13g2_mux2_1 _21059_ (.A0(_03476_),
    .A1(_03481_),
    .S(net10762),
    .X(_03482_));
 sg13g2_nand2_2 _21060_ (.Y(_03483_),
    .A(_08872_),
    .B(_03482_));
 sg13g2_nand2_1 _21061_ (.Y(_03484_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[1] ),
    .B(net10419));
 sg13g2_o21ai_1 _21062_ (.B1(_03484_),
    .Y(_03485_),
    .A1(net10419),
    .A2(_03483_));
 sg13g2_nor2_1 _21063_ (.A(net10425),
    .B(_03485_),
    .Y(_03486_));
 sg13g2_a21oi_1 _21064_ (.A1(_08682_),
    .A2(net10425),
    .Y(_01938_),
    .B1(_03486_));
 sg13g2_mux4_1 _21065_ (.S0(net10850),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][20] ),
    .S1(net10786),
    .X(_03487_));
 sg13g2_mux4_1 _21066_ (.S0(net10852),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][20] ),
    .S1(net10792),
    .X(_03488_));
 sg13g2_mux4_1 _21067_ (.S0(net10847),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][20] ),
    .S1(net10788),
    .X(_03489_));
 sg13g2_mux4_1 _21068_ (.S0(net10846),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][20] ),
    .S1(net10787),
    .X(_03490_));
 sg13g2_mux4_1 _21069_ (.S0(net10778),
    .A0(_03487_),
    .A1(_03488_),
    .A2(_03489_),
    .A3(_03490_),
    .S1(net10769),
    .X(_03491_));
 sg13g2_mux4_1 _21070_ (.S0(net10847),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][20] ),
    .S1(net10788),
    .X(_03492_));
 sg13g2_mux4_1 _21071_ (.S0(net10847),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][20] ),
    .S1(net10788),
    .X(_03493_));
 sg13g2_mux4_1 _21072_ (.S0(net10847),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][20] ),
    .S1(net10788),
    .X(_03494_));
 sg13g2_mux4_1 _21073_ (.S0(net10847),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][20] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][20] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][20] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][20] ),
    .S1(net10788),
    .X(_03495_));
 sg13g2_mux4_1 _21074_ (.S0(net10781),
    .A0(_03492_),
    .A1(_03493_),
    .A2(_03494_),
    .A3(_03495_),
    .S1(net10769),
    .X(_03496_));
 sg13g2_mux2_1 _21075_ (.A0(_03491_),
    .A1(_03496_),
    .S(net10773),
    .X(_03497_));
 sg13g2_a221oi_1 _21076_ (.B2(_03497_),
    .C1(net10426),
    .B1(net10262),
    .A1(net10685),
    .Y(_03498_),
    .A2(net10414));
 sg13g2_a21oi_1 _21077_ (.A1(_11862_),
    .A2(net10426),
    .Y(_01939_),
    .B1(_03498_));
 sg13g2_mux4_1 _21078_ (.S0(net10850),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][21] ),
    .S1(net10786),
    .X(_03499_));
 sg13g2_mux4_1 _21079_ (.S0(net10852),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][21] ),
    .S1(net10792),
    .X(_03500_));
 sg13g2_mux4_1 _21080_ (.S0(net10847),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][21] ),
    .S1(net10788),
    .X(_03501_));
 sg13g2_mux4_1 _21081_ (.S0(net10846),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][21] ),
    .S1(net10787),
    .X(_03502_));
 sg13g2_mux4_1 _21082_ (.S0(net10778),
    .A0(_03499_),
    .A1(_03500_),
    .A2(_03501_),
    .A3(_03502_),
    .S1(net10769),
    .X(_03503_));
 sg13g2_mux4_1 _21083_ (.S0(net10852),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][21] ),
    .S1(net10792),
    .X(_03504_));
 sg13g2_mux4_1 _21084_ (.S0(net10852),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][21] ),
    .S1(net10792),
    .X(_03505_));
 sg13g2_mux4_1 _21085_ (.S0(net10852),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][21] ),
    .S1(net10792),
    .X(_03506_));
 sg13g2_mux4_1 _21086_ (.S0(net10852),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][21] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][21] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][21] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][21] ),
    .S1(net10792),
    .X(_03507_));
 sg13g2_mux4_1 _21087_ (.S0(net10781),
    .A0(_03504_),
    .A1(_03505_),
    .A2(_03506_),
    .A3(_03507_),
    .S1(net10769),
    .X(_03508_));
 sg13g2_mux2_1 _21088_ (.A0(_03503_),
    .A1(_03508_),
    .S(net10773),
    .X(_03509_));
 sg13g2_a221oi_1 _21089_ (.B2(_03509_),
    .C1(net10426),
    .B1(net10262),
    .A1(net10684),
    .Y(_03510_),
    .A2(net10414));
 sg13g2_a21oi_1 _21090_ (.A1(_08801_),
    .A2(net10426),
    .Y(_01940_),
    .B1(_03510_));
 sg13g2_mux4_1 _21091_ (.S0(net10856),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][22] ),
    .S1(net10794),
    .X(_03511_));
 sg13g2_mux4_1 _21092_ (.S0(net10849),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][22] ),
    .S1(net10791),
    .X(_03512_));
 sg13g2_mux4_1 _21093_ (.S0(net10849),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][22] ),
    .S1(net10791),
    .X(_03513_));
 sg13g2_mux4_1 _21094_ (.S0(net10856),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][22] ),
    .S1(net10794),
    .X(_03514_));
 sg13g2_mux4_1 _21095_ (.S0(net10781),
    .A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S1(net10764),
    .X(_03515_));
 sg13g2_mux4_1 _21096_ (.S0(net10848),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][22] ),
    .S1(net10790),
    .X(_03516_));
 sg13g2_mux4_1 _21097_ (.S0(net10848),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][22] ),
    .S1(net10790),
    .X(_03517_));
 sg13g2_mux4_1 _21098_ (.S0(net10848),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][22] ),
    .S1(net10790),
    .X(_03518_));
 sg13g2_mux4_1 _21099_ (.S0(net10848),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][22] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][22] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][22] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][22] ),
    .S1(net10790),
    .X(_03519_));
 sg13g2_mux4_1 _21100_ (.S0(net10781),
    .A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S1(net10769),
    .X(_03520_));
 sg13g2_mux2_1 _21101_ (.A0(_03515_),
    .A1(_03520_),
    .S(net10773),
    .X(_03521_));
 sg13g2_a22oi_1 _21102_ (.Y(_03522_),
    .B1(net10262),
    .B2(_03521_),
    .A2(net10414),
    .A1(net10682));
 sg13g2_nand2_1 _21103_ (.Y(_03523_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[22] ),
    .B(net10426));
 sg13g2_o21ai_1 _21104_ (.B1(_03523_),
    .Y(_01941_),
    .A1(net10426),
    .A2(_03522_));
 sg13g2_mux4_1 _21105_ (.S0(net10855),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][23] ),
    .S1(net10794),
    .X(_03524_));
 sg13g2_mux4_1 _21106_ (.S0(net10855),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][23] ),
    .S1(net10793),
    .X(_03525_));
 sg13g2_mux4_1 _21107_ (.S0(net10855),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][23] ),
    .S1(net10794),
    .X(_03526_));
 sg13g2_mux4_1 _21108_ (.S0(net10855),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][23] ),
    .S1(net10794),
    .X(_03527_));
 sg13g2_mux4_1 _21109_ (.S0(net10775),
    .A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S1(net10764),
    .X(_03528_));
 sg13g2_mux4_1 _21110_ (.S0(net10848),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][23] ),
    .S1(net10789),
    .X(_03529_));
 sg13g2_mux4_1 _21111_ (.S0(net10848),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][23] ),
    .S1(net10789),
    .X(_03530_));
 sg13g2_mux4_1 _21112_ (.S0(net10848),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][23] ),
    .S1(net10789),
    .X(_03531_));
 sg13g2_mux4_1 _21113_ (.S0(net10848),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][23] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][23] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][23] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][23] ),
    .S1(net10789),
    .X(_03532_));
 sg13g2_mux4_1 _21114_ (.S0(net10781),
    .A0(_03529_),
    .A1(_03530_),
    .A2(_03531_),
    .A3(_03532_),
    .S1(net10769),
    .X(_03533_));
 sg13g2_mux2_1 _21115_ (.A0(_03528_),
    .A1(_03533_),
    .S(net10773),
    .X(_03534_));
 sg13g2_a221oi_1 _21116_ (.B2(_03534_),
    .C1(net10427),
    .B1(net10261),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[23] ),
    .Y(_03535_),
    .A2(net10414));
 sg13g2_a21oi_1 _21117_ (.A1(_11875_),
    .A2(net10427),
    .Y(_01942_),
    .B1(_03535_));
 sg13g2_mux4_1 _21118_ (.S0(net10856),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][24] ),
    .S1(net10794),
    .X(_03536_));
 sg13g2_mux4_1 _21119_ (.S0(net10856),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][24] ),
    .S1(net10794),
    .X(_03537_));
 sg13g2_mux4_1 _21120_ (.S0(net10849),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][24] ),
    .S1(net10791),
    .X(_03538_));
 sg13g2_mux4_1 _21121_ (.S0(net10856),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][24] ),
    .S1(net10794),
    .X(_03539_));
 sg13g2_mux4_1 _21122_ (.S0(net10781),
    .A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S1(net10764),
    .X(_03540_));
 sg13g2_mux4_1 _21123_ (.S0(net10849),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][24] ),
    .S1(net10791),
    .X(_03541_));
 sg13g2_mux4_1 _21124_ (.S0(net10849),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][24] ),
    .S1(net10791),
    .X(_03542_));
 sg13g2_mux4_1 _21125_ (.S0(net10849),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][24] ),
    .S1(net10791),
    .X(_03543_));
 sg13g2_mux4_1 _21126_ (.S0(net10849),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][24] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][24] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][24] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][24] ),
    .S1(net10791),
    .X(_03544_));
 sg13g2_mux4_1 _21127_ (.S0(net10781),
    .A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S1(net10769),
    .X(_03545_));
 sg13g2_mux2_1 _21128_ (.A0(_03540_),
    .A1(_03545_),
    .S(net10773),
    .X(_03546_));
 sg13g2_a221oi_1 _21129_ (.B2(_03546_),
    .C1(net10427),
    .B1(net10261),
    .A1(net10681),
    .Y(_03547_),
    .A2(net10414));
 sg13g2_a21oi_1 _21130_ (.A1(_08620_),
    .A2(net10427),
    .Y(_01943_),
    .B1(_03547_));
 sg13g2_buf_2 place10205 (.A(net10204),
    .X(net10205));
 sg13g2_mux4_1 _21132_ (.S0(net10859),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][25] ),
    .S1(net10797),
    .X(_03549_));
 sg13g2_mux4_1 _21133_ (.S0(net10860),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][25] ),
    .S1(net10798),
    .X(_03550_));
 sg13g2_mux4_1 _21134_ (.S0(net10860),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][25] ),
    .S1(net10798),
    .X(_03551_));
 sg13g2_buf_2 place10243 (.A(net10242),
    .X(net10243));
 sg13g2_buf_2 place10216 (.A(net10215),
    .X(net10216));
 sg13g2_mux4_1 _21137_ (.S0(net10859),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][25] ),
    .S1(net10797),
    .X(_03554_));
 sg13g2_mux4_1 _21138_ (.S0(net10776),
    .A0(_03549_),
    .A1(_03550_),
    .A2(_03551_),
    .A3(_03554_),
    .S1(net10766),
    .X(_03555_));
 sg13g2_mux4_1 _21139_ (.S0(net10865),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][25] ),
    .S1(net10803),
    .X(_03556_));
 sg13g2_mux4_1 _21140_ (.S0(net10865),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][25] ),
    .S1(net10804),
    .X(_03557_));
 sg13g2_mux4_1 _21141_ (.S0(net10866),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][25] ),
    .S1(net10805),
    .X(_03558_));
 sg13g2_mux4_1 _21142_ (.S0(net10865),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][25] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][25] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][25] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][25] ),
    .S1(net10804),
    .X(_03559_));
 sg13g2_mux4_1 _21143_ (.S0(net10775),
    .A0(_03556_),
    .A1(_03557_),
    .A2(_03558_),
    .A3(_03559_),
    .S1(net10765),
    .X(_03560_));
 sg13g2_mux2_1 _21144_ (.A0(_03555_),
    .A1(_03560_),
    .S(net10771),
    .X(_03561_));
 sg13g2_a22oi_1 _21145_ (.Y(_03562_),
    .B1(net10263),
    .B2(_03561_),
    .A2(net10415),
    .A1(net10680));
 sg13g2_nand2_1 _21146_ (.Y(_03563_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[25] ),
    .B(net10429));
 sg13g2_o21ai_1 _21147_ (.B1(_03563_),
    .Y(_01944_),
    .A1(net10429),
    .A2(_03562_));
 sg13g2_mux4_1 _21148_ (.S0(net10863),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][26] ),
    .S1(net10801),
    .X(_03564_));
 sg13g2_mux4_1 _21149_ (.S0(net10867),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][26] ),
    .S1(net10805),
    .X(_03565_));
 sg13g2_mux4_1 _21150_ (.S0(net10867),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][26] ),
    .S1(net10805),
    .X(_03566_));
 sg13g2_mux4_1 _21151_ (.S0(net10863),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][26] ),
    .S1(net10801),
    .X(_03567_));
 sg13g2_mux4_1 _21152_ (.S0(net10777),
    .A0(_03564_),
    .A1(_03565_),
    .A2(_03566_),
    .A3(_03567_),
    .S1(net10767),
    .X(_03568_));
 sg13g2_mux4_1 _21153_ (.S0(net10864),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][26] ),
    .S1(net10802),
    .X(_03569_));
 sg13g2_mux4_1 _21154_ (.S0(net10864),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][26] ),
    .S1(net10802),
    .X(_03570_));
 sg13g2_mux4_1 _21155_ (.S0(net10868),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][26] ),
    .S1(net10807),
    .X(_03571_));
 sg13g2_mux4_1 _21156_ (.S0(net10868),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][26] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][26] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][26] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][26] ),
    .S1(net10807),
    .X(_03572_));
 sg13g2_mux4_1 _21157_ (.S0(net10777),
    .A0(_03569_),
    .A1(_03570_),
    .A2(_03571_),
    .A3(_03572_),
    .S1(net10767),
    .X(_03573_));
 sg13g2_mux2_1 _21158_ (.A0(_03568_),
    .A1(_03573_),
    .S(net10774),
    .X(_03574_));
 sg13g2_a22oi_1 _21159_ (.Y(_03575_),
    .B1(net10263),
    .B2(_03574_),
    .A2(net10415),
    .A1(net10679));
 sg13g2_nand2_1 _21160_ (.Y(_03576_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[26] ),
    .B(net10428));
 sg13g2_o21ai_1 _21161_ (.B1(_03576_),
    .Y(_01945_),
    .A1(net10428),
    .A2(_03575_));
 sg13g2_mux4_1 _21162_ (.S0(net10865),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][27] ),
    .S1(net10804),
    .X(_03577_));
 sg13g2_mux4_1 _21163_ (.S0(net10865),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][27] ),
    .S1(net10804),
    .X(_03578_));
 sg13g2_mux4_1 _21164_ (.S0(net10865),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][27] ),
    .S1(net10804),
    .X(_03579_));
 sg13g2_mux4_1 _21165_ (.S0(net10865),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][27] ),
    .S1(net10804),
    .X(_03580_));
 sg13g2_mux4_1 _21166_ (.S0(net10776),
    .A0(_03577_),
    .A1(_03578_),
    .A2(_03579_),
    .A3(_03580_),
    .S1(net10766),
    .X(_03581_));
 sg13g2_mux4_1 _21167_ (.S0(net10866),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][27] ),
    .S1(net10806),
    .X(_03582_));
 sg13g2_mux4_1 _21168_ (.S0(net10866),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][27] ),
    .S1(net10806),
    .X(_03583_));
 sg13g2_mux4_1 _21169_ (.S0(net10866),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][27] ),
    .S1(net10806),
    .X(_03584_));
 sg13g2_mux4_1 _21170_ (.S0(net10866),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][27] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][27] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][27] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][27] ),
    .S1(net10806),
    .X(_03585_));
 sg13g2_mux4_1 _21171_ (.S0(net10775),
    .A0(_03582_),
    .A1(_03583_),
    .A2(_03584_),
    .A3(_03585_),
    .S1(net10765),
    .X(_03586_));
 sg13g2_mux2_1 _21172_ (.A0(_03581_),
    .A1(_03586_),
    .S(net10771),
    .X(_03587_));
 sg13g2_a22oi_1 _21173_ (.Y(_03588_),
    .B1(net10263),
    .B2(_03587_),
    .A2(net10415),
    .A1(net10678));
 sg13g2_nand2_1 _21174_ (.Y(_03589_),
    .A(net10508),
    .B(net10428));
 sg13g2_o21ai_1 _21175_ (.B1(_03589_),
    .Y(_01946_),
    .A1(net10428),
    .A2(_03588_));
 sg13g2_mux4_1 _21176_ (.S0(net10864),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][28] ),
    .S1(net10802),
    .X(_03590_));
 sg13g2_mux4_1 _21177_ (.S0(net10864),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][28] ),
    .S1(net10802),
    .X(_03591_));
 sg13g2_mux4_1 _21178_ (.S0(net10864),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][28] ),
    .S1(net10802),
    .X(_03592_));
 sg13g2_mux4_1 _21179_ (.S0(net10863),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][28] ),
    .S1(net10801),
    .X(_03593_));
 sg13g2_mux4_1 _21180_ (.S0(net10777),
    .A0(_03590_),
    .A1(_03591_),
    .A2(_03592_),
    .A3(_03593_),
    .S1(net10767),
    .X(_03594_));
 sg13g2_mux4_1 _21181_ (.S0(net10864),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][28] ),
    .S1(net10802),
    .X(_03595_));
 sg13g2_mux4_1 _21182_ (.S0(net10864),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][28] ),
    .S1(net10802),
    .X(_03596_));
 sg13g2_mux4_1 _21183_ (.S0(net10864),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][28] ),
    .S1(net10802),
    .X(_03597_));
 sg13g2_mux4_1 _21184_ (.S0(net10868),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][28] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][28] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][28] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][28] ),
    .S1(net10807),
    .X(_03598_));
 sg13g2_mux4_1 _21185_ (.S0(net10777),
    .A0(_03595_),
    .A1(_03596_),
    .A2(_03597_),
    .A3(_03598_),
    .S1(net10767),
    .X(_03599_));
 sg13g2_mux2_1 _21186_ (.A0(_03594_),
    .A1(_03599_),
    .S(net10774),
    .X(_03600_));
 sg13g2_a22oi_1 _21187_ (.Y(_03601_),
    .B1(net10263),
    .B2(_03600_),
    .A2(net10415),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[28] ));
 sg13g2_nand2_1 _21188_ (.Y(_03602_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[28] ),
    .B(net10428));
 sg13g2_o21ai_1 _21189_ (.B1(_03602_),
    .Y(_01947_),
    .A1(net10428),
    .A2(_03601_));
 sg13g2_mux4_1 _21190_ (.S0(net10859),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][29] ),
    .S1(net10797),
    .X(_03603_));
 sg13g2_mux4_1 _21191_ (.S0(net10860),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][29] ),
    .S1(net10798),
    .X(_03604_));
 sg13g2_mux4_1 _21192_ (.S0(net10860),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][29] ),
    .S1(net10798),
    .X(_03605_));
 sg13g2_mux4_1 _21193_ (.S0(net10859),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][29] ),
    .S1(net10797),
    .X(_03606_));
 sg13g2_mux4_1 _21194_ (.S0(net10776),
    .A0(_03603_),
    .A1(_03604_),
    .A2(_03605_),
    .A3(_03606_),
    .S1(net10766),
    .X(_03607_));
 sg13g2_mux4_1 _21195_ (.S0(net10860),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][29] ),
    .S1(net10798),
    .X(_03608_));
 sg13g2_mux4_1 _21196_ (.S0(net10860),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][29] ),
    .S1(net10798),
    .X(_03609_));
 sg13g2_mux4_1 _21197_ (.S0(net10860),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][29] ),
    .S1(net10798),
    .X(_03610_));
 sg13g2_mux4_1 _21198_ (.S0(net10859),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][29] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][29] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][29] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][29] ),
    .S1(net10797),
    .X(_03611_));
 sg13g2_mux4_1 _21199_ (.S0(net10776),
    .A0(_03608_),
    .A1(_03609_),
    .A2(_03610_),
    .A3(_03611_),
    .S1(net10766),
    .X(_03612_));
 sg13g2_mux2_1 _21200_ (.A0(_03607_),
    .A1(_03612_),
    .S(net10771),
    .X(_03613_));
 sg13g2_a22oi_1 _21201_ (.Y(_03614_),
    .B1(net10263),
    .B2(_03613_),
    .A2(net10415),
    .A1(net10676));
 sg13g2_nand2_1 _21202_ (.Y(_03615_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[29] ),
    .B(net10429));
 sg13g2_o21ai_1 _21203_ (.B1(_03615_),
    .Y(_01948_),
    .A1(net10429),
    .A2(_03614_));
 sg13g2_nor2_1 _21204_ (.A(net10419),
    .B(_08901_),
    .Y(_03616_));
 sg13g2_a21oi_1 _21205_ (.A1(net10675),
    .A2(net10419),
    .Y(_03617_),
    .B1(_03616_));
 sg13g2_nand2_1 _21206_ (.Y(_03618_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[2] ),
    .B(net10425));
 sg13g2_o21ai_1 _21207_ (.B1(_03618_),
    .Y(_01949_),
    .A1(net10425),
    .A2(_03617_));
 sg13g2_mux4_1 _21208_ (.S0(net10862),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][30] ),
    .S1(net10800),
    .X(_03619_));
 sg13g2_mux4_1 _21209_ (.S0(net10862),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][30] ),
    .S1(net10800),
    .X(_03620_));
 sg13g2_mux4_1 _21210_ (.S0(net10862),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][30] ),
    .S1(net10800),
    .X(_03621_));
 sg13g2_mux4_1 _21211_ (.S0(net10861),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][30] ),
    .S1(net10800),
    .X(_03622_));
 sg13g2_mux4_1 _21212_ (.S0(net10777),
    .A0(_03619_),
    .A1(_03620_),
    .A2(_03621_),
    .A3(_03622_),
    .S1(net10767),
    .X(_03623_));
 sg13g2_mux4_1 _21213_ (.S0(net10857),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][30] ),
    .S1(net10799),
    .X(_03624_));
 sg13g2_mux4_1 _21214_ (.S0(net10861),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][30] ),
    .S1(net10803),
    .X(_03625_));
 sg13g2_mux4_1 _21215_ (.S0(net10861),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][30] ),
    .S1(net10803),
    .X(_03626_));
 sg13g2_mux4_1 _21216_ (.S0(net10861),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][30] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][30] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][30] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][30] ),
    .S1(net10803),
    .X(_03627_));
 sg13g2_mux4_1 _21217_ (.S0(net10775),
    .A0(_03624_),
    .A1(_03625_),
    .A2(_03626_),
    .A3(_03627_),
    .S1(net10765),
    .X(_03628_));
 sg13g2_mux2_1 _21218_ (.A0(_03623_),
    .A1(_03628_),
    .S(net10774),
    .X(_03629_));
 sg13g2_a22oi_1 _21219_ (.Y(_03630_),
    .B1(net10263),
    .B2(_03629_),
    .A2(net10415),
    .A1(net10674));
 sg13g2_nand2_1 _21220_ (.Y(_03631_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[30] ),
    .B(net10429));
 sg13g2_o21ai_1 _21221_ (.B1(_03631_),
    .Y(_01950_),
    .A1(net10429),
    .A2(_03630_));
 sg13g2_mux4_1 _21222_ (.S0(net10862),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][31] ),
    .S1(net10800),
    .X(_03632_));
 sg13g2_mux4_1 _21223_ (.S0(net10862),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][31] ),
    .S1(net10800),
    .X(_03633_));
 sg13g2_mux4_1 _21224_ (.S0(net10862),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][31] ),
    .S1(net10800),
    .X(_03634_));
 sg13g2_mux4_1 _21225_ (.S0(net10862),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][31] ),
    .S1(net10800),
    .X(_03635_));
 sg13g2_mux4_1 _21226_ (.S0(net10777),
    .A0(_03632_),
    .A1(_03633_),
    .A2(_03634_),
    .A3(_03635_),
    .S1(net10767),
    .X(_03636_));
 sg13g2_mux4_1 _21227_ (.S0(net10857),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][31] ),
    .S1(net10795),
    .X(_03637_));
 sg13g2_mux4_1 _21228_ (.S0(net10857),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][31] ),
    .S1(net10795),
    .X(_03638_));
 sg13g2_mux4_1 _21229_ (.S0(net10845),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][31] ),
    .S1(net10795),
    .X(_03639_));
 sg13g2_mux4_1 _21230_ (.S0(net10857),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][31] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][31] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][31] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][31] ),
    .S1(net10799),
    .X(_03640_));
 sg13g2_mux4_1 _21231_ (.S0(net10776),
    .A0(_03637_),
    .A1(_03638_),
    .A2(_03639_),
    .A3(_03640_),
    .S1(net10766),
    .X(_03641_));
 sg13g2_mux2_1 _21232_ (.A0(_03636_),
    .A1(_03641_),
    .S(net10774),
    .X(_03642_));
 sg13g2_a22oi_1 _21233_ (.Y(_03643_),
    .B1(net10263),
    .B2(_03642_),
    .A2(net10415),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[31] ));
 sg13g2_nand2_1 _21234_ (.Y(_03644_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[31] ),
    .B(net10429));
 sg13g2_o21ai_1 _21235_ (.B1(_03644_),
    .Y(_01951_),
    .A1(net10428),
    .A2(_03643_));
 sg13g2_nand2_1 _21236_ (.Y(_03645_),
    .A(net10673),
    .B(net10419));
 sg13g2_o21ai_1 _21237_ (.B1(_03645_),
    .Y(_03646_),
    .A1(net10417),
    .A2(_08922_));
 sg13g2_nor2_1 _21238_ (.A(net10425),
    .B(_03646_),
    .Y(_03647_));
 sg13g2_a21oi_1 _21239_ (.A1(_08680_),
    .A2(net10425),
    .Y(_01952_),
    .B1(_03647_));
 sg13g2_nor2_1 _21240_ (.A(net10418),
    .B(_08939_),
    .Y(_03648_));
 sg13g2_a21oi_2 _21241_ (.B1(_03648_),
    .Y(_03649_),
    .A2(net10418),
    .A1(net10672));
 sg13g2_nand2_1 _21242_ (.Y(_03650_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[4] ),
    .B(net10424));
 sg13g2_o21ai_1 _21243_ (.B1(_03650_),
    .Y(_01953_),
    .A1(net10424),
    .A2(_03649_));
 sg13g2_mux4_1 _21244_ (.S0(net10832),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][5] ),
    .S1(net10809),
    .X(_03651_));
 sg13g2_mux4_1 _21245_ (.S0(net10832),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][5] ),
    .S1(net10809),
    .X(_03652_));
 sg13g2_mux4_1 _21246_ (.S0(net10832),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][5] ),
    .S1(net10809),
    .X(_03653_));
 sg13g2_mux4_1 _21247_ (.S0(net10830),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][5] ),
    .S1(net10814),
    .X(_03654_));
 sg13g2_mux4_1 _21248_ (.S0(net10780),
    .A0(_03651_),
    .A1(_03652_),
    .A2(_03653_),
    .A3(_03654_),
    .S1(net10768),
    .X(_03655_));
 sg13g2_mux4_1 _21249_ (.S0(net10842),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][5] ),
    .S1(net10824),
    .X(_03656_));
 sg13g2_mux4_1 _21250_ (.S0(net10842),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][5] ),
    .S1(net10824),
    .X(_03657_));
 sg13g2_mux4_1 _21251_ (.S0(net10842),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][5] ),
    .S1(net10824),
    .X(_03658_));
 sg13g2_mux4_1 _21252_ (.S0(net10844),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][5] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][5] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][5] ),
    .S1(net10826),
    .X(_03659_));
 sg13g2_mux4_1 _21253_ (.S0(net10780),
    .A0(_03656_),
    .A1(_03657_),
    .A2(_03658_),
    .A3(_03659_),
    .S1(net10762),
    .X(_03660_));
 sg13g2_mux2_1 _21254_ (.A0(_03655_),
    .A1(_03660_),
    .S(net10770),
    .X(_03661_));
 sg13g2_a22oi_1 _21255_ (.Y(_03662_),
    .B1(_03309_),
    .B2(_03661_),
    .A2(net10417),
    .A1(net10671));
 sg13g2_nand2_1 _21256_ (.Y(_03663_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[5] ),
    .B(net10423));
 sg13g2_o21ai_1 _21257_ (.B1(_03663_),
    .Y(_01954_),
    .A1(net10424),
    .A2(_03662_));
 sg13g2_mux4_1 _21258_ (.S0(net10837),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][6] ),
    .S1(net10819),
    .X(_03664_));
 sg13g2_mux4_1 _21259_ (.S0(net10837),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][6] ),
    .S1(net10819),
    .X(_03665_));
 sg13g2_mux4_1 _21260_ (.S0(net10837),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][6] ),
    .S1(net10819),
    .X(_03666_));
 sg13g2_mux4_1 _21261_ (.S0(net10837),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][6] ),
    .S1(net10819),
    .X(_03667_));
 sg13g2_mux4_1 _21262_ (.S0(net10783),
    .A0(_03664_),
    .A1(_03665_),
    .A2(_03666_),
    .A3(_03667_),
    .S1(net10763),
    .X(_03668_));
 sg13g2_mux4_1 _21263_ (.S0(net10837),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][6] ),
    .S1(net10819),
    .X(_03669_));
 sg13g2_mux4_1 _21264_ (.S0(net10837),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][6] ),
    .S1(net10819),
    .X(_03670_));
 sg13g2_mux4_1 _21265_ (.S0(net10837),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][6] ),
    .S1(net10819),
    .X(_03671_));
 sg13g2_mux4_1 _21266_ (.S0(net10835),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][6] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][6] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][6] ),
    .S1(net10818),
    .X(_03672_));
 sg13g2_mux4_1 _21267_ (.S0(net10783),
    .A0(_03669_),
    .A1(_03670_),
    .A2(_03671_),
    .A3(_03672_),
    .S1(net10763),
    .X(_03673_));
 sg13g2_mux2_1 _21268_ (.A0(_03668_),
    .A1(_03673_),
    .S(_00003_),
    .X(_03674_));
 sg13g2_a22oi_1 _21269_ (.Y(_03675_),
    .B1(_03309_),
    .B2(_03674_),
    .A2(net10417),
    .A1(net10670));
 sg13g2_nand2_1 _21270_ (.Y(_03676_),
    .A(net10502),
    .B(net10424));
 sg13g2_o21ai_1 _21271_ (.B1(_03676_),
    .Y(_01955_),
    .A1(net10424),
    .A2(_03675_));
 sg13g2_inv_4 _21272_ (.A(net10501),
    .Y(_03677_));
 sg13g2_mux4_1 _21273_ (.S0(net10843),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][7] ),
    .S1(net10825),
    .X(_03678_));
 sg13g2_mux4_1 _21274_ (.S0(net10843),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][7] ),
    .S1(net10825),
    .X(_03679_));
 sg13g2_mux4_1 _21275_ (.S0(net10843),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][7] ),
    .S1(net10825),
    .X(_03680_));
 sg13g2_mux4_1 _21276_ (.S0(net10843),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][7] ),
    .S1(net10825),
    .X(_03681_));
 sg13g2_mux4_1 _21277_ (.S0(net10783),
    .A0(_03678_),
    .A1(_03679_),
    .A2(_03680_),
    .A3(_03681_),
    .S1(net10763),
    .X(_03682_));
 sg13g2_mux4_1 _21278_ (.S0(net10838),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][7] ),
    .S1(net10820),
    .X(_03683_));
 sg13g2_mux4_1 _21279_ (.S0(net10838),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][7] ),
    .S1(net10820),
    .X(_03684_));
 sg13g2_mux4_1 _21280_ (.S0(net10838),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][7] ),
    .S1(net10820),
    .X(_03685_));
 sg13g2_mux4_1 _21281_ (.S0(net10839),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][7] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][7] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][7] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][7] ),
    .S1(net10821),
    .X(_03686_));
 sg13g2_mux4_1 _21282_ (.S0(net10783),
    .A0(_03683_),
    .A1(_03684_),
    .A2(_03685_),
    .A3(_03686_),
    .S1(net10763),
    .X(_03687_));
 sg13g2_mux2_1 _21283_ (.A0(_03682_),
    .A1(_03687_),
    .S(_00003_),
    .X(_03688_));
 sg13g2_a221oi_1 _21284_ (.B2(_03688_),
    .C1(net10423),
    .B1(_03309_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[7] ),
    .Y(_03689_),
    .A2(net10417));
 sg13g2_a21oi_1 _21285_ (.A1(_03677_),
    .A2(net10423),
    .Y(_01956_),
    .B1(_03689_));
 sg13g2_mux4_1 _21286_ (.S0(net10853),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][8] ),
    .S1(net10785),
    .X(_03690_));
 sg13g2_mux4_1 _21287_ (.S0(net10853),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][8] ),
    .S1(net10785),
    .X(_03691_));
 sg13g2_mux4_1 _21288_ (.S0(net10853),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][8] ),
    .S1(net10785),
    .X(_03692_));
 sg13g2_mux4_1 _21289_ (.S0(net10853),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][8] ),
    .S1(net10785),
    .X(_03693_));
 sg13g2_mux4_1 _21290_ (.S0(_00002_),
    .A0(_03690_),
    .A1(_03691_),
    .A2(_03692_),
    .A3(_03693_),
    .S1(net10764),
    .X(_03694_));
 sg13g2_mux4_1 _21291_ (.S0(net10853),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][8] ),
    .S1(net10785),
    .X(_03695_));
 sg13g2_mux4_1 _21292_ (.S0(net10853),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][8] ),
    .S1(net10785),
    .X(_03696_));
 sg13g2_mux4_1 _21293_ (.S0(net10853),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][8] ),
    .S1(net10784),
    .X(_03697_));
 sg13g2_mux4_1 _21294_ (.S0(net10853),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][8] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][8] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][8] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][8] ),
    .S1(net10785),
    .X(_03698_));
 sg13g2_mux4_1 _21295_ (.S0(_00002_),
    .A0(_03695_),
    .A1(_03696_),
    .A2(_03697_),
    .A3(_03698_),
    .S1(net10764),
    .X(_03699_));
 sg13g2_mux2_1 _21296_ (.A0(_03694_),
    .A1(_03699_),
    .S(net10774),
    .X(_03700_));
 sg13g2_a22oi_1 _21297_ (.Y(_03701_),
    .B1(_03309_),
    .B2(_03700_),
    .A2(net10416),
    .A1(net10669));
 sg13g2_nand2_1 _21298_ (.Y(_03702_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[8] ),
    .B(net10423));
 sg13g2_o21ai_1 _21299_ (.B1(_03702_),
    .Y(_01957_),
    .A1(net10423),
    .A2(_03701_));
 sg13g2_mux4_1 _21300_ (.S0(net10843),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][9] ),
    .S1(net10825),
    .X(_03703_));
 sg13g2_mux4_1 _21301_ (.S0(net10843),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][9] ),
    .S1(net10825),
    .X(_03704_));
 sg13g2_mux4_1 _21302_ (.S0(net10843),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][9] ),
    .S1(net10825),
    .X(_03705_));
 sg13g2_mux4_1 _21303_ (.S0(net10843),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][9] ),
    .S1(net10825),
    .X(_03706_));
 sg13g2_mux4_1 _21304_ (.S0(net10783),
    .A0(_03703_),
    .A1(_03704_),
    .A2(_03705_),
    .A3(_03706_),
    .S1(net10763),
    .X(_03707_));
 sg13g2_mux4_1 _21305_ (.S0(net10838),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][9] ),
    .S1(net10820),
    .X(_03708_));
 sg13g2_mux4_1 _21306_ (.S0(net10838),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][9] ),
    .S1(net10820),
    .X(_03709_));
 sg13g2_mux4_1 _21307_ (.S0(net10838),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][9] ),
    .S1(net10820),
    .X(_03710_));
 sg13g2_mux4_1 _21308_ (.S0(net10839),
    .A0(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][9] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][9] ),
    .A2(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][9] ),
    .A3(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][9] ),
    .S1(net10821),
    .X(_03711_));
 sg13g2_mux4_1 _21309_ (.S0(net10783),
    .A0(_03708_),
    .A1(_03709_),
    .A2(_03710_),
    .A3(_03711_),
    .S1(net10763),
    .X(_03712_));
 sg13g2_mux2_1 _21310_ (.A0(_03707_),
    .A1(_03712_),
    .S(_00003_),
    .X(_03713_));
 sg13g2_a221oi_1 _21311_ (.B2(_03713_),
    .C1(net10423),
    .B1(_03309_),
    .A1(net10668),
    .Y(_03714_),
    .A2(net10418));
 sg13g2_a21oi_1 _21312_ (.A1(_08779_),
    .A2(net10423),
    .Y(_01958_),
    .B1(_03714_));
 sg13g2_nand2_1 _21313_ (.Y(_03715_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_slli_srli_srai ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11] ));
 sg13g2_o21ai_1 _21314_ (.B1(_03715_),
    .Y(_03716_),
    .A1(net10632),
    .A2(_03274_));
 sg13g2_nor2_1 _21315_ (.A(net10704),
    .B(_03716_),
    .Y(_03717_));
 sg13g2_a22oi_1 _21316_ (.Y(_03718_),
    .B1(net10325),
    .B2(_08906_),
    .A2(_00109_),
    .A1(net10392));
 sg13g2_nor2_1 _21317_ (.A(_00109_),
    .B(net10325),
    .Y(_03719_));
 sg13g2_a21oi_1 _21318_ (.A1(net10392),
    .A2(_03716_),
    .Y(_03720_),
    .B1(_03719_));
 sg13g2_nand2b_1 _21319_ (.Y(_03721_),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_sh[0] ),
    .A_N(_03720_));
 sg13g2_o21ai_1 _21320_ (.B1(_03721_),
    .Y(_01990_),
    .A1(_03717_),
    .A2(_03718_));
 sg13g2_nor2_1 _21321_ (.A(net10632),
    .B(_03483_),
    .Y(_03722_));
 sg13g2_a21oi_2 _21322_ (.B1(_03722_),
    .Y(_03723_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.is_slli_srli_srai ));
 sg13g2_o21ai_1 _21323_ (.B1(net10392),
    .Y(_03724_),
    .A1(_00109_),
    .A2(net10325));
 sg13g2_nand3_1 _21324_ (.B(net10704),
    .C(net10325),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_sh[0] ),
    .Y(_03725_));
 sg13g2_nand2b_1 _21325_ (.Y(_03726_),
    .B(_03725_),
    .A_N(_03719_));
 sg13g2_a22oi_1 _21326_ (.Y(_03727_),
    .B1(_03726_),
    .B2(\u_ac_controller_soc_inst.u_picorv32.reg_sh[1] ),
    .A2(_08365_),
    .A1(net10704));
 sg13g2_o21ai_1 _21327_ (.B1(_03727_),
    .Y(_01991_),
    .A1(_03723_),
    .A2(_03724_));
 sg13g2_buf_16 clkbuf_leaf_334_clk (.X(clknet_leaf_334_clk),
    .A(clknet_8_116_0_clk));
 sg13g2_buf_2 place10161 (.A(net10160),
    .X(net10161));
 sg13g2_nor3_2 _21330_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[2] ),
    .B(_08231_),
    .C(_08259_),
    .Y(_03730_));
 sg13g2_buf_2 place10149 (.A(_04295_),
    .X(net10149));
 sg13g2_nand3b_1 _21332_ (.B(_03730_),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[0] ),
    .Y(_03732_),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[1] ));
 sg13g2_buf_2 place10150 (.A(net10149),
    .X(net10150));
 sg13g2_mux2_1 _21334_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[0] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[0] ),
    .S(_03732_),
    .X(_01993_));
 sg13g2_buf_2 place10153 (.A(net10152),
    .X(net10153));
 sg13g2_nand3b_1 _21336_ (.B(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[1] ),
    .C(_03730_),
    .Y(_03735_),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[0] ));
 sg13g2_buf_16 clkbuf_leaf_333_clk (.X(clknet_leaf_333_clk),
    .A(clknet_8_116_0_clk));
 sg13g2_mux2_1 _21338_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[2] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[10] ),
    .S(_03735_),
    .X(_01994_));
 sg13g2_buf_16 clkbuf_leaf_332_clk (.X(clknet_leaf_332_clk),
    .A(clknet_8_116_0_clk));
 sg13g2_mux2_1 _21340_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[3] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[11] ),
    .S(_03735_),
    .X(_01995_));
 sg13g2_buf_2 place10176 (.A(net10175),
    .X(net10176));
 sg13g2_mux2_1 _21342_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[4] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[12] ),
    .S(_03735_),
    .X(_01996_));
 sg13g2_buf_2 place10210 (.A(_11625_),
    .X(net10210));
 sg13g2_mux2_1 _21344_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[5] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[13] ),
    .S(_03735_),
    .X(_01997_));
 sg13g2_buf_2 place10178 (.A(net10174),
    .X(net10178));
 sg13g2_mux2_1 _21346_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[6] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[14] ),
    .S(_03735_),
    .X(_01998_));
 sg13g2_buf_16 clkbuf_leaf_335_clk (.X(clknet_leaf_335_clk),
    .A(clknet_8_116_0_clk));
 sg13g2_mux2_1 _21348_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[7] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[15] ),
    .S(_03735_),
    .X(_01999_));
 sg13g2_nand3_1 _21349_ (.B(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[1] ),
    .C(_03730_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[0] ),
    .Y(_03742_));
 sg13g2_buf_2 place10171 (.A(net10170),
    .X(net10171));
 sg13g2_mux2_1 _21351_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[0] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[16] ),
    .S(_03742_),
    .X(_02000_));
 sg13g2_buf_2 place10162 (.A(_11436_),
    .X(net10162));
 sg13g2_mux2_1 _21353_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[1] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[17] ),
    .S(_03742_),
    .X(_02001_));
 sg13g2_mux2_1 _21354_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[2] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[18] ),
    .S(_03742_),
    .X(_02002_));
 sg13g2_mux2_1 _21355_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[3] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[19] ),
    .S(_03742_),
    .X(_02003_));
 sg13g2_mux2_1 _21356_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[1] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[1] ),
    .S(_03732_),
    .X(_02004_));
 sg13g2_mux2_1 _21357_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[4] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[20] ),
    .S(_03742_),
    .X(_02005_));
 sg13g2_mux2_1 _21358_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[5] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[21] ),
    .S(_03742_),
    .X(_02006_));
 sg13g2_mux2_1 _21359_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[6] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[22] ),
    .S(_03742_),
    .X(_02007_));
 sg13g2_mux2_1 _21360_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[7] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[23] ),
    .S(_03742_),
    .X(_02008_));
 sg13g2_mux2_1 _21361_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[2] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[2] ),
    .S(_03732_),
    .X(_02009_));
 sg13g2_mux2_1 _21362_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[3] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[3] ),
    .S(_03732_),
    .X(_02010_));
 sg13g2_mux2_1 _21363_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[4] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[4] ),
    .S(_03732_),
    .X(_02011_));
 sg13g2_mux2_1 _21364_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[5] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[5] ),
    .S(_03732_),
    .X(_02012_));
 sg13g2_mux2_1 _21365_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[6] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[6] ),
    .S(_03732_),
    .X(_02013_));
 sg13g2_mux2_1 _21366_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[7] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[7] ),
    .S(_03732_),
    .X(_02014_));
 sg13g2_mux2_1 _21367_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[0] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[8] ),
    .S(_03735_),
    .X(_02015_));
 sg13g2_mux2_1 _21368_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[1] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[9] ),
    .S(_03735_),
    .X(_02016_));
 sg13g2_or3_1 _21369_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[12] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.state[5] ),
    .C(\u_ac_controller_soc_inst.u_spi_flash_mem.state[6] ),
    .X(_03745_));
 sg13g2_or3_1 _21370_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[1] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.state[9] ),
    .C(_03745_),
    .X(_03746_));
 sg13g2_buf_2 place10144 (.A(_05836_),
    .X(net10144));
 sg13g2_nor2_1 _21372_ (.A(net10469),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.state[4] ),
    .Y(_03748_));
 sg13g2_o21ai_1 _21373_ (.B1(net10470),
    .Y(_03749_),
    .A1(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[16] ),
    .A2(net9728));
 sg13g2_inv_1 _21374_ (.Y(_03750_),
    .A(_00099_));
 sg13g2_a22oi_1 _21375_ (.Y(_03751_),
    .B1(net10316),
    .B2(\u_ac_controller_soc_inst.cbus_addr[16] ),
    .A2(net10468),
    .A1(net10612));
 sg13g2_buf_2 place10157 (.A(net10156),
    .X(net10157));
 sg13g2_nand2b_1 _21377_ (.Y(_03753_),
    .B(net10297),
    .A_N(_03751_));
 sg13g2_nand4_1 _21378_ (.B(_03748_),
    .C(_03749_),
    .A(_03746_),
    .Y(_03754_),
    .D(_03753_));
 sg13g2_nand2b_2 _21379_ (.Y(_03755_),
    .B(_03748_),
    .A_N(_03746_));
 sg13g2_o21ai_1 _21380_ (.B1(_08215_),
    .Y(_03756_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[0] ),
    .A2(_03755_));
 sg13g2_nand2_2 _21381_ (.Y(_03757_),
    .A(_03750_),
    .B(_07982_));
 sg13g2_nand2b_2 _21382_ (.Y(_03758_),
    .B(_03757_),
    .A_N(_03756_));
 sg13g2_buf_2 place10202 (.A(_11808_),
    .X(net10202));
 sg13g2_buf_2 place10146 (.A(net10145),
    .X(net10146));
 sg13g2_mux2_1 _21385_ (.A0(_03754_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[0] ),
    .S(net9734),
    .X(_02035_));
 sg13g2_nand3_1 _21386_ (.B(_00098_),
    .C(net9728),
    .A(net10470),
    .Y(_03761_));
 sg13g2_nand2_1 _21387_ (.Y(_03762_),
    .A(_03755_),
    .B(_03761_));
 sg13g2_a22oi_1 _21388_ (.Y(_03763_),
    .B1(net10316),
    .B2(\u_ac_controller_soc_inst.cbus_addr[17] ),
    .A2(net10468),
    .A1(net10611));
 sg13g2_nand2_1 _21389_ (.Y(_03764_),
    .A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[22] ),
    .B(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[21] ));
 sg13g2_a21oi_1 _21390_ (.A1(net10469),
    .A2(_03764_),
    .Y(_03765_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[4] ));
 sg13g2_o21ai_1 _21391_ (.B1(_03765_),
    .Y(_03766_),
    .A1(net10302),
    .A2(_03763_));
 sg13g2_and3_1 _21392_ (.X(_03767_),
    .A(net10470),
    .B(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[17] ),
    .C(net9707));
 sg13g2_nor3_1 _21393_ (.A(_03762_),
    .B(_03766_),
    .C(_03767_),
    .Y(_03768_));
 sg13g2_nand2_1 _21394_ (.Y(_03769_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[1] ),
    .B(net9734));
 sg13g2_o21ai_1 _21395_ (.B1(_03769_),
    .Y(_02036_),
    .A1(net9734),
    .A2(_03768_));
 sg13g2_and2_1 _21396_ (.A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[22] ),
    .B(net10469),
    .X(_03770_));
 sg13g2_a22oi_1 _21397_ (.Y(_03771_),
    .B1(_03770_),
    .B2(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[21] ),
    .A2(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[18] ),
    .A1(net10470));
 sg13g2_a22oi_1 _21398_ (.Y(_03772_),
    .B1(net10316),
    .B2(\u_ac_controller_soc_inst.cbus_addr[18] ),
    .A2(net10468),
    .A1(\u_ac_controller_soc_inst.cbus_addr[10] ));
 sg13g2_nand2b_1 _21399_ (.Y(_03773_),
    .B(net10298),
    .A_N(_03772_));
 sg13g2_and3_1 _21400_ (.X(_03774_),
    .A(net10621),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.state[12] ),
    .C(net10297));
 sg13g2_o21ai_1 _21401_ (.B1(net9728),
    .Y(_03775_),
    .A1(net10470),
    .A2(_03774_));
 sg13g2_nand4_1 _21402_ (.B(_03771_),
    .C(_03773_),
    .A(_03755_),
    .Y(_03776_),
    .D(_03775_));
 sg13g2_mux2_1 _21403_ (.A0(_03776_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[2] ),
    .S(net9734),
    .X(_02037_));
 sg13g2_inv_1 _21404_ (.Y(_03777_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[3] ));
 sg13g2_buf_2 place10170 (.A(_10095_),
    .X(net10170));
 sg13g2_a22oi_1 _21406_ (.Y(_03779_),
    .B1(net10316),
    .B2(\u_ac_controller_soc_inst.cbus_addr[19] ),
    .A2(net10468),
    .A1(net10626));
 sg13g2_nand2_1 _21407_ (.Y(_03780_),
    .A(net10469),
    .B(_08226_));
 sg13g2_o21ai_1 _21408_ (.B1(_03780_),
    .Y(_03781_),
    .A1(net10469),
    .A2(_03746_));
 sg13g2_nor2_1 _21409_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[4] ),
    .B(_03781_),
    .Y(_03782_));
 sg13g2_o21ai_1 _21410_ (.B1(_03782_),
    .Y(_03783_),
    .A1(net10302),
    .A2(_03779_));
 sg13g2_nand3_1 _21411_ (.B(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[19] ),
    .C(net9707),
    .A(net10470),
    .Y(_03784_));
 sg13g2_nand4_1 _21412_ (.B(\u_ac_controller_soc_inst.u_spi_flash_mem.state[12] ),
    .C(net10298),
    .A(net10619),
    .Y(_03785_),
    .D(net9728));
 sg13g2_nand3_1 _21413_ (.B(_03784_),
    .C(_03785_),
    .A(_03761_),
    .Y(_03786_));
 sg13g2_nor3_2 _21414_ (.A(_03758_),
    .B(_03783_),
    .C(_03786_),
    .Y(_03787_));
 sg13g2_a21oi_1 _21415_ (.A1(_03777_),
    .A2(net9734),
    .Y(_02038_),
    .B1(_03787_));
 sg13g2_and3_2 _21416_ (.X(_03788_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[12] ),
    .B(net10297),
    .C(net9728));
 sg13g2_buf_2 place10206 (.A(net10203),
    .X(net10206));
 sg13g2_a22oi_1 _21418_ (.Y(_03790_),
    .B1(net10316),
    .B2(net10624),
    .A2(net10468),
    .A1(\u_ac_controller_soc_inst.cbus_addr[12] ));
 sg13g2_nor2_1 _21419_ (.A(net10301),
    .B(_03790_),
    .Y(_03791_));
 sg13g2_a221oi_1 _21420_ (.B2(\u_ac_controller_soc_inst.cbus_addr[4] ),
    .C1(_03791_),
    .B1(_03788_),
    .A1(_08264_),
    .Y(_03792_),
    .A2(_03770_));
 sg13g2_nor2b_1 _21421_ (.A(_03762_),
    .B_N(_03792_),
    .Y(_03793_));
 sg13g2_nand2_1 _21422_ (.Y(_03794_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[4] ),
    .B(_03758_));
 sg13g2_o21ai_1 _21423_ (.B1(_03794_),
    .Y(_02039_),
    .A1(net9734),
    .A2(_03793_));
 sg13g2_a22oi_1 _21424_ (.Y(_03795_),
    .B1(net10316),
    .B2(net10623),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.state[6] ),
    .A1(net10625));
 sg13g2_and2_1 _21425_ (.A(_08217_),
    .B(_03782_),
    .X(_03796_));
 sg13g2_o21ai_1 _21426_ (.B1(_03796_),
    .Y(_03797_),
    .A1(net10302),
    .A2(_03795_));
 sg13g2_a21oi_2 _21427_ (.B1(_03797_),
    .Y(_03798_),
    .A2(_03788_),
    .A1(net10616));
 sg13g2_nand2_1 _21428_ (.Y(_03799_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[5] ),
    .B(net9734));
 sg13g2_o21ai_1 _21429_ (.B1(_03799_),
    .Y(_02040_),
    .A1(net9734),
    .A2(_03798_));
 sg13g2_a22oi_1 _21430_ (.Y(_03800_),
    .B1(net10316),
    .B2(\u_ac_controller_soc_inst.cbus_addr[22] ),
    .A2(net10468),
    .A1(\u_ac_controller_soc_inst.cbus_addr[14] ));
 sg13g2_nor2_1 _21431_ (.A(net10301),
    .B(_03800_),
    .Y(_03801_));
 sg13g2_a221oi_1 _21432_ (.B2(net10614),
    .C1(_03801_),
    .B1(_03788_),
    .A1(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[21] ),
    .Y(_03802_),
    .A2(net10469));
 sg13g2_nor2b_1 _21433_ (.A(_03762_),
    .B_N(_03802_),
    .Y(_03803_));
 sg13g2_nand2_1 _21434_ (.Y(_03804_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[6] ),
    .B(_03758_));
 sg13g2_o21ai_1 _21435_ (.B1(_03804_),
    .Y(_02041_),
    .A1(_03758_),
    .A2(_03803_));
 sg13g2_a22oi_1 _21436_ (.Y(_03805_),
    .B1(net10316),
    .B2(net10622),
    .A2(net10468),
    .A1(\u_ac_controller_soc_inst.cbus_addr[15] ));
 sg13g2_o21ai_1 _21437_ (.B1(_03796_),
    .Y(_03806_),
    .A1(net10302),
    .A2(_03805_));
 sg13g2_a21oi_2 _21438_ (.B1(_03806_),
    .Y(_03807_),
    .A2(_03788_),
    .A1(net10613));
 sg13g2_nand2_1 _21439_ (.Y(_03808_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[7] ),
    .B(_03758_));
 sg13g2_o21ai_1 _21440_ (.B1(_03808_),
    .Y(_02042_),
    .A1(_03758_),
    .A2(_03807_));
 sg13g2_nor2_1 _21441_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[0] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[1] ),
    .Y(_03809_));
 sg13g2_nand3_1 _21442_ (.B(_08240_),
    .C(_03809_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[2] ),
    .Y(_03810_));
 sg13g2_buf_2 place10145 (.A(_05836_),
    .X(net10145));
 sg13g2_nor2_2 _21444_ (.A(_08231_),
    .B(_03810_),
    .Y(_03812_));
 sg13g2_buf_16 clkbuf_leaf_337_clk (.X(clknet_leaf_337_clk),
    .A(clknet_8_94_0_clk));
 sg13g2_buf_16 clkbuf_leaf_336_clk (.X(clknet_leaf_336_clk),
    .A(clknet_8_113_0_clk));
 sg13g2_buf_2 place10137 (.A(net10134),
    .X(net10137));
 sg13g2_inv_4 _21448_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_inc ),
    .Y(_03816_));
 sg13g2_buf_2 place10136 (.A(net10134),
    .X(net10136));
 sg13g2_buf_2 place10135 (.A(net10134),
    .X(net10135));
 sg13g2_mux2_1 _21451_ (.A0(_08031_),
    .A1(_08108_),
    .S(net10312),
    .X(_03819_));
 sg13g2_buf_2 place10421 (.A(net10420),
    .X(net10421));
 sg13g2_o21ai_1 _21453_ (.B1(net9663),
    .Y(_03821_),
    .A1(net10312),
    .A2(_08105_));
 sg13g2_a22oi_1 _21454_ (.Y(_02050_),
    .B1(_03821_),
    .B2(_07788_),
    .A2(_03819_),
    .A1(net9663));
 sg13g2_or2_1 _21455_ (.X(_03822_),
    .B(_03810_),
    .A(_08231_));
 sg13g2_buf_2 place10165 (.A(_11413_),
    .X(net10165));
 sg13g2_buf_2 place10152 (.A(_04295_),
    .X(net10152));
 sg13g2_buf_2 place10134 (.A(_09852_),
    .X(net10134));
 sg13g2_nor2_2 _21459_ (.A(net10471),
    .B(net10300),
    .Y(_03826_));
 sg13g2_buf_2 place10151 (.A(net10150),
    .X(net10151));
 sg13g2_buf_2 place10169 (.A(net10168),
    .X(net10169));
 sg13g2_nor2_1 _21462_ (.A(net10484),
    .B(net10311),
    .Y(_03829_));
 sg13g2_a22oi_1 _21463_ (.Y(_03830_),
    .B1(_03829_),
    .B2(net10291),
    .A2(_03826_),
    .A1(net10626));
 sg13g2_buf_16 clkbuf_leaf_340_clk (.X(clknet_leaf_340_clk),
    .A(clknet_8_117_0_clk));
 sg13g2_buf_16 clkbuf_leaf_338_clk (.X(clknet_leaf_338_clk),
    .A(clknet_8_95_0_clk));
 sg13g2_nor2_1 _21466_ (.A(net10311),
    .B(net10291),
    .Y(_03833_));
 sg13g2_o21ai_1 _21467_ (.B1(net10484),
    .Y(_03834_),
    .A1(net9655),
    .A2(_03833_));
 sg13g2_o21ai_1 _21468_ (.B1(_03834_),
    .Y(_02051_),
    .A1(net9655),
    .A2(_03830_));
 sg13g2_o21ai_1 _21469_ (.B1(net10312),
    .Y(_03835_),
    .A1(_07739_),
    .A2(net10300));
 sg13g2_o21ai_1 _21470_ (.B1(_03835_),
    .Y(_03836_),
    .A1(net10311),
    .A2(_08033_));
 sg13g2_a21o_1 _21471_ (.A2(net10291),
    .A1(net10484),
    .B1(net10311),
    .X(_03837_));
 sg13g2_a21oi_1 _21472_ (.A1(net9663),
    .A2(_03837_),
    .Y(_03838_),
    .B1(net10483));
 sg13g2_a21oi_1 _21473_ (.A1(net9663),
    .A2(_03836_),
    .Y(_02052_),
    .B1(_03838_));
 sg13g2_nor3_1 _21474_ (.A(net10482),
    .B(net10311),
    .C(_08033_),
    .Y(_03839_));
 sg13g2_a21oi_1 _21475_ (.A1(net10625),
    .A2(_03826_),
    .Y(_03840_),
    .B1(_03839_));
 sg13g2_and2_1 _21476_ (.A(net10471),
    .B(_08033_),
    .X(_03841_));
 sg13g2_o21ai_1 _21477_ (.B1(net10482),
    .Y(_03842_),
    .A1(net9655),
    .A2(_03841_));
 sg13g2_o21ai_1 _21478_ (.B1(_03842_),
    .Y(_02053_),
    .A1(net9655),
    .A2(_03840_));
 sg13g2_buf_2 place10133 (.A(net10132),
    .X(net10133));
 sg13g2_mux2_1 _21480_ (.A0(_07729_),
    .A1(_08018_),
    .S(net10472),
    .X(_03844_));
 sg13g2_nand2_1 _21481_ (.Y(_03845_),
    .A(net10472),
    .B(_08106_));
 sg13g2_a21oi_1 _21482_ (.A1(net9664),
    .A2(_03845_),
    .Y(_03846_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[14] ));
 sg13g2_a21oi_1 _21483_ (.A1(net9664),
    .A2(_03844_),
    .Y(_02054_),
    .B1(_03846_));
 sg13g2_nor2_1 _21484_ (.A(net10472),
    .B(_08045_),
    .Y(_03847_));
 sg13g2_a21oi_1 _21485_ (.A1(net10472),
    .A2(_08019_),
    .Y(_03848_),
    .B1(_03847_));
 sg13g2_o21ai_1 _21486_ (.B1(net9664),
    .Y(_03849_),
    .A1(net10312),
    .A2(_08018_));
 sg13g2_a22oi_1 _21487_ (.Y(_02055_),
    .B1(_03849_),
    .B2(_08029_),
    .A2(_03848_),
    .A1(net9664));
 sg13g2_nor2_1 _21488_ (.A(net10472),
    .B(_07727_),
    .Y(_03850_));
 sg13g2_a21oi_1 _21489_ (.A1(net10472),
    .A2(_08020_),
    .Y(_03851_),
    .B1(_03850_));
 sg13g2_nand2_1 _21490_ (.Y(_03852_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[16] ),
    .B(net9657));
 sg13g2_o21ai_1 _21491_ (.B1(_03852_),
    .Y(_02056_),
    .A1(net9657),
    .A2(_03851_));
 sg13g2_mux2_1 _21492_ (.A0(_07998_),
    .A1(_08098_),
    .S(net10312),
    .X(_03853_));
 sg13g2_o21ai_1 _21493_ (.B1(net9664),
    .Y(_03854_),
    .A1(net10312),
    .A2(_08006_));
 sg13g2_a22oi_1 _21494_ (.Y(_02057_),
    .B1(_03854_),
    .B2(_07986_),
    .A2(_03853_),
    .A1(net9664));
 sg13g2_nor2_1 _21495_ (.A(_07760_),
    .B(net10300),
    .Y(_03855_));
 sg13g2_nand3_1 _21496_ (.B(net10472),
    .C(_07998_),
    .A(net10481),
    .Y(_03856_));
 sg13g2_o21ai_1 _21497_ (.B1(_03856_),
    .Y(_03857_),
    .A1(net10472),
    .A2(_03855_));
 sg13g2_o21ai_1 _21498_ (.B1(net9664),
    .Y(_03858_),
    .A1(net10312),
    .A2(_08007_));
 sg13g2_a22oi_1 _21499_ (.Y(_02058_),
    .B1(_03858_),
    .B2(_08096_),
    .A2(_03857_),
    .A1(net9664));
 sg13g2_mux2_1 _21500_ (.A0(_08116_),
    .A1(_08100_),
    .S(net10313),
    .X(_03859_));
 sg13g2_a21o_1 _21501_ (.A2(_07998_),
    .A1(net10481),
    .B1(net10312),
    .X(_03860_));
 sg13g2_a21oi_1 _21502_ (.A1(net9663),
    .A2(_03860_),
    .Y(_03861_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19] ));
 sg13g2_a21oi_1 _21503_ (.A1(net9663),
    .A2(_03859_),
    .Y(_02059_),
    .B1(_03861_));
 sg13g2_nor2_1 _21504_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20] ),
    .B(net10313),
    .Y(_03862_));
 sg13g2_a22oi_1 _21505_ (.Y(_03863_),
    .B1(_03862_),
    .B2(_08116_),
    .A2(_03826_),
    .A1(net10624));
 sg13g2_nor2_1 _21506_ (.A(net10313),
    .B(_08116_),
    .Y(_03864_));
 sg13g2_o21ai_1 _21507_ (.B1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20] ),
    .Y(_03865_),
    .A1(net9657),
    .A2(_03864_));
 sg13g2_o21ai_1 _21508_ (.B1(_03865_),
    .Y(_02060_),
    .A1(net9657),
    .A2(_03863_));
 sg13g2_nor2_1 _21509_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21] ),
    .B(net10315),
    .Y(_03866_));
 sg13g2_a22oi_1 _21510_ (.Y(_03867_),
    .B1(_03866_),
    .B2(_08000_),
    .A2(net10197),
    .A1(net10623));
 sg13g2_nor2_1 _21511_ (.A(net10314),
    .B(_08000_),
    .Y(_03868_));
 sg13g2_o21ai_1 _21512_ (.B1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21] ),
    .Y(_03869_),
    .A1(net9656),
    .A2(_03868_));
 sg13g2_o21ai_1 _21513_ (.B1(_03869_),
    .Y(_02061_),
    .A1(net9656),
    .A2(_03867_));
 sg13g2_nor2_1 _21514_ (.A(net10480),
    .B(net10315),
    .Y(_03870_));
 sg13g2_a22oi_1 _21515_ (.Y(_03871_),
    .B1(_03870_),
    .B2(_08002_),
    .A2(_03826_),
    .A1(\u_ac_controller_soc_inst.cbus_addr[22] ));
 sg13g2_nor2_1 _21516_ (.A(net10315),
    .B(_08002_),
    .Y(_03872_));
 sg13g2_o21ai_1 _21517_ (.B1(net10480),
    .Y(_03873_),
    .A1(net9657),
    .A2(_03872_));
 sg13g2_o21ai_1 _21518_ (.B1(_03873_),
    .Y(_02062_),
    .A1(net9657),
    .A2(_03871_));
 sg13g2_nand2_1 _21519_ (.Y(_03874_),
    .A(net10480),
    .B(_08002_));
 sg13g2_nor3_1 _21520_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23] ),
    .B(net10315),
    .C(_03874_),
    .Y(_03875_));
 sg13g2_a21oi_1 _21521_ (.A1(net10622),
    .A2(_03826_),
    .Y(_03876_),
    .B1(_03875_));
 sg13g2_a21oi_1 _21522_ (.A1(net10471),
    .A2(_03874_),
    .Y(_03877_),
    .B1(net9657));
 sg13g2_nand2b_1 _21523_ (.Y(_03878_),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23] ),
    .A_N(_03877_));
 sg13g2_o21ai_1 _21524_ (.B1(_03878_),
    .Y(_02063_),
    .A1(net9657),
    .A2(_03876_));
 sg13g2_nor2_1 _21525_ (.A(_08082_),
    .B(net10471),
    .Y(_03879_));
 sg13g2_a22oi_1 _21526_ (.Y(_03880_),
    .B1(net10297),
    .B2(_03879_),
    .A2(net10471),
    .A1(_00125_));
 sg13g2_nand2_1 _21527_ (.Y(_03881_),
    .A(net10479),
    .B(net9654));
 sg13g2_o21ai_1 _21528_ (.B1(_03881_),
    .Y(_02064_),
    .A1(net9654),
    .A2(_03880_));
 sg13g2_nor2b_1 _21529_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[3] ),
    .B_N(net10479),
    .Y(_03882_));
 sg13g2_a22oi_1 _21530_ (.Y(_03883_),
    .B1(net10197),
    .B2(net10619),
    .A2(_03882_),
    .A1(net10471));
 sg13g2_nor2_1 _21531_ (.A(net10479),
    .B(net10311),
    .Y(_03884_));
 sg13g2_o21ai_1 _21532_ (.B1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[3] ),
    .Y(_03885_),
    .A1(net9655),
    .A2(_03884_));
 sg13g2_o21ai_1 _21533_ (.B1(_03885_),
    .Y(_02065_),
    .A1(net9654),
    .A2(_03883_));
 sg13g2_o21ai_1 _21534_ (.B1(net10313),
    .Y(_03886_),
    .A1(_07707_),
    .A2(net10301));
 sg13g2_o21ai_1 _21535_ (.B1(_03886_),
    .Y(_03887_),
    .A1(net10313),
    .A2(_07990_));
 sg13g2_nand2_1 _21536_ (.Y(_03888_),
    .A(net10471),
    .B(_08123_));
 sg13g2_a21oi_1 _21537_ (.A1(_03812_),
    .A2(_03888_),
    .Y(_03889_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[4] ));
 sg13g2_a21oi_1 _21538_ (.A1(net9663),
    .A2(_03887_),
    .Y(_02066_),
    .B1(_03889_));
 sg13g2_buf_2 place10132 (.A(net10130),
    .X(net10132));
 sg13g2_nor2_1 _21540_ (.A(net10476),
    .B(net10314),
    .Y(_03891_));
 sg13g2_a22oi_1 _21541_ (.Y(_03892_),
    .B1(_03891_),
    .B2(_08064_),
    .A2(net10197),
    .A1(net10616));
 sg13g2_nor2_1 _21542_ (.A(net10314),
    .B(_08064_),
    .Y(_03893_));
 sg13g2_o21ai_1 _21543_ (.B1(net10476),
    .Y(_03894_),
    .A1(_03822_),
    .A2(_03893_));
 sg13g2_o21ai_1 _21544_ (.B1(_03894_),
    .Y(_02067_),
    .A1(_03822_),
    .A2(_03892_));
 sg13g2_nor3_1 _21545_ (.A(net10475),
    .B(net10314),
    .C(_08075_),
    .Y(_03895_));
 sg13g2_a21oi_1 _21546_ (.A1(net10614),
    .A2(net10197),
    .Y(_03896_),
    .B1(_03895_));
 sg13g2_a21oi_1 _21547_ (.A1(net10476),
    .A2(_08064_),
    .Y(_03897_),
    .B1(net10314));
 sg13g2_o21ai_1 _21548_ (.B1(net10475),
    .Y(_03898_),
    .A1(_03822_),
    .A2(_03897_));
 sg13g2_o21ai_1 _21549_ (.B1(_03898_),
    .Y(_02068_),
    .A1(net9656),
    .A2(_03896_));
 sg13g2_nor2_1 _21550_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[7] ),
    .B(_03816_),
    .Y(_03899_));
 sg13g2_a22oi_1 _21551_ (.Y(_03900_),
    .B1(_03899_),
    .B2(_08066_),
    .A2(net10197),
    .A1(net10613));
 sg13g2_nor2_1 _21552_ (.A(_03816_),
    .B(_08066_),
    .Y(_03901_));
 sg13g2_o21ai_1 _21553_ (.B1(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[7] ),
    .Y(_03902_),
    .A1(net9654),
    .A2(_03901_));
 sg13g2_o21ai_1 _21554_ (.B1(_03902_),
    .Y(_02069_),
    .A1(net9654),
    .A2(_03900_));
 sg13g2_nor2_1 _21555_ (.A(net10474),
    .B(net10315),
    .Y(_03903_));
 sg13g2_a22oi_1 _21556_ (.Y(_03904_),
    .B1(_03903_),
    .B2(_07994_),
    .A2(net10197),
    .A1(net10612));
 sg13g2_nor2_1 _21557_ (.A(net10315),
    .B(_07994_),
    .Y(_03905_));
 sg13g2_o21ai_1 _21558_ (.B1(net10474),
    .Y(_03906_),
    .A1(net9658),
    .A2(_03905_));
 sg13g2_o21ai_1 _21559_ (.B1(_03906_),
    .Y(_02070_),
    .A1(net9656),
    .A2(_03904_));
 sg13g2_nor3_1 _21560_ (.A(net10473),
    .B(net10315),
    .C(_08142_),
    .Y(_03907_));
 sg13g2_a21oi_1 _21561_ (.A1(\u_ac_controller_soc_inst.cbus_addr[9] ),
    .A2(net10197),
    .Y(_03908_),
    .B1(_03907_));
 sg13g2_a21oi_1 _21562_ (.A1(net10474),
    .A2(_07994_),
    .Y(_03909_),
    .B1(net10315));
 sg13g2_o21ai_1 _21563_ (.B1(net10473),
    .Y(_03910_),
    .A1(net9659),
    .A2(_03909_));
 sg13g2_o21ai_1 _21564_ (.B1(_03910_),
    .Y(_02071_),
    .A1(net9659),
    .A2(_03908_));
 sg13g2_or2_1 _21565_ (.X(_03911_),
    .B(_08151_),
    .A(net10469));
 sg13g2_a22oi_1 _21566_ (.Y(_02072_),
    .B1(_03911_),
    .B2(_08215_),
    .A2(_03822_),
    .A1(_03816_));
 sg13g2_inv_1 _21567_ (.Y(_03912_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_wait ));
 sg13g2_a21oi_1 _21568_ (.A1(_07744_),
    .A2(_03810_),
    .Y(_03913_),
    .B1(_08231_));
 sg13g2_nand3_1 _21569_ (.B(_07744_),
    .C(_03812_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_inc ),
    .Y(_03914_));
 sg13g2_o21ai_1 _21570_ (.B1(_03914_),
    .Y(_02074_),
    .A1(_03912_),
    .A2(_03913_));
 sg13g2_mux2_1 _21571_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[0] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[0] ),
    .S(net9659),
    .X(_02075_));
 sg13g2_mux2_1 _21572_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[10] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[10] ),
    .S(net9660),
    .X(_02076_));
 sg13g2_mux2_1 _21573_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[11] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[11] ),
    .S(net9660),
    .X(_02077_));
 sg13g2_mux2_1 _21574_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[12] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[12] ),
    .S(net9660),
    .X(_02078_));
 sg13g2_mux2_1 _21575_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[13] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[13] ),
    .S(net9660),
    .X(_02079_));
 sg13g2_buf_2 place10148 (.A(net10147),
    .X(net10148));
 sg13g2_mux2_1 _21577_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[14] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[14] ),
    .S(net9661),
    .X(_02080_));
 sg13g2_mux2_1 _21578_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[15] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[15] ),
    .S(net9662),
    .X(_02081_));
 sg13g2_mux2_1 _21579_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[16] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[16] ),
    .S(net9658),
    .X(_02082_));
 sg13g2_mux2_1 _21580_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[17] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[17] ),
    .S(net9662),
    .X(_02083_));
 sg13g2_mux2_1 _21581_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[18] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[18] ),
    .S(net9662),
    .X(_02084_));
 sg13g2_mux2_1 _21582_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[19] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[19] ),
    .S(net9662),
    .X(_02085_));
 sg13g2_mux2_1 _21583_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[1] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[1] ),
    .S(net9659),
    .X(_02086_));
 sg13g2_mux2_1 _21584_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[20] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[20] ),
    .S(net9661),
    .X(_02087_));
 sg13g2_mux2_1 _21585_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[21] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[21] ),
    .S(net9659),
    .X(_02088_));
 sg13g2_mux2_1 _21586_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[22] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[22] ),
    .S(net9662),
    .X(_02089_));
 sg13g2_buf_2 place10131 (.A(net10130),
    .X(net10131));
 sg13g2_mux2_1 _21588_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[23] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[23] ),
    .S(net9662),
    .X(_02090_));
 sg13g2_mux2_1 _21589_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[0] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[24] ),
    .S(net9659),
    .X(_02091_));
 sg13g2_mux2_1 _21590_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[1] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[25] ),
    .S(net9659),
    .X(_02092_));
 sg13g2_mux2_1 _21591_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[2] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[26] ),
    .S(net9661),
    .X(_02093_));
 sg13g2_mux2_1 _21592_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[3] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[27] ),
    .S(net9662),
    .X(_02094_));
 sg13g2_mux2_1 _21593_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[4] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[28] ),
    .S(net9661),
    .X(_02095_));
 sg13g2_mux2_1 _21594_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[5] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[29] ),
    .S(net9659),
    .X(_02096_));
 sg13g2_nand2_1 _21595_ (.Y(_03917_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[2] ),
    .B(_03812_));
 sg13g2_o21ai_1 _21596_ (.B1(_03917_),
    .Y(_02097_),
    .A1(_08431_),
    .A2(_03812_));
 sg13g2_mux2_1 _21597_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[6] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[30] ),
    .S(net9660),
    .X(_02098_));
 sg13g2_mux2_1 _21598_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[7] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[31] ),
    .S(net9661),
    .X(_02099_));
 sg13g2_nand2_1 _21599_ (.Y(_03918_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[3] ),
    .B(_03812_));
 sg13g2_o21ai_1 _21600_ (.B1(_03918_),
    .Y(_02100_),
    .A1(_08436_),
    .A2(_03812_));
 sg13g2_mux2_1 _21601_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[4] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[4] ),
    .S(net9658),
    .X(_02101_));
 sg13g2_mux2_1 _21602_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[5] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[5] ),
    .S(net9660),
    .X(_02102_));
 sg13g2_mux2_1 _21603_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[6] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[6] ),
    .S(net9658),
    .X(_02103_));
 sg13g2_mux2_1 _21604_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[7] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[7] ),
    .S(net9660),
    .X(_02104_));
 sg13g2_mux2_1 _21605_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[8] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[8] ),
    .S(net9658),
    .X(_02105_));
 sg13g2_mux2_1 _21606_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[9] ),
    .A1(\u_ac_controller_soc_inst.spi_flash_rdata[9] ),
    .S(net9660),
    .X(_02106_));
 sg13g2_and2_1 _21607_ (.A(_08171_),
    .B(_08571_),
    .X(_03919_));
 sg13g2_o21ai_1 _21608_ (.B1(_08180_),
    .Y(_03920_),
    .A1(net10466),
    .A2(_00090_));
 sg13g2_o21ai_1 _21609_ (.B1(_03920_),
    .Y(_03921_),
    .A1(net10467),
    .A2(_08180_));
 sg13g2_nand3_1 _21610_ (.B(_03919_),
    .C(_03921_),
    .A(net10461),
    .Y(_03922_));
 sg13g2_buf_2 place10138 (.A(net10137),
    .X(net10138));
 sg13g2_buf_2 place10155 (.A(net10154),
    .X(net10155));
 sg13g2_buf_2 place10154 (.A(net10153),
    .X(net10154));
 sg13g2_buf_2 place10156 (.A(net10152),
    .X(net10156));
 sg13g2_nor2b_1 _21615_ (.A(_08197_),
    .B_N(spi_flash_io0_di),
    .Y(_03927_));
 sg13g2_a21oi_1 _21616_ (.A1(spi_flash_io1_di),
    .A2(net10457),
    .Y(_03928_),
    .B1(_03927_));
 sg13g2_nand2_1 _21617_ (.Y(_03929_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[0] ),
    .B(_03922_));
 sg13g2_o21ai_1 _21618_ (.B1(_03929_),
    .Y(_02119_),
    .A1(_03922_),
    .A2(_03928_));
 sg13g2_nor2b_1 _21619_ (.A(net10457),
    .B_N(spi_flash_io1_di),
    .Y(_03930_));
 sg13g2_a21oi_1 _21620_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[0] ),
    .A2(net10457),
    .Y(_03931_),
    .B1(_03930_));
 sg13g2_nand2_1 _21621_ (.Y(_03932_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[1] ),
    .B(net10160));
 sg13g2_o21ai_1 _21622_ (.B1(_03932_),
    .Y(_02120_),
    .A1(net10160),
    .A2(_03931_));
 sg13g2_nor2_2 _21623_ (.A(net10462),
    .B(net10456),
    .Y(_03933_));
 sg13g2_buf_2 place10130 (.A(_09868_),
    .X(net10130));
 sg13g2_buf_16 clkbuf_leaf_342_clk (.X(clknet_leaf_342_clk),
    .A(clknet_8_94_0_clk));
 sg13g2_and2_1 _21626_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[1] ),
    .B(net10458),
    .X(_03936_));
 sg13g2_a221oi_1 _21627_ (.B2(_03933_),
    .C1(_03936_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[0] ),
    .A1(net10463),
    .Y(_03937_),
    .A2(spi_flash_io2_di));
 sg13g2_nand2_1 _21628_ (.Y(_03938_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[2] ),
    .B(net10160));
 sg13g2_o21ai_1 _21629_ (.B1(_03938_),
    .Y(_02121_),
    .A1(net10160),
    .A2(_03937_));
 sg13g2_and2_1 _21630_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[2] ),
    .B(net10458),
    .X(_03939_));
 sg13g2_a221oi_1 _21631_ (.B2(_03933_),
    .C1(_03939_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[1] ),
    .A1(net10463),
    .Y(_03940_),
    .A2(spi_flash_io3_di));
 sg13g2_nand2_1 _21632_ (.Y(_03941_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[3] ),
    .B(net10160));
 sg13g2_o21ai_1 _21633_ (.B1(_03941_),
    .Y(_02122_),
    .A1(net10160),
    .A2(_03940_));
 sg13g2_and2_1 _21634_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[3] ),
    .B(net10458),
    .X(_03942_));
 sg13g2_a221oi_1 _21635_ (.B2(_03933_),
    .C1(_03942_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[2] ),
    .A1(net10463),
    .Y(_03943_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[0] ));
 sg13g2_nand2_1 _21636_ (.Y(_03944_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[4] ),
    .B(net10161));
 sg13g2_o21ai_1 _21637_ (.B1(_03944_),
    .Y(_02123_),
    .A1(net10161),
    .A2(_03943_));
 sg13g2_and2_1 _21638_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[4] ),
    .B(net10458),
    .X(_03945_));
 sg13g2_a221oi_1 _21639_ (.B2(_03933_),
    .C1(_03945_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[3] ),
    .A1(net10463),
    .Y(_03946_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[1] ));
 sg13g2_nand2_1 _21640_ (.Y(_03947_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[5] ),
    .B(net10161));
 sg13g2_o21ai_1 _21641_ (.B1(_03947_),
    .Y(_02124_),
    .A1(net10161),
    .A2(_03946_));
 sg13g2_and2_1 _21642_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[5] ),
    .B(net10458),
    .X(_03948_));
 sg13g2_a221oi_1 _21643_ (.B2(_03933_),
    .C1(_03948_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[4] ),
    .A1(net10463),
    .Y(_03949_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[2] ));
 sg13g2_nand2_1 _21644_ (.Y(_03950_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[6] ),
    .B(net10161));
 sg13g2_o21ai_1 _21645_ (.B1(_03950_),
    .Y(_02125_),
    .A1(net10161),
    .A2(_03949_));
 sg13g2_and2_1 _21646_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[6] ),
    .B(net10458),
    .X(_03951_));
 sg13g2_a221oi_1 _21647_ (.B2(_03933_),
    .C1(_03951_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[5] ),
    .A1(net10463),
    .Y(_03952_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[3] ));
 sg13g2_nand2_1 _21648_ (.Y(_03953_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[7] ),
    .B(net10161));
 sg13g2_o21ai_1 _21649_ (.B1(_03953_),
    .Y(_02126_),
    .A1(net10161),
    .A2(_03952_));
 sg13g2_inv_1 _21650_ (.Y(_03954_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[0] ));
 sg13g2_nand3b_1 _21651_ (.B(_00090_),
    .C(_08180_),
    .Y(_03955_),
    .A_N(net10466));
 sg13g2_o21ai_1 _21652_ (.B1(_03955_),
    .Y(_03956_),
    .A1(net10467),
    .A2(_08180_));
 sg13g2_nand3_1 _21653_ (.B(_08171_),
    .C(_03956_),
    .A(_08563_),
    .Y(_03957_));
 sg13g2_nand2_1 _21654_ (.Y(_03958_),
    .A(_03919_),
    .B(_03957_));
 sg13g2_a21oi_2 _21655_ (.B1(_00095_),
    .Y(_03959_),
    .A2(_03958_),
    .A1(net9729));
 sg13g2_buf_16 clkbuf_leaf_341_clk (.X(clknet_leaf_341_clk),
    .A(clknet_8_117_0_clk));
 sg13g2_nand3_1 _21657_ (.B(net9706),
    .C(net9683),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[0] ),
    .Y(_03961_));
 sg13g2_o21ai_1 _21658_ (.B1(_03961_),
    .Y(_02128_),
    .A1(_03954_),
    .A2(net9683));
 sg13g2_inv_1 _21659_ (.Y(_03962_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[1] ));
 sg13g2_inv_2 _21660_ (.Y(_03963_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[1] ));
 sg13g2_nand3_1 _21661_ (.B(net10456),
    .C(net9729),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[0] ),
    .Y(_03964_));
 sg13g2_o21ai_1 _21662_ (.B1(_03964_),
    .Y(_03965_),
    .A1(_03963_),
    .A2(net9729));
 sg13g2_nand2_1 _21663_ (.Y(_03966_),
    .A(net9683),
    .B(_03965_));
 sg13g2_o21ai_1 _21664_ (.B1(_03966_),
    .Y(_02129_),
    .A1(_03962_),
    .A2(net9683));
 sg13g2_buf_2 place10139 (.A(_09852_),
    .X(net10139));
 sg13g2_nor3_1 _21666_ (.A(net10463),
    .B(_03954_),
    .C(net10456),
    .Y(_03968_));
 sg13g2_a21oi_1 _21667_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[1] ),
    .A2(net10456),
    .Y(_03969_),
    .B1(_03968_));
 sg13g2_nand2_1 _21668_ (.Y(_03970_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[2] ),
    .B(net9705));
 sg13g2_o21ai_1 _21669_ (.B1(_03970_),
    .Y(_03971_),
    .A1(net9706),
    .A2(_03969_));
 sg13g2_mux2_1 _21670_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[2] ),
    .A1(_03971_),
    .S(net9683),
    .X(_02130_));
 sg13g2_buf_2 place10147 (.A(net10145),
    .X(net10147));
 sg13g2_nor3_1 _21672_ (.A(net10463),
    .B(_03962_),
    .C(net10458),
    .Y(_03973_));
 sg13g2_a21oi_1 _21673_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[2] ),
    .A2(net10458),
    .Y(_03974_),
    .B1(_03973_));
 sg13g2_nand2_1 _21674_ (.Y(_03975_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[3] ),
    .B(net9706));
 sg13g2_o21ai_1 _21675_ (.B1(_03975_),
    .Y(_03976_),
    .A1(net9706),
    .A2(_03974_));
 sg13g2_mux2_1 _21676_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[3] ),
    .A1(_03976_),
    .S(net9683),
    .X(_02131_));
 sg13g2_and2_1 _21677_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[3] ),
    .B(net10456),
    .X(_03977_));
 sg13g2_a221oi_1 _21678_ (.B2(net10260),
    .C1(_03977_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[2] ),
    .A1(net10462),
    .Y(_03978_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[0] ));
 sg13g2_nor2_1 _21679_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[4] ),
    .B(_08209_),
    .Y(_03979_));
 sg13g2_a21oi_1 _21680_ (.A1(net9729),
    .A2(_03978_),
    .Y(_03980_),
    .B1(_03979_));
 sg13g2_mux2_1 _21681_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[4] ),
    .A1(_03980_),
    .S(_03959_),
    .X(_02132_));
 sg13g2_and2_1 _21682_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[4] ),
    .B(net10456),
    .X(_03981_));
 sg13g2_a221oi_1 _21683_ (.B2(net10260),
    .C1(_03981_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[3] ),
    .A1(net10462),
    .Y(_03982_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[1] ));
 sg13g2_nor2_1 _21684_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[5] ),
    .B(net9729),
    .Y(_03983_));
 sg13g2_a21oi_1 _21685_ (.A1(net9729),
    .A2(_03982_),
    .Y(_03984_),
    .B1(_03983_));
 sg13g2_mux2_1 _21686_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[5] ),
    .A1(_03984_),
    .S(net9683),
    .X(_02133_));
 sg13g2_and2_1 _21687_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[5] ),
    .B(net10457),
    .X(_03985_));
 sg13g2_a221oi_1 _21688_ (.B2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[4] ),
    .C1(_03985_),
    .B1(net10260),
    .A1(net10462),
    .Y(_03986_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[2] ));
 sg13g2_nor2_1 _21689_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[6] ),
    .B(net9726),
    .Y(_03987_));
 sg13g2_a21oi_1 _21690_ (.A1(net9729),
    .A2(_03986_),
    .Y(_03988_),
    .B1(_03987_));
 sg13g2_mux2_1 _21691_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[6] ),
    .A1(_03988_),
    .S(_03959_),
    .X(_02134_));
 sg13g2_and2_1 _21692_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[6] ),
    .B(net10457),
    .X(_03989_));
 sg13g2_a221oi_1 _21693_ (.B2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[5] ),
    .C1(_03989_),
    .B1(net10260),
    .A1(net10462),
    .Y(_03990_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[3] ));
 sg13g2_nor2_2 _21694_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[7] ),
    .B(net9727),
    .Y(_03991_));
 sg13g2_a21oi_1 _21695_ (.A1(net9729),
    .A2(_03990_),
    .Y(_03992_),
    .B1(_03991_));
 sg13g2_mux2_1 _21696_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[7] ),
    .A1(_03992_),
    .S(_03959_),
    .X(_02135_));
 sg13g2_nand2_1 _21697_ (.Y(_03993_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[30] ),
    .B(net9807));
 sg13g2_o21ai_1 _21698_ (.B1(_03993_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[30] ),
    .A1(net9807),
    .A2(_09178_));
 sg13g2_inv_2 _21699_ (.Y(_03994_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[10] ));
 sg13g2_nand2_1 _21700_ (.Y(_03995_),
    .A(net9703),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[30] ));
 sg13g2_o21ai_1 _21701_ (.B1(_03995_),
    .Y(_01714_),
    .A1(_03994_),
    .A2(net9703));
 sg13g2_mux2_1 _21702_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12] ),
    .A1(_08474_),
    .S(_08490_),
    .X(_01715_));
 sg13g2_inv_2 _21703_ (.Y(_03996_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[13] ));
 sg13g2_nand2_2 _21704_ (.Y(_03997_),
    .A(_08468_),
    .B(_08490_));
 sg13g2_o21ai_1 _21705_ (.B1(_03997_),
    .Y(_01716_),
    .A1(_03996_),
    .A2(net9700));
 sg13g2_inv_2 _21706_ (.Y(_03998_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[14] ));
 sg13g2_nand2_2 _21707_ (.Y(_03999_),
    .A(_08480_),
    .B(_08490_));
 sg13g2_o21ai_1 _21708_ (.B1(_03999_),
    .Y(_01717_),
    .A1(_03998_),
    .A2(net9700));
 sg13g2_nand2_1 _21709_ (.Y(_04000_),
    .A(net9805),
    .B(_09208_));
 sg13g2_o21ai_1 _21710_ (.B1(_04000_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[31] ),
    .A1(_11547_),
    .A2(net9805));
 sg13g2_inv_8 _21711_ (.Y(_04001_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20] ));
 sg13g2_nand2_1 _21712_ (.Y(_04002_),
    .A(net9701),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[31] ));
 sg13g2_o21ai_1 _21713_ (.B1(_04002_),
    .Y(_01718_),
    .A1(_04001_),
    .A2(net9701));
 sg13g2_mux2_1 _21714_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[25] ),
    .A1(_09012_),
    .S(_08417_),
    .X(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[25] ));
 sg13g2_mux2_1 _21715_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[5] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[25] ),
    .S(net9702),
    .X(_01719_));
 sg13g2_nand2_1 _21716_ (.Y(_04003_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[26] ),
    .B(net9809));
 sg13g2_o21ai_1 _21717_ (.B1(_04003_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[26] ),
    .A1(net9809),
    .A2(_09042_));
 sg13g2_mux2_1 _21718_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[6] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[26] ),
    .S(net9702),
    .X(_01720_));
 sg13g2_nand2_1 _21719_ (.Y(_04004_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27] ),
    .B(_07936_));
 sg13g2_o21ai_1 _21720_ (.B1(_04004_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[27] ),
    .A1(_07936_),
    .A2(_09074_));
 sg13g2_inv_2 _21721_ (.Y(_04005_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[7] ));
 sg13g2_nand2_1 _21722_ (.Y(_04006_),
    .A(net9702),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[27] ));
 sg13g2_o21ai_1 _21723_ (.B1(_04006_),
    .Y(_01721_),
    .A1(_04005_),
    .A2(net9703));
 sg13g2_nand2_1 _21724_ (.Y(_04007_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[28] ),
    .B(net9807));
 sg13g2_o21ai_1 _21725_ (.B1(_04007_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[28] ),
    .A1(_07936_),
    .A2(_09106_));
 sg13g2_inv_1 _21726_ (.Y(_04008_),
    .A(net10663));
 sg13g2_nand2_1 _21727_ (.Y(_04009_),
    .A(net9703),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[28] ));
 sg13g2_o21ai_1 _21728_ (.B1(_04009_),
    .Y(_01722_),
    .A1(_04008_),
    .A2(net9703));
 sg13g2_nand2_1 _21729_ (.Y(_04010_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[29] ),
    .B(net9806));
 sg13g2_o21ai_1 _21730_ (.B1(_04010_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[29] ),
    .A1(net9806),
    .A2(_09378_));
 sg13g2_inv_4 _21731_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[9] ),
    .Y(_04011_));
 sg13g2_nand2_1 _21732_ (.Y(_04012_),
    .A(net9703),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[29] ));
 sg13g2_o21ai_1 _21733_ (.B1(_04012_),
    .Y(_01723_),
    .A1(_04011_),
    .A2(net9703));
 sg13g2_mux2_1 _21734_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[7] ),
    .A1(_09217_),
    .S(net9805),
    .X(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[7] ));
 sg13g2_mux2_1 _21735_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[0] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[7] ),
    .S(net9702),
    .X(_01724_));
 sg13g2_mux2_1 _21736_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[8] ),
    .A1(_08979_),
    .S(net9805),
    .X(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[8] ));
 sg13g2_mux2_1 _21737_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[1] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[8] ),
    .S(net9704),
    .X(_01725_));
 sg13g2_mux2_1 _21738_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[9] ),
    .A1(_09016_),
    .S(_08417_),
    .X(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[9] ));
 sg13g2_mux2_1 _21739_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[2] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[9] ),
    .S(net9704),
    .X(_01726_));
 sg13g2_nand2_1 _21740_ (.Y(_04013_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[10] ),
    .B(net9809));
 sg13g2_o21ai_1 _21741_ (.B1(_04013_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[10] ),
    .A1(net9809),
    .A2(_09046_));
 sg13g2_mux2_1 _21742_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[3] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[10] ),
    .S(net9704),
    .X(_01727_));
 sg13g2_nand2_1 _21743_ (.Y(_04014_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[11] ),
    .B(net9809));
 sg13g2_o21ai_1 _21744_ (.B1(_04014_),
    .Y(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[11] ),
    .A1(net9809),
    .A2(_09078_));
 sg13g2_mux2_1 _21745_ (.A0(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[4] ),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[11] ),
    .S(net9704),
    .X(_01728_));
 sg13g2_nand3b_1 _21746_ (.B(_08490_),
    .C(_08449_),
    .Y(_04015_),
    .A_N(_08460_));
 sg13g2_buf_2 place10128 (.A(net10126),
    .X(net10128));
 sg13g2_and3_2 _21748_ (.X(_04017_),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[0] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[1] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[2] ));
 sg13g2_nand2_1 _21749_ (.Y(_04018_),
    .A(_08415_),
    .B(_08428_));
 sg13g2_nor3_1 _21750_ (.A(net9810),
    .B(_08434_),
    .C(_04018_),
    .Y(_04019_));
 sg13g2_a21oi_1 _21751_ (.A1(net9811),
    .A2(_04017_),
    .Y(_04020_),
    .B1(_04019_));
 sg13g2_or2_1 _21752_ (.X(_04021_),
    .B(_04020_),
    .A(_08441_));
 sg13g2_or2_1 _21753_ (.X(_04022_),
    .B(_04021_),
    .A(_04015_));
 sg13g2_nand2_1 _21754_ (.Y(_04023_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_auipc ),
    .B(net9699));
 sg13g2_o21ai_1 _21755_ (.B1(_04023_),
    .Y(_01734_),
    .A1(_08455_),
    .A2(_04022_));
 sg13g2_buf_2 place10126 (.A(_10111_),
    .X(net10126));
 sg13g2_inv_1 _21757_ (.Y(_04025_),
    .A(_04020_));
 sg13g2_nand2_1 _21758_ (.Y(_04026_),
    .A(_08455_),
    .B(_08460_));
 sg13g2_nor3_2 _21759_ (.A(_08449_),
    .B(_08581_),
    .C(_04026_),
    .Y(_04027_));
 sg13g2_nand3_1 _21760_ (.B(_04025_),
    .C(_04027_),
    .A(_08441_),
    .Y(_04028_));
 sg13g2_o21ai_1 _21761_ (.B1(_04028_),
    .Y(_01742_),
    .A1(net10362),
    .A2(net9700));
 sg13g2_nor4_1 _21762_ (.A(_08468_),
    .B(_08474_),
    .C(_08480_),
    .D(_04021_),
    .Y(_04029_));
 sg13g2_a22oi_1 _21763_ (.Y(_04030_),
    .B1(_04027_),
    .B2(_04029_),
    .A2(_08581_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_jalr ));
 sg13g2_inv_1 _21764_ (.Y(_01743_),
    .A(_04030_));
 sg13g2_nor2b_1 _21765_ (.A(_04022_),
    .B_N(_08455_),
    .Y(_04031_));
 sg13g2_a21o_1 _21766_ (.A2(net9699),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_lui ),
    .B1(_04031_),
    .X(_01748_));
 sg13g2_mux2_1 _21767_ (.A0(_11545_),
    .A1(_04018_),
    .S(net9804),
    .X(_04032_));
 sg13g2_nor3_2 _21768_ (.A(_00115_),
    .B(_08441_),
    .C(_04032_),
    .Y(_04033_));
 sg13g2_nand2b_1 _21769_ (.Y(_04034_),
    .B(_04033_),
    .A_N(_08455_));
 sg13g2_nand2_1 _21770_ (.Y(_04035_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_alu_reg_imm ),
    .B(net9699));
 sg13g2_o21ai_1 _21771_ (.B1(_04035_),
    .Y(_01772_),
    .A1(_04015_),
    .A2(_04034_));
 sg13g2_nand2_1 _21772_ (.Y(_04036_),
    .A(_08455_),
    .B(_04033_));
 sg13g2_nand2_1 _21773_ (.Y(_04037_),
    .A(\u_ac_controller_soc_inst.u_picorv32.is_alu_reg_reg ),
    .B(net9699));
 sg13g2_o21ai_1 _21774_ (.B1(_04037_),
    .Y(_01773_),
    .A1(_04015_),
    .A2(_04036_));
 sg13g2_or2_1 _21775_ (.X(_04038_),
    .B(_08460_),
    .A(_08449_));
 sg13g2_nor3_1 _21776_ (.A(net9699),
    .B(_04034_),
    .C(_04038_),
    .Y(_04039_));
 sg13g2_a21o_1 _21777_ (.A2(net9699),
    .A1(\u_ac_controller_soc_inst.u_picorv32.is_lb_lh_lw_lbu_lhu ),
    .B1(_04039_),
    .X(_01777_));
 sg13g2_nor3_1 _21778_ (.A(net9699),
    .B(_04036_),
    .C(_04038_),
    .Y(_04040_));
 sg13g2_a21o_1 _21779_ (.A2(net9699),
    .A1(\u_ac_controller_soc_inst.u_picorv32.is_sb_sh_sw ),
    .B1(_04040_),
    .X(_01778_));
 sg13g2_nor2_1 _21780_ (.A(\u_ac_controller_soc_inst.sram_ready ),
    .B(net11004),
    .Y(_04041_));
 sg13g2_and2_1 _21781_ (.A(_07907_),
    .B(_04041_),
    .X(_00143_));
 sg13g2_inv_1 _21782_ (.Y(_04042_),
    .A(_00139_));
 sg13g2_buf_2 place10143 (.A(net10142),
    .X(net10143));
 sg13g2_buf_2 place10142 (.A(net10141),
    .X(net10142));
 sg13g2_buf_2 place10141 (.A(_09852_),
    .X(net10141));
 sg13g2_nor2b_1 _21786_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[10] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10] ),
    .Y(_04046_));
 sg13g2_buf_2 place10127 (.A(net10126),
    .X(net10127));
 sg13g2_buf_2 place10140 (.A(net10139),
    .X(net10140));
 sg13g2_inv_1 _21789_ (.Y(_04049_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[8] ));
 sg13g2_buf_16 clkbuf_leaf_344_clk (.X(clknet_leaf_344_clk),
    .A(clknet_8_94_0_clk));
 sg13g2_inv_4 _21791_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[7] ),
    .Y(_04051_));
 sg13g2_buf_16 clkbuf_leaf_343_clk (.X(clknet_leaf_343_clk),
    .A(clknet_8_94_0_clk));
 sg13g2_inv_4 _21793_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[5] ),
    .Y(_04053_));
 sg13g2_buf_2 place10118 (.A(_10171_),
    .X(net10118));
 sg13g2_inv_1 _21795_ (.Y(_04055_),
    .A(net10761));
 sg13g2_buf_2 place10119 (.A(net10118),
    .X(net10119));
 sg13g2_inv_1 _21797_ (.Y(_04057_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[4] ));
 sg13g2_inv_1 _21798_ (.Y(_04058_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[3] ));
 sg13g2_inv_1 _21799_ (.Y(_04059_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[2] ));
 sg13g2_buf_2 place10117 (.A(_10171_),
    .X(net10117));
 sg13g2_nor2_1 _21801_ (.A(_04059_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2] ),
    .Y(_04061_));
 sg13g2_buf_2 place10125 (.A(net10122),
    .X(net10125));
 sg13g2_inv_1 _21803_ (.Y(_04063_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[1] ));
 sg13g2_buf_2 place10121 (.A(net10120),
    .X(net10121));
 sg13g2_nor2b_1 _21805_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[0] ),
    .Y(_04065_));
 sg13g2_nand2_1 _21806_ (.Y(_04066_),
    .A(_04063_),
    .B(_04065_));
 sg13g2_o21ai_1 _21807_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[1] ),
    .Y(_04067_),
    .A1(_04063_),
    .A2(_04065_));
 sg13g2_a22oi_1 _21808_ (.Y(_04068_),
    .B1(_04066_),
    .B2(_04067_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2] ),
    .A1(_04059_));
 sg13g2_buf_2 place10124 (.A(net10122),
    .X(net10124));
 sg13g2_inv_2 _21810_ (.Y(_04070_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[3] ));
 sg13g2_o21ai_1 _21811_ (.B1(_04070_),
    .Y(_04071_),
    .A1(_04061_),
    .A2(_04068_));
 sg13g2_nor3_1 _21812_ (.A(_04070_),
    .B(_04061_),
    .C(_04068_),
    .Y(_04072_));
 sg13g2_a221oi_1 _21813_ (.B2(_04071_),
    .C1(_04072_),
    .B1(_04058_),
    .A1(net10761),
    .Y(_04073_),
    .A2(_04057_));
 sg13g2_a221oi_1 _21814_ (.B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[4] ),
    .C1(_04073_),
    .B1(_04055_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[5] ),
    .Y(_04074_),
    .A2(_04053_));
 sg13g2_buf_2 place10120 (.A(net10119),
    .X(net10120));
 sg13g2_buf_2 place10122 (.A(_10171_),
    .X(net10122));
 sg13g2_nand2b_1 _21817_ (.Y(_04077_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[6] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[6] ));
 sg13g2_o21ai_1 _21818_ (.B1(_04077_),
    .Y(_04078_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[5] ),
    .A2(_04053_));
 sg13g2_nand2b_1 _21819_ (.Y(_04079_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[6] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[6] ));
 sg13g2_o21ai_1 _21820_ (.B1(_04079_),
    .Y(_04080_),
    .A1(_04074_),
    .A2(_04078_));
 sg13g2_o21ai_1 _21821_ (.B1(_04080_),
    .Y(_04081_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[7] ),
    .A2(_04051_));
 sg13g2_inv_2 _21822_ (.Y(_04082_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[8] ));
 sg13g2_a22oi_1 _21823_ (.Y(_04083_),
    .B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[7] ),
    .B2(_04051_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[8] ),
    .A1(_04082_));
 sg13g2_a22oi_1 _21824_ (.Y(_04084_),
    .B1(_04081_),
    .B2(_04083_),
    .A2(_04049_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[8] ));
 sg13g2_inv_1 _21825_ (.Y(_04085_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[9] ));
 sg13g2_buf_2 place10123 (.A(net10122),
    .X(net10123));
 sg13g2_nand2_1 _21827_ (.Y(_04087_),
    .A(_04085_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9] ));
 sg13g2_nor2_1 _21828_ (.A(_04085_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9] ),
    .Y(_04088_));
 sg13g2_a21oi_1 _21829_ (.A1(_04084_),
    .A2(_04087_),
    .Y(_04089_),
    .B1(_04088_));
 sg13g2_inv_2 _21830_ (.Y(_04090_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[11] ));
 sg13g2_nor2b_1 _21831_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[10] ),
    .Y(_04091_));
 sg13g2_nor2_1 _21832_ (.A(_04090_),
    .B(_04091_),
    .Y(_04092_));
 sg13g2_buf_2 place10116 (.A(net10115),
    .X(net10116));
 sg13g2_inv_1 _21834_ (.Y(_04094_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[12] ));
 sg13g2_buf_2 place10109 (.A(net10107),
    .X(net10109));
 sg13g2_o21ai_1 _21836_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[11] ),
    .Y(_04096_),
    .A1(_04094_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[12] ));
 sg13g2_a221oi_1 _21837_ (.B2(_04092_),
    .C1(_04096_),
    .B1(_04089_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[11] ),
    .Y(_04097_),
    .A2(_04046_));
 sg13g2_inv_1 _21838_ (.Y(_04098_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[12] ));
 sg13g2_nor3_1 _21839_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[11] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9] ),
    .C(_04046_),
    .Y(_04099_));
 sg13g2_nor3_1 _21840_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[11] ),
    .B(_04085_),
    .C(_04046_),
    .Y(_04100_));
 sg13g2_o21ai_1 _21841_ (.B1(_04084_),
    .Y(_04101_),
    .A1(_04099_),
    .A2(_04100_));
 sg13g2_inv_1 _21842_ (.Y(_04102_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9] ));
 sg13g2_a22oi_1 _21843_ (.Y(_04103_),
    .B1(_04100_),
    .B2(_04102_),
    .A2(_04091_),
    .A1(_04090_));
 sg13g2_a22oi_1 _21844_ (.Y(_04104_),
    .B1(_04101_),
    .B2(_04103_),
    .A2(_04098_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[12] ));
 sg13g2_buf_2 place10164 (.A(net10163),
    .X(net10164));
 sg13g2_buf_2 place10114 (.A(net10113),
    .X(net10114));
 sg13g2_nand2b_1 _21847_ (.Y(_04107_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[29] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[29] ));
 sg13g2_buf_2 place10113 (.A(net10112),
    .X(net10113));
 sg13g2_buf_2 place10112 (.A(net10111),
    .X(net10112));
 sg13g2_xnor2_1 _21850_ (.Y(_04110_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[28] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[28] ));
 sg13g2_inv_1 _21851_ (.Y(_04111_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[31] ));
 sg13g2_buf_2 place10108 (.A(net10107),
    .X(net10108));
 sg13g2_nor2_1 _21853_ (.A(_04111_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[31] ),
    .Y(_04113_));
 sg13g2_nor2b_1 _21854_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[29] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[29] ),
    .Y(_04114_));
 sg13g2_buf_2 place10110 (.A(net10107),
    .X(net10110));
 sg13g2_buf_2 place10107 (.A(_10253_),
    .X(net10107));
 sg13g2_nor2b_1 _21857_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[30] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[30] ),
    .Y(_04117_));
 sg13g2_inv_1 _21858_ (.Y(_04118_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[30] ));
 sg13g2_nand2_1 _21859_ (.Y(_04119_),
    .A(_04111_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[31] ));
 sg13g2_o21ai_1 _21860_ (.B1(_04119_),
    .Y(_04120_),
    .A1(_04118_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[30] ));
 sg13g2_nor4_1 _21861_ (.A(_04113_),
    .B(_04114_),
    .C(_04117_),
    .D(_04120_),
    .Y(_04121_));
 sg13g2_buf_2 place10115 (.A(net10111),
    .X(net10115));
 sg13g2_buf_16 clkbuf_leaf_346_clk (.X(clknet_leaf_346_clk),
    .A(clknet_8_117_0_clk));
 sg13g2_xor2_1 _21864_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[24] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24] ),
    .X(_04124_));
 sg13g2_buf_2 place10104 (.A(net10103),
    .X(net10104));
 sg13g2_buf_2 place10106 (.A(net10105),
    .X(net10106));
 sg13g2_xor2_1 _21867_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[26] ),
    .X(_04127_));
 sg13g2_buf_2 place10105 (.A(_10335_),
    .X(net10105));
 sg13g2_buf_2 place10103 (.A(_10335_),
    .X(net10103));
 sg13g2_xor2_1 _21870_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[25] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[25] ),
    .X(_04130_));
 sg13g2_buf_2 place10099 (.A(net10097),
    .X(net10099));
 sg13g2_buf_2 place10098 (.A(net10097),
    .X(net10098));
 sg13g2_xor2_1 _21873_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[27] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[27] ),
    .X(_04133_));
 sg13g2_nor4_1 _21874_ (.A(_04124_),
    .B(_04127_),
    .C(_04130_),
    .D(_04133_),
    .Y(_04134_));
 sg13g2_and4_2 _21875_ (.A(_04107_),
    .B(_04110_),
    .C(_04121_),
    .D(_04134_),
    .X(_04135_));
 sg13g2_buf_2 place10101 (.A(net10100),
    .X(net10101));
 sg13g2_buf_2 place10100 (.A(net10097),
    .X(net10100));
 sg13g2_xor2_1 _21878_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[23] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[23] ),
    .X(_04138_));
 sg13g2_buf_2 place10102 (.A(net10101),
    .X(net10102));
 sg13g2_buf_16 clkbuf_leaf_348_clk (.X(clknet_leaf_348_clk),
    .A(clknet_8_119_0_clk));
 sg13g2_nor2b_1 _21881_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[22] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22] ),
    .Y(_04141_));
 sg13g2_nor2b_1 _21882_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[22] ),
    .Y(_04142_));
 sg13g2_buf_2 place10203 (.A(net10202),
    .X(net10203));
 sg13g2_buf_2 place10093 (.A(net10092),
    .X(net10093));
 sg13g2_nor2b_1 _21885_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[21] ),
    .Y(_04145_));
 sg13g2_nor4_1 _21886_ (.A(_04138_),
    .B(_04141_),
    .C(_04142_),
    .D(_04145_),
    .Y(_04146_));
 sg13g2_nor2b_1 _21887_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[21] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21] ),
    .Y(_04147_));
 sg13g2_buf_2 place10096 (.A(net10092),
    .X(net10096));
 sg13g2_buf_2 place10095 (.A(net10092),
    .X(net10095));
 sg13g2_xor2_1 _21890_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[20] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[20] ),
    .X(_04150_));
 sg13g2_buf_2 place10088 (.A(_10415_),
    .X(net10088));
 sg13g2_inv_2 _21892_ (.Y(_04152_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[16] ));
 sg13g2_buf_2 place10092 (.A(_10415_),
    .X(net10092));
 sg13g2_buf_2 place10091 (.A(net10090),
    .X(net10091));
 sg13g2_nand2b_1 _21895_ (.Y(_04155_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[17] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[17] ));
 sg13g2_o21ai_1 _21896_ (.B1(_04155_),
    .Y(_04156_),
    .A1(_04152_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[16] ));
 sg13g2_nor2b_1 _21897_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[16] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[16] ),
    .Y(_04157_));
 sg13g2_nor4_1 _21898_ (.A(_04147_),
    .B(_04150_),
    .C(_04156_),
    .D(_04157_),
    .Y(_04158_));
 sg13g2_inv_2 _21899_ (.Y(_04159_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[17] ));
 sg13g2_buf_2 place10204 (.A(net10203),
    .X(net10204));
 sg13g2_buf_2 place10094 (.A(net10092),
    .X(net10094));
 sg13g2_nand2_1 _21902_ (.Y(_04162_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[18] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[18] ));
 sg13g2_or2_1 _21903_ (.X(_04163_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[18] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[18] ));
 sg13g2_buf_2 place10082 (.A(net10081),
    .X(net10082));
 sg13g2_buf_2 place10158 (.A(net10156),
    .X(net10158));
 sg13g2_xor2_1 _21906_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[19] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[19] ),
    .X(_04166_));
 sg13g2_a221oi_1 _21907_ (.B2(_04163_),
    .C1(_04166_),
    .B1(_04162_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[17] ),
    .Y(_04167_),
    .A2(_04159_));
 sg13g2_and4_2 _21908_ (.A(_04135_),
    .B(_04146_),
    .C(_04158_),
    .D(_04167_),
    .X(_04168_));
 sg13g2_buf_2 place10244 (.A(_07931_),
    .X(net10244));
 sg13g2_buf_2 place10080 (.A(net10079),
    .X(net10080));
 sg13g2_xnor2_1 _21911_ (.Y(_04171_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[15] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[15] ));
 sg13g2_buf_2 place10087 (.A(net10086),
    .X(net10087));
 sg13g2_buf_2 place10081 (.A(net10079),
    .X(net10081));
 sg13g2_xnor2_1 _21914_ (.Y(_04174_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[14] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14] ));
 sg13g2_buf_2 place10086 (.A(_10568_),
    .X(net10086));
 sg13g2_buf_2 place10079 (.A(_10568_),
    .X(net10079));
 sg13g2_nand2b_1 _21917_ (.Y(_04177_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[13] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[13] ));
 sg13g2_nand3_1 _21918_ (.B(_04174_),
    .C(_04177_),
    .A(_04171_),
    .Y(_04178_));
 sg13g2_inv_1 _21919_ (.Y(_04179_),
    .A(_04178_));
 sg13g2_nand2_1 _21920_ (.Y(_04180_),
    .A(_04094_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[12] ));
 sg13g2_nand3_1 _21921_ (.B(_04179_),
    .C(_04180_),
    .A(_04168_),
    .Y(_04181_));
 sg13g2_nor3_2 _21922_ (.A(_04097_),
    .B(_04104_),
    .C(_04181_),
    .Y(_04182_));
 sg13g2_inv_1 _21923_ (.Y(_04183_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[28] ));
 sg13g2_inv_2 _21924_ (.Y(_04184_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[27] ));
 sg13g2_inv_1 _21925_ (.Y(_04185_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[27] ));
 sg13g2_inv_1 _21926_ (.Y(_04186_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26] ));
 sg13g2_nand2_1 _21927_ (.Y(_04187_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[26] ),
    .B(_04186_));
 sg13g2_nor2b_1 _21928_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[24] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24] ),
    .Y(_04188_));
 sg13g2_nand2_1 _21929_ (.Y(_04189_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[25] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24] ));
 sg13g2_o21ai_1 _21930_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[25] ),
    .Y(_04190_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[24] ),
    .A2(_04189_));
 sg13g2_o21ai_1 _21931_ (.B1(_04190_),
    .Y(_04191_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[25] ),
    .A2(_04188_));
 sg13g2_o21ai_1 _21932_ (.B1(_04191_),
    .Y(_04192_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[26] ),
    .A2(_04186_));
 sg13g2_a22oi_1 _21933_ (.Y(_04193_),
    .B1(_04187_),
    .B2(_04192_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[27] ),
    .A1(_04185_));
 sg13g2_a221oi_1 _21934_ (.B2(_04184_),
    .C1(_04193_),
    .B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[27] ),
    .A1(_04183_),
    .Y(_04194_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[28] ));
 sg13g2_o21ai_1 _21935_ (.B1(_04107_),
    .Y(_04195_),
    .A1(_04183_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[28] ));
 sg13g2_o21ai_1 _21936_ (.B1(_04121_),
    .Y(_04196_),
    .A1(_04194_),
    .A2(_04195_));
 sg13g2_inv_2 _21937_ (.Y(_04197_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[20] ));
 sg13g2_inv_2 _21938_ (.Y(_04198_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[18] ));
 sg13g2_inv_1 _21939_ (.Y(_04199_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[19] ));
 sg13g2_o21ai_1 _21940_ (.B1(_04199_),
    .Y(_04200_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[18] ),
    .A2(_04198_));
 sg13g2_nand2_2 _21941_ (.Y(_04201_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[19] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[18] ));
 sg13g2_o21ai_1 _21942_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[19] ),
    .Y(_04202_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[18] ),
    .A2(_04201_));
 sg13g2_a22oi_1 _21943_ (.Y(_04203_),
    .B1(_04200_),
    .B2(_04202_),
    .A2(_04167_),
    .A1(_04156_));
 sg13g2_o21ai_1 _21944_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[20] ),
    .Y(_04204_),
    .A1(_04197_),
    .A2(_04203_));
 sg13g2_nand2_1 _21945_ (.Y(_04205_),
    .A(_04197_),
    .B(_04203_));
 sg13g2_a21oi_1 _21946_ (.A1(_04204_),
    .A2(_04205_),
    .Y(_04206_),
    .B1(_04147_));
 sg13g2_nand2b_1 _21947_ (.Y(_04207_),
    .B(_04146_),
    .A_N(_04206_));
 sg13g2_nand2_1 _21948_ (.Y(_04208_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[23] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22] ));
 sg13g2_o21ai_1 _21949_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[23] ),
    .Y(_04209_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[22] ),
    .A2(_04208_));
 sg13g2_o21ai_1 _21950_ (.B1(_04209_),
    .Y(_04210_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[23] ),
    .A2(_04141_));
 sg13g2_nand2_1 _21951_ (.Y(_04211_),
    .A(_04207_),
    .B(_04210_));
 sg13g2_nand2b_1 _21952_ (.Y(_04212_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[13] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[13] ));
 sg13g2_nor2b_1 _21953_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[14] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14] ),
    .Y(_04213_));
 sg13g2_nand2_1 _21954_ (.Y(_04214_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[15] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14] ));
 sg13g2_o21ai_1 _21955_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[15] ),
    .Y(_04215_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[14] ),
    .A2(_04214_));
 sg13g2_o21ai_1 _21956_ (.B1(_04215_),
    .Y(_04216_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[15] ),
    .A2(_04213_));
 sg13g2_o21ai_1 _21957_ (.B1(_04216_),
    .Y(_04217_),
    .A1(_04178_),
    .A2(_04212_));
 sg13g2_nand2_2 _21958_ (.Y(_04218_),
    .A(net11038),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_enable ));
 sg13g2_o21ai_1 _21959_ (.B1(_04119_),
    .Y(_04219_),
    .A1(_04113_),
    .A2(_04117_));
 sg13g2_nand2b_1 _21960_ (.Y(_04220_),
    .B(_04219_),
    .A_N(_04218_));
 sg13g2_a221oi_1 _21961_ (.B2(_04168_),
    .C1(_04220_),
    .B1(_04217_),
    .A1(_04135_),
    .Y(_04221_),
    .A2(_04211_));
 sg13g2_nand3b_1 _21962_ (.B(_04196_),
    .C(_04221_),
    .Y(_04222_),
    .A_N(_04182_));
 sg13g2_buf_2 place10085 (.A(net10084),
    .X(net10085));
 sg13g2_buf_2 place10083 (.A(net10081),
    .X(net10083));
 sg13g2_nor2_1 _21965_ (.A(_04042_),
    .B(net9628),
    .Y(_00144_));
 sg13g2_and4_2 _21966_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[3] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[1] ),
    .D(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0] ),
    .X(_04225_));
 sg13g2_buf_2 place10071 (.A(net10070),
    .X(net10071));
 sg13g2_nand4_1 _21968_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[5] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[4] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[6] ),
    .Y(_04227_),
    .D(_04225_));
 sg13g2_buf_2 place10077 (.A(net10074),
    .X(net10077));
 sg13g2_nor3_2 _21970_ (.A(_04082_),
    .B(_04051_),
    .C(_04227_),
    .Y(_04229_));
 sg13g2_and2_1 _21971_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9] ),
    .B(_04229_),
    .X(_04230_));
 sg13g2_xnor2_1 _21972_ (.Y(_04231_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10] ),
    .B(_04230_));
 sg13g2_nor2_1 _21973_ (.A(net9627),
    .B(_04231_),
    .Y(_00145_));
 sg13g2_nand2_1 _21974_ (.Y(_04232_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10] ),
    .B(_04230_));
 sg13g2_xnor2_1 _21975_ (.Y(_04233_),
    .A(_04090_),
    .B(_04232_));
 sg13g2_nor2_1 _21976_ (.A(net9627),
    .B(_04233_),
    .Y(_00146_));
 sg13g2_and4_2 _21977_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[11] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9] ),
    .D(_04229_),
    .X(_04234_));
 sg13g2_buf_2 place10166 (.A(_10103_),
    .X(net10166));
 sg13g2_xnor2_1 _21979_ (.Y(_04236_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[12] ),
    .B(_04234_));
 sg13g2_nor2_1 _21980_ (.A(net9627),
    .B(_04236_),
    .Y(_00147_));
 sg13g2_nand2_1 _21981_ (.Y(_04237_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[12] ),
    .B(_04234_));
 sg13g2_xor2_1 _21982_ (.B(_04237_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[13] ),
    .X(_04238_));
 sg13g2_nor2_1 _21983_ (.A(net9627),
    .B(_04238_),
    .Y(_00148_));
 sg13g2_and3_2 _21984_ (.X(_04239_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[13] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[12] ),
    .C(_04234_));
 sg13g2_buf_2 place10076 (.A(net10075),
    .X(net10076));
 sg13g2_xnor2_1 _21986_ (.Y(_04241_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14] ),
    .B(_04239_));
 sg13g2_nor2_1 _21987_ (.A(net9627),
    .B(_04241_),
    .Y(_00149_));
 sg13g2_inv_2 _21988_ (.Y(_04242_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[15] ));
 sg13g2_nand2_1 _21989_ (.Y(_04243_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14] ),
    .B(_04239_));
 sg13g2_xnor2_1 _21990_ (.Y(_04244_),
    .A(_04242_),
    .B(_04243_));
 sg13g2_nor2_1 _21991_ (.A(_04222_),
    .B(_04244_),
    .Y(_00150_));
 sg13g2_nand2b_1 _21992_ (.Y(_04245_),
    .B(_04239_),
    .A_N(_04214_));
 sg13g2_xnor2_1 _21993_ (.Y(_04246_),
    .A(_04152_),
    .B(_04245_));
 sg13g2_nor2_1 _21994_ (.A(_04222_),
    .B(_04246_),
    .Y(_00151_));
 sg13g2_nand4_1 _21995_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[15] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[16] ),
    .Y(_04247_),
    .D(_04239_));
 sg13g2_xnor2_1 _21996_ (.Y(_04248_),
    .A(_04159_),
    .B(_04247_));
 sg13g2_nor2_1 _21997_ (.A(net9630),
    .B(_04248_),
    .Y(_00152_));
 sg13g2_or2_1 _21998_ (.X(_04249_),
    .B(_04247_),
    .A(_04159_));
 sg13g2_buf_2 place10070 (.A(_10648_),
    .X(net10070));
 sg13g2_xnor2_1 _22000_ (.Y(_04251_),
    .A(_04198_),
    .B(_04249_));
 sg13g2_nor2_1 _22001_ (.A(net9630),
    .B(_04251_),
    .Y(_00153_));
 sg13g2_buf_2 place10073 (.A(net10072),
    .X(net10073));
 sg13g2_nor2_1 _22003_ (.A(_04198_),
    .B(_04249_),
    .Y(_04253_));
 sg13g2_xnor2_1 _22004_ (.Y(_04254_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[19] ),
    .B(_04253_));
 sg13g2_nor2_1 _22005_ (.A(net9630),
    .B(_04254_),
    .Y(_00154_));
 sg13g2_xnor2_1 _22006_ (.Y(_04255_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[1] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0] ));
 sg13g2_nor2_1 _22007_ (.A(net9628),
    .B(_04255_),
    .Y(_00155_));
 sg13g2_nor2_1 _22008_ (.A(_04201_),
    .B(_04249_),
    .Y(_04256_));
 sg13g2_xnor2_1 _22009_ (.Y(_04257_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[20] ),
    .B(_04256_));
 sg13g2_nor2_1 _22010_ (.A(net9630),
    .B(_04257_),
    .Y(_00156_));
 sg13g2_nor3_2 _22011_ (.A(_04197_),
    .B(_04201_),
    .C(_04249_),
    .Y(_04258_));
 sg13g2_xnor2_1 _22012_ (.Y(_04259_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21] ),
    .B(_04258_));
 sg13g2_nor2_1 _22013_ (.A(net9630),
    .B(_04259_),
    .Y(_00157_));
 sg13g2_nand2_1 _22014_ (.Y(_04260_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21] ),
    .B(_04258_));
 sg13g2_xor2_1 _22015_ (.B(_04260_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22] ),
    .X(_04261_));
 sg13g2_nor2_1 _22016_ (.A(net9630),
    .B(_04261_),
    .Y(_00158_));
 sg13g2_inv_2 _22017_ (.Y(_04262_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[23] ));
 sg13g2_nand3_1 _22018_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21] ),
    .C(_04258_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22] ),
    .Y(_04263_));
 sg13g2_buf_2 place10072 (.A(net10070),
    .X(net10072));
 sg13g2_xnor2_1 _22020_ (.Y(_04265_),
    .A(_04262_),
    .B(_04263_));
 sg13g2_nor2_1 _22021_ (.A(net9629),
    .B(_04265_),
    .Y(_00159_));
 sg13g2_nor2_1 _22022_ (.A(_04262_),
    .B(_04263_),
    .Y(_04266_));
 sg13g2_xnor2_1 _22023_ (.Y(_04267_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24] ),
    .B(_04266_));
 sg13g2_nor2_1 _22024_ (.A(net9629),
    .B(_04267_),
    .Y(_00160_));
 sg13g2_nand2_1 _22025_ (.Y(_04268_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24] ),
    .B(_04266_));
 sg13g2_xor2_1 _22026_ (.B(_04268_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[25] ),
    .X(_04269_));
 sg13g2_nor2_1 _22027_ (.A(net9629),
    .B(_04269_),
    .Y(_00161_));
 sg13g2_nor3_2 _22028_ (.A(_04262_),
    .B(_04189_),
    .C(_04263_),
    .Y(_04270_));
 sg13g2_xnor2_1 _22029_ (.Y(_04271_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26] ),
    .B(_04270_));
 sg13g2_nor2_1 _22030_ (.A(net9629),
    .B(_04271_),
    .Y(_00162_));
 sg13g2_nand2_1 _22031_ (.Y(_04272_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26] ),
    .B(_04270_));
 sg13g2_xnor2_1 _22032_ (.Y(_04273_),
    .A(_04184_),
    .B(_04272_));
 sg13g2_nor2_1 _22033_ (.A(net9631),
    .B(_04273_),
    .Y(_00163_));
 sg13g2_buf_2 place10074 (.A(_10648_),
    .X(net10074));
 sg13g2_nor2_1 _22035_ (.A(_04184_),
    .B(_04272_),
    .Y(_04275_));
 sg13g2_xnor2_1 _22036_ (.Y(_04276_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[28] ),
    .B(_04275_));
 sg13g2_nor2_1 _22037_ (.A(net9631),
    .B(_04276_),
    .Y(_00164_));
 sg13g2_and4_2 _22038_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[28] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[27] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26] ),
    .D(_04270_),
    .X(_04277_));
 sg13g2_xnor2_1 _22039_ (.Y(_04278_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[29] ),
    .B(_04277_));
 sg13g2_nor2_1 _22040_ (.A(net9631),
    .B(_04278_),
    .Y(_00165_));
 sg13g2_nand2_1 _22041_ (.Y(_04279_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[1] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0] ));
 sg13g2_xor2_1 _22042_ (.B(_04279_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2] ),
    .X(_04280_));
 sg13g2_nor2_1 _22043_ (.A(net9628),
    .B(_04280_),
    .Y(_00166_));
 sg13g2_and2_1 _22044_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[29] ),
    .B(_04277_),
    .X(_04281_));
 sg13g2_xnor2_1 _22045_ (.Y(_04282_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[30] ),
    .B(_04281_));
 sg13g2_nor2_1 _22046_ (.A(net9631),
    .B(_04282_),
    .Y(_00167_));
 sg13g2_a21oi_1 _22047_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[30] ),
    .A2(_04281_),
    .Y(_04283_),
    .B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[31] ));
 sg13g2_nor2_1 _22048_ (.A(net9631),
    .B(_04283_),
    .Y(_00168_));
 sg13g2_nand3_1 _22049_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[1] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2] ),
    .Y(_04284_));
 sg13g2_xnor2_1 _22050_ (.Y(_04285_),
    .A(_04070_),
    .B(_04284_));
 sg13g2_nor2_1 _22051_ (.A(net9628),
    .B(_04285_),
    .Y(_00169_));
 sg13g2_xnor2_1 _22052_ (.Y(_04286_),
    .A(net10761),
    .B(_04225_));
 sg13g2_nor2_1 _22053_ (.A(net9628),
    .B(_04286_),
    .Y(_00170_));
 sg13g2_nand2_1 _22054_ (.Y(_04287_),
    .A(net10761),
    .B(_04225_));
 sg13g2_xnor2_1 _22055_ (.Y(_04288_),
    .A(_04053_),
    .B(_04287_));
 sg13g2_nor2_1 _22056_ (.A(net9628),
    .B(_04288_),
    .Y(_00171_));
 sg13g2_nand3_1 _22057_ (.B(net10761),
    .C(_04225_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[5] ),
    .Y(_04289_));
 sg13g2_xor2_1 _22058_ (.B(_04289_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[6] ),
    .X(_04290_));
 sg13g2_nor2_1 _22059_ (.A(net9628),
    .B(_04290_),
    .Y(_00172_));
 sg13g2_xnor2_1 _22060_ (.Y(_04291_),
    .A(_04051_),
    .B(_04227_));
 sg13g2_nor2_1 _22061_ (.A(net9628),
    .B(_04291_),
    .Y(_00173_));
 sg13g2_nor2_1 _22062_ (.A(_04051_),
    .B(_04227_),
    .Y(_04292_));
 sg13g2_xnor2_1 _22063_ (.Y(_04293_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[8] ),
    .B(_04292_));
 sg13g2_nor2_1 _22064_ (.A(net9627),
    .B(_04293_),
    .Y(_00174_));
 sg13g2_xnor2_1 _22065_ (.Y(_04294_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9] ),
    .B(_04229_));
 sg13g2_nor2_1 _22066_ (.A(net9627),
    .B(_04294_),
    .Y(_00175_));
 sg13g2_nand2_2 _22067_ (.Y(_04295_),
    .A(\u_ac_controller_soc_inst.cbus_valid ),
    .B(_07886_));
 sg13g2_buf_2 place10075 (.A(net10074),
    .X(net10075));
 sg13g2_buf_2 place10069 (.A(_10648_),
    .X(net10069));
 sg13g2_buf_2 place10063 (.A(net10061),
    .X(net10063));
 sg13g2_buf_2 place10065 (.A(net10064),
    .X(net10065));
 sg13g2_buf_2 place10061 (.A(_10730_),
    .X(net10061));
 sg13g2_buf_2 place10962 (.A(net10960),
    .X(net10962));
 sg13g2_inv_1 _22074_ (.Y(_04302_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[34] ));
 sg13g2_buf_2 place10068 (.A(net10064),
    .X(net10068));
 sg13g2_nand3_1 _22076_ (.B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[33] ),
    .C(net10236),
    .A(net10749),
    .Y(_04304_));
 sg13g2_o21ai_1 _22077_ (.B1(_04304_),
    .Y(_04305_),
    .A1(net10749),
    .A2(_04302_));
 sg13g2_buf_2 place10798 (.A(net10797),
    .X(net10798));
 sg13g2_buf_2 place10062 (.A(net10061),
    .X(net10062));
 sg13g2_buf_2 place10064 (.A(_10730_),
    .X(net10064));
 sg13g2_a22oi_1 _22081_ (.Y(_04309_),
    .B1(_04305_),
    .B2(net10736),
    .A2(net10149),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[34] ));
 sg13g2_nor2_1 _22082_ (.A(net10979),
    .B(_04309_),
    .Y(_00380_));
 sg13g2_inv_1 _22083_ (.Y(_04310_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[35] ));
 sg13g2_nand3_1 _22084_ (.B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[34] ),
    .C(net10236),
    .A(net10749),
    .Y(_04311_));
 sg13g2_o21ai_1 _22085_ (.B1(_04311_),
    .Y(_04312_),
    .A1(net10749),
    .A2(_04310_));
 sg13g2_a22oi_1 _22086_ (.Y(_04313_),
    .B1(_04312_),
    .B2(net10736),
    .A2(net10149),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[35] ));
 sg13g2_nor2_1 _22087_ (.A(net10979),
    .B(_04313_),
    .Y(_00381_));
 sg13g2_nor2_1 _22088_ (.A(\u_ac_controller_soc_inst.cbus_addr[27] ),
    .B(\u_ac_controller_soc_inst.cbus_addr[26] ),
    .Y(_04314_));
 sg13g2_and4_1 _22089_ (.A(_00104_),
    .B(_04314_),
    .C(_07926_),
    .D(_07895_),
    .X(_04315_));
 sg13g2_o21ai_1 _22090_ (.B1(_07718_),
    .Y(_04316_),
    .A1(_00105_),
    .A2(_04315_));
 sg13g2_nand2b_1 _22091_ (.Y(_04317_),
    .B(_07887_),
    .A_N(\u_ac_controller_soc_inst.spi_sensor_ready ));
 sg13g2_o21ai_1 _22092_ (.B1(spi_sensor_cs_n),
    .Y(_04318_),
    .A1(_04316_),
    .A2(_04317_));
 sg13g2_inv_2 _22093_ (.Y(_04319_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[2] ));
 sg13g2_buf_2 place10067 (.A(net10065),
    .X(net10067));
 sg13g2_nor2b_1 _22095_ (.A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[3] ),
    .Y(_04321_));
 sg13g2_buf_2 place10060 (.A(_10730_),
    .X(net10060));
 sg13g2_xor2_1 _22097_ (.B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[5] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[5] ),
    .X(_04323_));
 sg13g2_buf_2 place10066 (.A(net10065),
    .X(net10066));
 sg13g2_nor2b_1 _22099_ (.A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[4] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[4] ),
    .Y(_04325_));
 sg13g2_nor2b_1 _22100_ (.A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[4] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[4] ),
    .Y(_04326_));
 sg13g2_nor4_1 _22101_ (.A(_04321_),
    .B(_04323_),
    .C(_04325_),
    .D(_04326_),
    .Y(_04327_));
 sg13g2_buf_16 clkbuf_leaf_349_clk (.X(clknet_leaf_349_clk),
    .A(clknet_8_118_0_clk));
 sg13g2_nor2b_1 _22103_ (.A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[3] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3] ),
    .Y(_04329_));
 sg13g2_nor3_1 _22104_ (.A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[1] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[0] ),
    .C(_04329_),
    .Y(_04330_));
 sg13g2_nand3_1 _22105_ (.B(_04327_),
    .C(_04330_),
    .A(_04319_),
    .Y(_04331_));
 sg13g2_nand3_1 _22106_ (.B(_04318_),
    .C(_04331_),
    .A(net11037),
    .Y(_00394_));
 sg13g2_buf_2 place10053 (.A(net10052),
    .X(net10053));
 sg13g2_buf_2 place10089 (.A(net10088),
    .X(net10089));
 sg13g2_xor2_1 _22109_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[27] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[27] ),
    .X(_04334_));
 sg13g2_buf_2 place10052 (.A(_10810_),
    .X(net10052));
 sg13g2_buf_2 place10059 (.A(net10055),
    .X(net10059));
 sg13g2_xor2_1 _22112_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[26] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[26] ),
    .X(_04337_));
 sg13g2_buf_2 place10058 (.A(net10056),
    .X(net10058));
 sg13g2_buf_2 place10056 (.A(net10055),
    .X(net10056));
 sg13g2_nor2b_1 _22115_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[25] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[25] ),
    .Y(_04340_));
 sg13g2_nor3_1 _22116_ (.A(_04334_),
    .B(_04337_),
    .C(_04340_),
    .Y(_04341_));
 sg13g2_buf_2 place10051 (.A(_10810_),
    .X(net10051));
 sg13g2_buf_2 place10055 (.A(_10810_),
    .X(net10055));
 sg13g2_nand2b_2 _22119_ (.Y(_04344_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[30] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[30] ));
 sg13g2_inv_2 _22120_ (.Y(_04345_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[30] ));
 sg13g2_nand2_1 _22121_ (.Y(_04346_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[30] ),
    .B(_04345_));
 sg13g2_buf_2 place10054 (.A(net10052),
    .X(net10054));
 sg13g2_buf_2 place10057 (.A(net10056),
    .X(net10057));
 sg13g2_inv_2 _22124_ (.Y(_04349_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[29] ));
 sg13g2_buf_2 place10048 (.A(net10045),
    .X(net10048));
 sg13g2_xor2_1 _22126_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[31] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[31] ),
    .X(_04351_));
 sg13g2_a21oi_1 _22127_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[29] ),
    .A2(_04349_),
    .Y(_04352_),
    .B1(_04351_));
 sg13g2_nand3_1 _22128_ (.B(_04346_),
    .C(_04352_),
    .A(_04344_),
    .Y(_04353_));
 sg13g2_buf_2 place10050 (.A(net10049),
    .X(net10050));
 sg13g2_buf_2 place10880 (.A(net10878),
    .X(net10880));
 sg13g2_xor2_1 _22131_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[28] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[28] ),
    .X(_04356_));
 sg13g2_buf_2 place10045 (.A(_10891_),
    .X(net10045));
 sg13g2_inv_1 _22133_ (.Y(_04358_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[24] ));
 sg13g2_nor2b_1 _22134_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[25] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[25] ),
    .Y(_04359_));
 sg13g2_a21o_1 _22135_ (.A2(_04358_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[24] ),
    .B1(_04359_),
    .X(_04360_));
 sg13g2_nand2b_1 _22136_ (.Y(_04361_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[29] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[29] ));
 sg13g2_o21ai_1 _22137_ (.B1(_04361_),
    .Y(_04362_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[24] ),
    .A2(_04358_));
 sg13g2_nor4_1 _22138_ (.A(_04353_),
    .B(_04356_),
    .C(_04360_),
    .D(_04362_),
    .Y(_04363_));
 sg13g2_and2_1 _22139_ (.A(_04341_),
    .B(_04363_),
    .X(_04364_));
 sg13g2_buf_2 place10049 (.A(_10891_),
    .X(net10049));
 sg13g2_buf_2 place10043 (.A(net10042),
    .X(net10043));
 sg13g2_nor2b_1 _22142_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[22] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22] ),
    .Y(_04367_));
 sg13g2_nand2b_1 _22143_ (.Y(_04368_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[22] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22] ));
 sg13g2_buf_2 place10042 (.A(_10891_),
    .X(net10042));
 sg13g2_inv_4 _22145_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[21] ),
    .Y(_04370_));
 sg13g2_buf_2 place10044 (.A(net10042),
    .X(net10044));
 sg13g2_buf_2 place10046 (.A(net10045),
    .X(net10046));
 sg13g2_xor2_1 _22148_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[23] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[23] ),
    .X(_04373_));
 sg13g2_a21oi_1 _22149_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[21] ),
    .A2(_04370_),
    .Y(_04374_),
    .B1(_04373_));
 sg13g2_nand3b_1 _22150_ (.B(_04368_),
    .C(_04374_),
    .Y(_04375_),
    .A_N(_04367_));
 sg13g2_inv_1 _22151_ (.Y(_04376_),
    .A(_04375_));
 sg13g2_buf_2 place10047 (.A(net10046),
    .X(net10047));
 sg13g2_buf_2 place10037 (.A(net10036),
    .X(net10037));
 sg13g2_xor2_1 _22154_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[19] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[19] ),
    .X(_04379_));
 sg13g2_buf_2 place10041 (.A(net10040),
    .X(net10041));
 sg13g2_buf_2 place10035 (.A(net10034),
    .X(net10035));
 sg13g2_xor2_1 _22157_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[18] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[18] ),
    .X(_04382_));
 sg13g2_buf_2 place10034 (.A(net10032),
    .X(net10034));
 sg13g2_buf_2 place10090 (.A(net10088),
    .X(net10090));
 sg13g2_nor2b_1 _22160_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[17] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[17] ),
    .Y(_04385_));
 sg13g2_nor3_2 _22161_ (.A(_04379_),
    .B(_04382_),
    .C(_04385_),
    .Y(_04386_));
 sg13g2_nor2_1 _22162_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[21] ),
    .B(_04370_),
    .Y(_04387_));
 sg13g2_buf_2 place10036 (.A(net10032),
    .X(net10036));
 sg13g2_buf_2 place10028 (.A(net10027),
    .X(net10028));
 sg13g2_xor2_1 _22165_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[20] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[20] ),
    .X(_04390_));
 sg13g2_buf_2 place10040 (.A(net10038),
    .X(net10040));
 sg13g2_buf_2 place10039 (.A(net10038),
    .X(net10039));
 sg13g2_nor2b_1 _22168_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[16] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[16] ),
    .Y(_04393_));
 sg13g2_inv_1 _22169_ (.Y(_04394_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[16] ));
 sg13g2_nand2b_1 _22170_ (.Y(_04395_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[17] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[17] ));
 sg13g2_o21ai_1 _22171_ (.B1(_04395_),
    .Y(_04396_),
    .A1(_04394_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[16] ));
 sg13g2_nor4_1 _22172_ (.A(_04387_),
    .B(_04390_),
    .C(_04393_),
    .D(_04396_),
    .Y(_04397_));
 sg13g2_nand4_1 _22173_ (.B(_04376_),
    .C(_04386_),
    .A(_04364_),
    .Y(_04398_),
    .D(_04397_));
 sg13g2_buf_2 place10078 (.A(net10077),
    .X(net10078));
 sg13g2_buf_2 place10031 (.A(net10030),
    .X(net10031));
 sg13g2_xor2_1 _22176_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[11] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[11] ),
    .X(_04401_));
 sg13g2_buf_2 place10016 (.A(_11164_),
    .X(net10016));
 sg13g2_buf_2 place10021 (.A(net10020),
    .X(net10021));
 sg13g2_xor2_1 _22179_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[10] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[10] ),
    .X(_04404_));
 sg13g2_buf_16 clkbuf_leaf_352_clk (.X(clknet_leaf_352_clk),
    .A(clknet_8_118_0_clk));
 sg13g2_buf_16 clkbuf_leaf_350_clk (.X(clknet_leaf_350_clk),
    .A(clknet_8_118_0_clk));
 sg13g2_nor2b_1 _22182_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[9] ),
    .Y(_04407_));
 sg13g2_nor3_1 _22183_ (.A(_04401_),
    .B(_04404_),
    .C(_04407_),
    .Y(_04408_));
 sg13g2_buf_2 place10024 (.A(net10023),
    .X(net10024));
 sg13g2_buf_2 place10004 (.A(_11244_),
    .X(net10004));
 sg13g2_xnor2_1 _22186_ (.Y(_04411_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[15] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[15] ));
 sg13g2_buf_2 place10038 (.A(_11003_),
    .X(net10038));
 sg13g2_buf_2 place10015 (.A(net10014),
    .X(net10015));
 sg13g2_xnor2_1 _22189_ (.Y(_04414_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[14] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14] ));
 sg13g2_buf_16 clkbuf_leaf_355_clk (.X(clknet_leaf_355_clk),
    .A(clknet_8_124_0_clk));
 sg13g2_buf_16 clkbuf_leaf_353_clk (.X(clknet_leaf_353_clk),
    .A(clknet_8_118_0_clk));
 sg13g2_nand2b_1 _22192_ (.Y(_04417_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[13] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13] ));
 sg13g2_nand3_1 _22193_ (.B(_04414_),
    .C(_04417_),
    .A(_04411_),
    .Y(_04418_));
 sg13g2_buf_2 place9997 (.A(net9996),
    .X(net9997));
 sg13g2_buf_2 place10013 (.A(_11164_),
    .X(net10013));
 sg13g2_xor2_1 _22196_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[12] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[12] ),
    .X(_04421_));
 sg13g2_inv_4 _22197_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[8] ),
    .Y(_04422_));
 sg13g2_buf_2 place10008 (.A(net10007),
    .X(net10008));
 sg13g2_nand2b_1 _22199_ (.Y(_04424_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[9] ));
 sg13g2_o21ai_1 _22200_ (.B1(_04424_),
    .Y(_04425_),
    .A1(_04422_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[8] ));
 sg13g2_nor2b_1 _22201_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[13] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13] ),
    .Y(_04426_));
 sg13g2_a21o_1 _22202_ (.A2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[8] ),
    .A1(_04422_),
    .B1(_04426_),
    .X(_04427_));
 sg13g2_nor4_1 _22203_ (.A(_04418_),
    .B(_04421_),
    .C(_04425_),
    .D(_04427_),
    .Y(_04428_));
 sg13g2_and2_1 _22204_ (.A(_04408_),
    .B(_04428_),
    .X(_04429_));
 sg13g2_buf_2 place10014 (.A(net10013),
    .X(net10014));
 sg13g2_buf_16 clkbuf_leaf_356_clk (.X(clknet_leaf_356_clk),
    .A(clknet_8_124_0_clk));
 sg13g2_xor2_1 _22207_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[2] ),
    .X(_04432_));
 sg13g2_buf_2 place10006 (.A(net10005),
    .X(net10006));
 sg13g2_buf_2 place9990 (.A(_05426_),
    .X(net9990));
 sg13g2_nor2b_1 _22210_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[5] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[5] ),
    .Y(_04435_));
 sg13g2_buf_2 place9998 (.A(_11324_),
    .X(net9998));
 sg13g2_buf_2 place10005 (.A(net10004),
    .X(net10005));
 sg13g2_xnor2_1 _22213_ (.Y(_04438_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[7] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[7] ));
 sg13g2_buf_16 clkbuf_leaf_365_clk (.X(clknet_leaf_365_clk),
    .A(clknet_8_126_0_clk));
 sg13g2_buf_2 place9995 (.A(net9994),
    .X(net9995));
 sg13g2_xnor2_1 _22216_ (.Y(_04441_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[6] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[6] ));
 sg13g2_nand2b_1 _22217_ (.Y(_04442_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[5] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[5] ));
 sg13g2_nand3_1 _22218_ (.B(_04441_),
    .C(_04442_),
    .A(_04438_),
    .Y(_04443_));
 sg13g2_buf_2 place9996 (.A(net9994),
    .X(net9996));
 sg13g2_xnor2_1 _22220_ (.Y(_04445_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[0] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[0] ));
 sg13g2_buf_2 place9989 (.A(_05426_),
    .X(net9989));
 sg13g2_buf_2 place9987 (.A(_05789_),
    .X(net9987));
 sg13g2_nand2b_1 _22223_ (.Y(_04448_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[4] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[4] ));
 sg13g2_inv_2 _22224_ (.Y(_04449_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[4] ));
 sg13g2_nand2_1 _22225_ (.Y(_04450_),
    .A(_04449_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[4] ));
 sg13g2_buf_16 clkbuf_leaf_362_clk (.X(clknet_leaf_362_clk),
    .A(clknet_8_125_0_clk));
 sg13g2_buf_16 clkbuf_leaf_360_clk (.X(clknet_leaf_360_clk),
    .A(clknet_8_125_0_clk));
 sg13g2_xor2_1 _22228_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[1] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[1] ),
    .X(_04453_));
 sg13g2_buf_16 clkbuf_leaf_357_clk (.X(clknet_leaf_357_clk),
    .A(clknet_8_125_0_clk));
 sg13g2_buf_16 clkbuf_leaf_359_clk (.X(clknet_leaf_359_clk),
    .A(clknet_8_119_0_clk));
 sg13g2_xor2_1 _22231_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[3] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[3] ),
    .X(_04456_));
 sg13g2_nor2_1 _22232_ (.A(_04453_),
    .B(_04456_),
    .Y(_04457_));
 sg13g2_nand4_1 _22233_ (.B(_04448_),
    .C(_04450_),
    .A(_04445_),
    .Y(_04458_),
    .D(_04457_));
 sg13g2_nor4_1 _22234_ (.A(_04432_),
    .B(_04435_),
    .C(_04443_),
    .D(_04458_),
    .Y(_04459_));
 sg13g2_nand3b_1 _22235_ (.B(_04429_),
    .C(_04459_),
    .Y(_04460_),
    .A_N(_04398_));
 sg13g2_buf_16 clkbuf_leaf_358_clk (.X(clknet_leaf_358_clk),
    .A(clknet_8_119_0_clk));
 sg13g2_inv_2 _22237_ (.Y(_04462_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[3] ));
 sg13g2_inv_1 _22238_ (.Y(_04463_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[2] ));
 sg13g2_nor2_1 _22239_ (.A(_04463_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2] ),
    .Y(_04464_));
 sg13g2_inv_2 _22240_ (.Y(_04465_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[1] ));
 sg13g2_nor2b_1 _22241_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[0] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[0] ),
    .Y(_04466_));
 sg13g2_nand2_1 _22242_ (.Y(_04467_),
    .A(_04465_),
    .B(_04466_));
 sg13g2_o21ai_1 _22243_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[1] ),
    .Y(_04468_),
    .A1(_04465_),
    .A2(_04466_));
 sg13g2_a22oi_1 _22244_ (.Y(_04469_),
    .B1(_04467_),
    .B2(_04468_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2] ),
    .A1(_04463_));
 sg13g2_nor3_1 _22245_ (.A(_04462_),
    .B(_04464_),
    .C(_04469_),
    .Y(_04470_));
 sg13g2_o21ai_1 _22246_ (.B1(_04462_),
    .Y(_04471_),
    .A1(_04464_),
    .A2(_04469_));
 sg13g2_a21oi_1 _22247_ (.A1(_04449_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[4] ),
    .Y(_04472_),
    .B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[3] ));
 sg13g2_nand2b_1 _22248_ (.Y(_04473_),
    .B(_04448_),
    .A_N(_04435_));
 sg13g2_a221oi_1 _22249_ (.B2(_04472_),
    .C1(_04473_),
    .B1(_04471_),
    .A1(_04450_),
    .Y(_04474_),
    .A2(_04470_));
 sg13g2_nor2b_1 _22250_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[6] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[6] ),
    .Y(_04475_));
 sg13g2_nand2_2 _22251_ (.Y(_04476_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[7] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[6] ));
 sg13g2_o21ai_1 _22252_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[7] ),
    .Y(_04477_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[6] ),
    .A2(_04476_));
 sg13g2_o21ai_1 _22253_ (.B1(_04477_),
    .Y(_04478_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[7] ),
    .A2(_04475_));
 sg13g2_o21ai_1 _22254_ (.B1(_04478_),
    .Y(_04479_),
    .A1(_04443_),
    .A2(_04474_));
 sg13g2_and2_1 _22255_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[11] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[10] ),
    .X(_04480_));
 sg13g2_buf_16 clkbuf_leaf_366_clk (.X(clknet_leaf_366_clk),
    .A(clknet_8_126_0_clk));
 sg13g2_inv_1 _22257_ (.Y(_04482_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[10] ));
 sg13g2_inv_1 _22258_ (.Y(_04483_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[11] ));
 sg13g2_nand2b_1 _22259_ (.Y(_04484_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[10] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[10] ));
 sg13g2_a21oi_1 _22260_ (.A1(_04483_),
    .A2(_04484_),
    .Y(_04485_),
    .B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[11] ));
 sg13g2_a221oi_1 _22261_ (.B2(_04482_),
    .C1(_04485_),
    .B1(_04480_),
    .A1(_04408_),
    .Y(_04486_),
    .A2(_04425_));
 sg13g2_inv_1 _22262_ (.Y(_04487_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[12] ));
 sg13g2_o21ai_1 _22263_ (.B1(_04487_),
    .Y(_04488_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[12] ),
    .A2(_04486_));
 sg13g2_nand2_1 _22264_ (.Y(_04489_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[12] ),
    .B(_04486_));
 sg13g2_a21oi_1 _22265_ (.A1(_04488_),
    .A2(_04489_),
    .Y(_04490_),
    .B1(_04426_));
 sg13g2_nor2b_1 _22266_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[14] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14] ),
    .Y(_04491_));
 sg13g2_nand2_1 _22267_ (.Y(_04492_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[15] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14] ));
 sg13g2_o21ai_1 _22268_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[15] ),
    .Y(_04493_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[14] ),
    .A2(_04492_));
 sg13g2_o21ai_1 _22269_ (.B1(_04493_),
    .Y(_04494_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[15] ),
    .A2(_04491_));
 sg13g2_o21ai_1 _22270_ (.B1(_04494_),
    .Y(_04495_),
    .A1(_04418_),
    .A2(_04490_));
 sg13g2_a21oi_1 _22271_ (.A1(_04429_),
    .A2(_04479_),
    .Y(_04496_),
    .B1(_04495_));
 sg13g2_nand2_1 _22272_ (.Y(_04497_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[31] ),
    .B(_04344_));
 sg13g2_inv_2 _22273_ (.Y(_04498_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[31] ));
 sg13g2_o21ai_1 _22274_ (.B1(_04498_),
    .Y(_04499_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[31] ),
    .A2(_04344_));
 sg13g2_nand2b_1 _22275_ (.Y(_04500_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[18] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[18] ));
 sg13g2_nand2b_1 _22276_ (.Y(_04501_),
    .B(_04500_),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[19] ));
 sg13g2_nand2_2 _22277_ (.Y(_04502_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[19] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[18] ));
 sg13g2_o21ai_1 _22278_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[19] ),
    .Y(_04503_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[18] ),
    .A2(_04502_));
 sg13g2_a22oi_1 _22279_ (.Y(_04504_),
    .B1(_04501_),
    .B2(_04503_),
    .A2(_04396_),
    .A1(_04386_));
 sg13g2_inv_2 _22280_ (.Y(_04505_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[20] ));
 sg13g2_o21ai_1 _22281_ (.B1(_04505_),
    .Y(_04506_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[20] ),
    .A2(_04504_));
 sg13g2_nand2_1 _22282_ (.Y(_04507_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[20] ),
    .B(_04504_));
 sg13g2_a21oi_1 _22283_ (.A1(_04506_),
    .A2(_04507_),
    .Y(_04508_),
    .B1(_04387_));
 sg13g2_nand2_1 _22284_ (.Y(_04509_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[23] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22] ));
 sg13g2_o21ai_1 _22285_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[23] ),
    .Y(_04510_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[22] ),
    .A2(_04509_));
 sg13g2_o21ai_1 _22286_ (.B1(_04510_),
    .Y(_04511_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[23] ),
    .A2(_04367_));
 sg13g2_o21ai_1 _22287_ (.B1(_04511_),
    .Y(_04512_),
    .A1(_04375_),
    .A2(_04508_));
 sg13g2_and2_1 _22288_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[27] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[26] ),
    .X(_04513_));
 sg13g2_buf_2 place9992 (.A(net9991),
    .X(net9992));
 sg13g2_inv_1 _22290_ (.Y(_04515_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[26] ));
 sg13g2_inv_1 _22291_ (.Y(_04516_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[27] ));
 sg13g2_nand2b_1 _22292_ (.Y(_04517_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[26] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[26] ));
 sg13g2_a21oi_1 _22293_ (.A1(_04516_),
    .A2(_04517_),
    .Y(_04518_),
    .B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[27] ));
 sg13g2_a221oi_1 _22294_ (.B2(_04515_),
    .C1(_04518_),
    .B1(_04513_),
    .A1(_04341_),
    .Y(_04519_),
    .A2(_04360_));
 sg13g2_nor2_1 _22295_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[28] ),
    .B(_04519_),
    .Y(_04520_));
 sg13g2_nand2_1 _22296_ (.Y(_04521_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[28] ),
    .B(_04519_));
 sg13g2_o21ai_1 _22297_ (.B1(_04521_),
    .Y(_04522_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[28] ),
    .A2(_04520_));
 sg13g2_a21oi_1 _22298_ (.A1(_04361_),
    .A2(_04522_),
    .Y(_04523_),
    .B1(_04353_));
 sg13g2_a221oi_1 _22299_ (.B2(_04364_),
    .C1(_04523_),
    .B1(_04512_),
    .A1(_04497_),
    .Y(_04524_),
    .A2(_04499_));
 sg13g2_o21ai_1 _22300_ (.B1(_04524_),
    .Y(_04525_),
    .A1(_04398_),
    .A2(_04496_));
 sg13g2_buf_2 place10029 (.A(_11043_),
    .X(net10029));
 sg13g2_nand2_2 _22302_ (.Y(_04527_),
    .A(_04460_),
    .B(_04525_));
 sg13g2_buf_2 place9991 (.A(net9990),
    .X(net9991));
 sg13g2_buf_2 place9986 (.A(_07054_),
    .X(net9986));
 sg13g2_buf_2 place10027 (.A(net10025),
    .X(net10027));
 sg13g2_nand3_1 _22306_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfering ),
    .C(_00096_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.start_bit ),
    .Y(_04531_));
 sg13g2_buf_2 place10012 (.A(net10011),
    .X(net10012));
 sg13g2_buf_2 place10030 (.A(net10029),
    .X(net10030));
 sg13g2_nor2b_1 _22309_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[1] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[1] ),
    .Y(_04534_));
 sg13g2_nand2b_1 _22310_ (.Y(_04535_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[1] ),
    .A_N(net10733));
 sg13g2_buf_2 place10020 (.A(net10018),
    .X(net10020));
 sg13g2_xor2_1 _22312_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[2] ),
    .X(_04537_));
 sg13g2_buf_2 place9988 (.A(net9987),
    .X(net9988));
 sg13g2_xor2_1 _22314_ (.B(net10734),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[0] ),
    .X(_04539_));
 sg13g2_nand2b_2 _22315_ (.Y(_04540_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfering ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.start_bit ));
 sg13g2_nor4_1 _22316_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.stop_bit ),
    .B(_04537_),
    .C(_04539_),
    .D(_04540_),
    .Y(_04541_));
 sg13g2_nand3b_1 _22317_ (.B(_04535_),
    .C(_04541_),
    .Y(_04542_),
    .A_N(_04534_));
 sg13g2_or2_1 _22318_ (.X(_04543_),
    .B(_04542_),
    .A(_04460_));
 sg13g2_buf_16 clkbuf_leaf_367_clk (.X(clknet_leaf_367_clk),
    .A(clknet_8_121_0_clk));
 sg13g2_nand2_1 _22320_ (.Y(_04545_),
    .A(_04531_),
    .B(_04543_));
 sg13g2_inv_8 _22321_ (.Y(_04546_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout ));
 sg13g2_nor3_1 _22322_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_ready ),
    .B(_04546_),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_done ),
    .Y(_04547_));
 sg13g2_nand2_2 _22323_ (.Y(_04548_),
    .A(_08412_),
    .B(_04547_));
 sg13g2_nand2_2 _22324_ (.Y(_04549_),
    .A(net11056),
    .B(_04548_));
 sg13g2_and2_1 _22325_ (.A(_07881_),
    .B(_07895_),
    .X(_04550_));
 sg13g2_buf_2 place10007 (.A(net10004),
    .X(net10007));
 sg13g2_nand2_2 _22327_ (.Y(_04552_),
    .A(_07882_),
    .B(_04550_));
 sg13g2_nor3_2 _22328_ (.A(\u_ac_controller_soc_inst.cbus_wstrb[1] ),
    .B(\u_ac_controller_soc_inst.cbus_wstrb[2] ),
    .C(\u_ac_controller_soc_inst.cbus_wstrb[3] ),
    .Y(_04553_));
 sg13g2_nand2b_2 _22329_ (.Y(_04554_),
    .B(_04553_),
    .A_N(\u_ac_controller_soc_inst.cbus_wstrb[0] ));
 sg13g2_buf_2 place9994 (.A(_11324_),
    .X(net9994));
 sg13g2_nand2b_2 _22331_ (.Y(_04556_),
    .B(_04554_),
    .A_N(_08410_));
 sg13g2_buf_2 place9983 (.A(net9982),
    .X(net9983));
 sg13g2_nor4_2 _22333_ (.A(net10606),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_ready ),
    .C(_04552_),
    .Y(_04558_),
    .D(_04556_));
 sg13g2_nor2b_2 _22334_ (.A(\u_ac_controller_soc_inst.cbus_wstrb[0] ),
    .B_N(_04553_),
    .Y(_04559_));
 sg13g2_nor4_1 _22335_ (.A(net10615),
    .B(net10617),
    .C(net10606),
    .D(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_ready ),
    .Y(_04560_));
 sg13g2_nor4_1 _22336_ (.A(net10613),
    .B(net10614),
    .C(net10612),
    .D(\u_ac_controller_soc_inst.cbus_addr[9] ),
    .Y(_04561_));
 sg13g2_nor2_2 _22337_ (.A(net10618),
    .B(net10459),
    .Y(_04562_));
 sg13g2_nand4_1 _22338_ (.B(_04560_),
    .C(_04561_),
    .A(_04559_),
    .Y(_04563_),
    .D(_04562_));
 sg13g2_buf_2 place10018 (.A(_11164_),
    .X(net10018));
 sg13g2_nor3_2 _22340_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync ),
    .B(_08410_),
    .C(_04563_),
    .Y(_04565_));
 sg13g2_o21ai_1 _22341_ (.B1(_00097_),
    .Y(_04566_),
    .A1(_04558_),
    .A2(_04565_));
 sg13g2_buf_2 place10019 (.A(net10018),
    .X(net10019));
 sg13g2_nand2b_2 _22343_ (.Y(_04568_),
    .B(_04566_),
    .A_N(_04549_));
 sg13g2_buf_2 place9982 (.A(_09877_),
    .X(net9982));
 sg13g2_a21o_2 _22345_ (.A2(_04545_),
    .A1(_04527_),
    .B1(_04568_),
    .X(_04570_));
 sg13g2_buf_2 place10017 (.A(net10016),
    .X(net10017));
 sg13g2_nor2_2 _22347_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.stop_bit ),
    .B(_04540_),
    .Y(_04572_));
 sg13g2_inv_4 _22348_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2] ),
    .Y(_04573_));
 sg13g2_inv_4 _22349_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[0] ),
    .Y(_04574_));
 sg13g2_nor2_1 _22350_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[0] ),
    .B(_04574_),
    .Y(_04575_));
 sg13g2_a21oi_1 _22351_ (.A1(_04535_),
    .A2(_04575_),
    .Y(_04576_),
    .B1(_04534_));
 sg13g2_o21ai_1 _22352_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[2] ),
    .Y(_04577_),
    .A1(_04573_),
    .A2(_04576_));
 sg13g2_nand2_1 _22353_ (.Y(_04578_),
    .A(_04573_),
    .B(_04576_));
 sg13g2_nand2_2 _22354_ (.Y(_04579_),
    .A(_04577_),
    .B(_04578_));
 sg13g2_nand2_2 _22355_ (.Y(_04580_),
    .A(_04572_),
    .B(_04579_));
 sg13g2_or2_1 _22356_ (.X(_04581_),
    .B(_04540_),
    .A(_00096_));
 sg13g2_buf_2 place9985 (.A(_09877_),
    .X(net9985));
 sg13g2_and2_1 _22358_ (.A(_04580_),
    .B(_04581_),
    .X(_04583_));
 sg13g2_buf_2 place9984 (.A(net9983),
    .X(net9984));
 sg13g2_o21ai_1 _22360_ (.B1(_04527_),
    .Y(_04585_),
    .A1(_04525_),
    .A2(_04580_));
 sg13g2_or2_1 _22361_ (.X(_04586_),
    .B(_04585_),
    .A(_04583_));
 sg13g2_buf_16 clkbuf_leaf_369_clk (.X(clknet_leaf_369_clk),
    .A(clknet_8_126_0_clk));
 sg13g2_nor3_1 _22363_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[0] ),
    .B(_04460_),
    .C(_04580_),
    .Y(_04588_));
 sg13g2_a21oi_1 _22364_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[0] ),
    .A2(_04586_),
    .Y(_04589_),
    .B1(_04588_));
 sg13g2_nor2_1 _22365_ (.A(_04570_),
    .B(_04589_),
    .Y(_00401_));
 sg13g2_nor2_1 _22366_ (.A(_04460_),
    .B(_04580_),
    .Y(_04590_));
 sg13g2_buf_16 clkbuf_leaf_368_clk (.X(clknet_leaf_368_clk),
    .A(clknet_8_121_0_clk));
 sg13g2_nor2_2 _22368_ (.A(_04574_),
    .B(net10733),
    .Y(_04592_));
 sg13g2_nand2_1 _22369_ (.Y(_04593_),
    .A(_04590_),
    .B(_04592_));
 sg13g2_o21ai_1 _22370_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[1] ),
    .Y(_04594_),
    .A1(_04588_),
    .A2(_04586_));
 sg13g2_a21oi_1 _22371_ (.A1(_04593_),
    .A2(_04594_),
    .Y(_00402_),
    .B1(_04570_));
 sg13g2_and2_1 _22372_ (.A(net10734),
    .B(net10733),
    .X(_04595_));
 sg13g2_buf_2 place9980 (.A(net9979),
    .X(net9980));
 sg13g2_xnor2_1 _22374_ (.Y(_04597_),
    .A(_00136_),
    .B(_04595_));
 sg13g2_a22oi_1 _22375_ (.Y(_04598_),
    .B1(_04597_),
    .B2(_04590_),
    .A2(_04586_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2] ));
 sg13g2_nor2_1 _22376_ (.A(_04570_),
    .B(_04598_),
    .Y(_00403_));
 sg13g2_inv_1 _22377_ (.Y(_04599_),
    .A(_04525_));
 sg13g2_and3_1 _22378_ (.X(_04600_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.start_bit ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfering ),
    .C(_00096_));
 sg13g2_nand2_1 _22379_ (.Y(_04601_),
    .A(_00135_),
    .B(_04600_));
 sg13g2_o21ai_1 _22380_ (.B1(_04601_),
    .Y(_04602_),
    .A1(net10732),
    .A2(_04583_));
 sg13g2_nand2_1 _22381_ (.Y(_04603_),
    .A(_04531_),
    .B(_04583_));
 sg13g2_nand2_2 _22382_ (.Y(_04604_),
    .A(_04527_),
    .B(_04603_));
 sg13g2_a22oi_1 _22383_ (.Y(_04605_),
    .B1(_04604_),
    .B2(net10732),
    .A2(_04602_),
    .A1(_04599_));
 sg13g2_nor2_1 _22384_ (.A(_04568_),
    .B(_04605_),
    .Y(_00404_));
 sg13g2_a21oi_1 _22385_ (.A1(_04531_),
    .A2(_04583_),
    .Y(_04606_),
    .B1(_04460_));
 sg13g2_or2_1 _22386_ (.X(_04607_),
    .B(_04606_),
    .A(_04568_));
 sg13g2_buf_2 place10032 (.A(_11003_),
    .X(net10032));
 sg13g2_buf_2 place9978 (.A(_09894_),
    .X(net9978));
 sg13g2_nor2_1 _22389_ (.A(_04449_),
    .B(_04462_),
    .Y(_04610_));
 sg13g2_nand4_1 _22390_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[1] ),
    .C(net10732),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2] ),
    .Y(_04611_),
    .D(_04610_));
 sg13g2_a221oi_1 _22391_ (.B2(_04583_),
    .C1(_04611_),
    .B1(_04531_),
    .A1(_04460_),
    .Y(_04612_),
    .A2(_04525_));
 sg13g2_buf_2 place10010 (.A(net10004),
    .X(net10010));
 sg13g2_and2_1 _22393_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[5] ),
    .B(_04612_),
    .X(_04614_));
 sg13g2_buf_2 place10009 (.A(net10007),
    .X(net10009));
 sg13g2_nor2_2 _22395_ (.A(_04422_),
    .B(_04476_),
    .Y(_04616_));
 sg13g2_nand3_1 _22396_ (.B(_04614_),
    .C(_04616_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9] ),
    .Y(_04617_));
 sg13g2_xor2_1 _22397_ (.B(_04617_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[10] ),
    .X(_04618_));
 sg13g2_nor2_1 _22398_ (.A(net9709),
    .B(_04618_),
    .Y(_00405_));
 sg13g2_nand4_1 _22399_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9] ),
    .C(_04614_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[10] ),
    .Y(_04619_),
    .D(_04616_));
 sg13g2_xnor2_1 _22400_ (.Y(_04620_),
    .A(_04483_),
    .B(_04619_));
 sg13g2_nor2_1 _22401_ (.A(net9709),
    .B(_04620_),
    .Y(_00406_));
 sg13g2_nand4_1 _22402_ (.B(_04480_),
    .C(_04614_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9] ),
    .Y(_04621_),
    .D(_04616_));
 sg13g2_xnor2_1 _22403_ (.Y(_04622_),
    .A(_04487_),
    .B(_04621_));
 sg13g2_nor2_1 _22404_ (.A(net9708),
    .B(_04622_),
    .Y(_00407_));
 sg13g2_and2_1 _22405_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[12] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9] ),
    .X(_04623_));
 sg13g2_and4_1 _22406_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[5] ),
    .B(_04480_),
    .C(_04616_),
    .D(_04623_),
    .X(_04624_));
 sg13g2_and2_1 _22407_ (.A(_04612_),
    .B(_04624_),
    .X(_04625_));
 sg13g2_buf_2 place9993 (.A(_11462_),
    .X(net9993));
 sg13g2_xnor2_1 _22409_ (.Y(_04627_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13] ),
    .B(_04625_));
 sg13g2_nor2_1 _22410_ (.A(net9709),
    .B(_04627_),
    .Y(_00408_));
 sg13g2_nand2_1 _22411_ (.Y(_04628_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13] ),
    .B(_04625_));
 sg13g2_xor2_1 _22412_ (.B(_04628_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14] ),
    .X(_04629_));
 sg13g2_nor2_1 _22413_ (.A(net9709),
    .B(_04629_),
    .Y(_00409_));
 sg13g2_nand3_1 _22414_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13] ),
    .C(_04625_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14] ),
    .Y(_04630_));
 sg13g2_xor2_1 _22415_ (.B(_04630_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[15] ),
    .X(_04631_));
 sg13g2_nor2_1 _22416_ (.A(net9709),
    .B(_04631_),
    .Y(_00410_));
 sg13g2_nor2_1 _22417_ (.A(_04492_),
    .B(_04628_),
    .Y(_04632_));
 sg13g2_xnor2_1 _22418_ (.Y(_04633_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[16] ),
    .B(_04632_));
 sg13g2_nor2_1 _22419_ (.A(net9709),
    .B(_04633_),
    .Y(_00411_));
 sg13g2_and4_1 _22420_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[16] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[15] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14] ),
    .D(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13] ),
    .X(_04634_));
 sg13g2_nand2_1 _22421_ (.Y(_04635_),
    .A(_04625_),
    .B(_04634_));
 sg13g2_xor2_1 _22422_ (.B(_04635_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[17] ),
    .X(_04636_));
 sg13g2_nor2_1 _22423_ (.A(net9709),
    .B(_04636_),
    .Y(_00412_));
 sg13g2_and4_2 _22424_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[17] ),
    .B(_04612_),
    .C(_04624_),
    .D(_04634_),
    .X(_04637_));
 sg13g2_buf_2 place9979 (.A(net9978),
    .X(net9979));
 sg13g2_xnor2_1 _22426_ (.Y(_04639_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[18] ),
    .B(_04637_));
 sg13g2_nor2_1 _22427_ (.A(net9711),
    .B(_04639_),
    .Y(_00413_));
 sg13g2_buf_2 place10011 (.A(_11244_),
    .X(net10011));
 sg13g2_nand2_1 _22429_ (.Y(_04641_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[18] ),
    .B(_04637_));
 sg13g2_xor2_1 _22430_ (.B(_04641_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[19] ),
    .X(_04642_));
 sg13g2_nor2_1 _22431_ (.A(net9711),
    .B(_04642_),
    .Y(_00414_));
 sg13g2_and2_1 _22432_ (.A(_04527_),
    .B(_04603_),
    .X(_04643_));
 sg13g2_buf_2 place9981 (.A(_09894_),
    .X(net9981));
 sg13g2_nand2_1 _22434_ (.Y(_04645_),
    .A(net10732),
    .B(_04643_));
 sg13g2_xnor2_1 _22435_ (.Y(_04646_),
    .A(_04465_),
    .B(_04645_));
 sg13g2_nor2_1 _22436_ (.A(net9708),
    .B(_04646_),
    .Y(_00415_));
 sg13g2_nand2b_1 _22437_ (.Y(_04647_),
    .B(_04637_),
    .A_N(_04502_));
 sg13g2_xnor2_1 _22438_ (.Y(_04648_),
    .A(_04505_),
    .B(_04647_));
 sg13g2_nor2_1 _22439_ (.A(net9711),
    .B(_04648_),
    .Y(_00416_));
 sg13g2_or2_1 _22440_ (.X(_04649_),
    .B(_04647_),
    .A(_04505_));
 sg13g2_xnor2_1 _22441_ (.Y(_04650_),
    .A(_04370_),
    .B(_04649_));
 sg13g2_nor2_1 _22442_ (.A(net9711),
    .B(_04650_),
    .Y(_00417_));
 sg13g2_nor3_2 _22443_ (.A(_04370_),
    .B(_04505_),
    .C(_04502_),
    .Y(_04651_));
 sg13g2_nand2_1 _22444_ (.Y(_04652_),
    .A(_04637_),
    .B(_04651_));
 sg13g2_xor2_1 _22445_ (.B(_04652_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22] ),
    .X(_04653_));
 sg13g2_nor2_1 _22446_ (.A(net9711),
    .B(_04653_),
    .Y(_00418_));
 sg13g2_nand3_1 _22447_ (.B(_04637_),
    .C(_04651_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22] ),
    .Y(_04654_));
 sg13g2_xor2_1 _22448_ (.B(_04654_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[23] ),
    .X(_04655_));
 sg13g2_nor2_1 _22449_ (.A(net9711),
    .B(_04655_),
    .Y(_00419_));
 sg13g2_nand3_1 _22450_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22] ),
    .C(_04651_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[23] ),
    .Y(_04656_));
 sg13g2_inv_1 _22451_ (.Y(_04657_),
    .A(_04656_));
 sg13g2_and2_1 _22452_ (.A(_04637_),
    .B(_04657_),
    .X(_04658_));
 sg13g2_xnor2_1 _22453_ (.Y(_04659_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[24] ),
    .B(_04658_));
 sg13g2_nor2_1 _22454_ (.A(net9711),
    .B(_04659_),
    .Y(_00420_));
 sg13g2_nand2_1 _22455_ (.Y(_04660_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[24] ),
    .B(_04658_));
 sg13g2_xor2_1 _22456_ (.B(_04660_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[25] ),
    .X(_04661_));
 sg13g2_nor2_1 _22457_ (.A(net9711),
    .B(_04661_),
    .Y(_00421_));
 sg13g2_and4_2 _22458_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[25] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[24] ),
    .C(_04637_),
    .D(_04657_),
    .X(_04662_));
 sg13g2_buf_16 clkbuf_leaf_371_clk (.X(clknet_leaf_371_clk),
    .A(clknet_8_121_0_clk));
 sg13g2_xnor2_1 _22460_ (.Y(_04664_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[26] ),
    .B(_04662_));
 sg13g2_nor2_1 _22461_ (.A(net9710),
    .B(_04664_),
    .Y(_00422_));
 sg13g2_nand2_1 _22462_ (.Y(_04665_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[26] ),
    .B(_04662_));
 sg13g2_xnor2_1 _22463_ (.Y(_04666_),
    .A(_04516_),
    .B(_04665_));
 sg13g2_nor2_1 _22464_ (.A(net9710),
    .B(_04666_),
    .Y(_00423_));
 sg13g2_buf_16 clkbuf_leaf_370_clk (.X(clknet_leaf_370_clk),
    .A(clknet_8_124_0_clk));
 sg13g2_nand2_1 _22466_ (.Y(_04668_),
    .A(_04513_),
    .B(_04662_));
 sg13g2_xor2_1 _22467_ (.B(_04668_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[28] ),
    .X(_04669_));
 sg13g2_nor2_1 _22468_ (.A(net9710),
    .B(_04669_),
    .Y(_00424_));
 sg13g2_nand3_1 _22469_ (.B(_04513_),
    .C(_04662_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[28] ),
    .Y(_04670_));
 sg13g2_xnor2_1 _22470_ (.Y(_04671_),
    .A(_04349_),
    .B(_04670_));
 sg13g2_nor2_1 _22471_ (.A(net9710),
    .B(_04671_),
    .Y(_00425_));
 sg13g2_nand3_1 _22472_ (.B(net10732),
    .C(_04643_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[1] ),
    .Y(_04672_));
 sg13g2_xor2_1 _22473_ (.B(_04672_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2] ),
    .X(_04673_));
 sg13g2_nor2_1 _22474_ (.A(net9708),
    .B(_04673_),
    .Y(_00426_));
 sg13g2_nand4_1 _22475_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[28] ),
    .C(_04513_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[29] ),
    .Y(_04674_),
    .D(_04662_));
 sg13g2_xnor2_1 _22476_ (.Y(_04675_),
    .A(_04345_),
    .B(_04674_));
 sg13g2_nor2_1 _22477_ (.A(net9710),
    .B(_04675_),
    .Y(_00427_));
 sg13g2_o21ai_1 _22478_ (.B1(_04498_),
    .Y(_04676_),
    .A1(_04345_),
    .A2(_04674_));
 sg13g2_nor2b_1 _22479_ (.A(net9710),
    .B_N(_04676_),
    .Y(_00428_));
 sg13g2_nand4_1 _22480_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[1] ),
    .C(net10732),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2] ),
    .Y(_04677_),
    .D(_04643_));
 sg13g2_xnor2_1 _22481_ (.Y(_04678_),
    .A(_04462_),
    .B(_04677_));
 sg13g2_nor2_1 _22482_ (.A(_04607_),
    .B(_04678_),
    .Y(_00429_));
 sg13g2_nor2_1 _22483_ (.A(_04462_),
    .B(_04677_),
    .Y(_04679_));
 sg13g2_xnor2_1 _22484_ (.Y(_04680_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[4] ),
    .B(_04679_));
 sg13g2_nor2_1 _22485_ (.A(_04607_),
    .B(_04680_),
    .Y(_00430_));
 sg13g2_xnor2_1 _22486_ (.Y(_04681_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[5] ),
    .B(_04612_));
 sg13g2_nor2_1 _22487_ (.A(_04607_),
    .B(_04681_),
    .Y(_00431_));
 sg13g2_xnor2_1 _22488_ (.Y(_04682_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[6] ),
    .B(_04614_));
 sg13g2_nor2_1 _22489_ (.A(net9708),
    .B(_04682_),
    .Y(_00432_));
 sg13g2_nand2_1 _22490_ (.Y(_04683_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[6] ),
    .B(_04614_));
 sg13g2_xor2_1 _22491_ (.B(_04683_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[7] ),
    .X(_04684_));
 sg13g2_nor2_1 _22492_ (.A(net9708),
    .B(_04684_),
    .Y(_00433_));
 sg13g2_nand2b_1 _22493_ (.Y(_04685_),
    .B(_04614_),
    .A_N(_04476_));
 sg13g2_xnor2_1 _22494_ (.Y(_04686_),
    .A(_04422_),
    .B(_04685_));
 sg13g2_nor2_1 _22495_ (.A(net9708),
    .B(_04686_),
    .Y(_00434_));
 sg13g2_nand2_1 _22496_ (.Y(_04687_),
    .A(_04614_),
    .B(_04616_));
 sg13g2_xor2_1 _22497_ (.B(_04687_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9] ),
    .X(_04688_));
 sg13g2_nor2_1 _22498_ (.A(net9709),
    .B(_04688_),
    .Y(_00435_));
 sg13g2_nand2_1 _22499_ (.Y(_04689_),
    .A(_04566_),
    .B(_04604_));
 sg13g2_mux4_1 _22500_ (.S0(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[0] ),
    .A0(net10605),
    .A1(\u_ac_controller_soc_inst.cbus_wdata[1] ),
    .A2(\u_ac_controller_soc_inst.cbus_wdata[2] ),
    .A3(\u_ac_controller_soc_inst.cbus_wdata[3] ),
    .S1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[1] ),
    .X(_04690_));
 sg13g2_mux4_1 _22501_ (.S0(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[0] ),
    .A0(\u_ac_controller_soc_inst.cbus_wdata[4] ),
    .A1(\u_ac_controller_soc_inst.cbus_wdata[5] ),
    .A2(\u_ac_controller_soc_inst.cbus_wdata[6] ),
    .A3(\u_ac_controller_soc_inst.cbus_wdata[7] ),
    .S1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[1] ),
    .X(_04691_));
 sg13g2_nand2b_1 _22502_ (.Y(_04692_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2] ),
    .A_N(_04691_));
 sg13g2_o21ai_1 _22503_ (.B1(_04692_),
    .Y(_04693_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2] ),
    .A2(_04690_));
 sg13g2_nand4_1 _22504_ (.B(_04543_),
    .C(_04579_),
    .A(_04572_),
    .Y(_04694_),
    .D(_04693_));
 sg13g2_a21oi_1 _22505_ (.A1(_04531_),
    .A2(_04694_),
    .Y(_04695_),
    .B1(_04556_));
 sg13g2_a22oi_1 _22506_ (.Y(_04696_),
    .B1(_04527_),
    .B2(_04695_),
    .A2(_04558_),
    .A1(_00097_));
 sg13g2_o21ai_1 _22507_ (.B1(_04696_),
    .Y(_04697_),
    .A1(ser_tx),
    .A2(_04689_));
 sg13g2_nand2b_1 _22508_ (.Y(_00447_),
    .B(_04697_),
    .A_N(_04549_));
 sg13g2_o21ai_1 _22509_ (.B1(_04566_),
    .Y(_04698_),
    .A1(_04525_),
    .A2(_04531_));
 sg13g2_a21oi_1 _22510_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.start_bit ),
    .A2(_04604_),
    .Y(_04699_),
    .B1(_04698_));
 sg13g2_nor2_1 _22511_ (.A(_04549_),
    .B(_04699_),
    .Y(_00448_));
 sg13g2_o21ai_1 _22512_ (.B1(_04460_),
    .Y(_04700_),
    .A1(_04525_),
    .A2(_04581_));
 sg13g2_inv_1 _22513_ (.Y(_04701_),
    .A(_04700_));
 sg13g2_o21ai_1 _22514_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.stop_bit ),
    .Y(_04702_),
    .A1(_04583_),
    .A2(_04701_));
 sg13g2_nand2b_1 _22515_ (.Y(_04703_),
    .B(_04580_),
    .A_N(_04581_));
 sg13g2_o21ai_1 _22516_ (.B1(_04543_),
    .Y(_04704_),
    .A1(_04525_),
    .A2(_04703_));
 sg13g2_inv_1 _22517_ (.Y(_04705_),
    .A(_04704_));
 sg13g2_a221oi_1 _22518_ (.B2(_04705_),
    .C1(_04568_),
    .B1(_04702_),
    .A1(_04527_),
    .Y(_00449_),
    .A2(_04600_));
 sg13g2_buf_2 place9974 (.A(_10119_),
    .X(net9974));
 sg13g2_buf_2 place10084 (.A(_10568_),
    .X(net10084));
 sg13g2_buf_2 place9999 (.A(net9998),
    .X(net9999));
 sg13g2_nand4_1 _22522_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[16] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[15] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[17] ),
    .Y(_04709_),
    .D(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[14] ));
 sg13g2_nand2_1 _22523_ (.Y(_04710_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[19] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[18] ));
 sg13g2_nor2_1 _22524_ (.A(_04709_),
    .B(_04710_),
    .Y(_04711_));
 sg13g2_and3_2 _22525_ (.X(_04712_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[21] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[20] ),
    .C(_04711_));
 sg13g2_buf_2 place9977 (.A(net9976),
    .X(net9977));
 sg13g2_buf_2 place10003 (.A(net10002),
    .X(net10003));
 sg13g2_buf_2 place9976 (.A(net9975),
    .X(net9976));
 sg13g2_nand4_1 _22529_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[25] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[24] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[26] ),
    .Y(_04716_),
    .D(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[23] ));
 sg13g2_inv_1 _22530_ (.Y(_04717_),
    .A(_04716_));
 sg13g2_nand4_1 _22531_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[22] ),
    .C(_04712_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[27] ),
    .Y(_04718_),
    .D(_04717_));
 sg13g2_buf_2 place10000 (.A(net9999),
    .X(net10000));
 sg13g2_and2_1 _22533_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[7] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[6] ),
    .X(_04720_));
 sg13g2_buf_2 place9975 (.A(net9974),
    .X(net9975));
 sg13g2_nand4_1 _22535_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[9] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[8] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[10] ),
    .Y(_04722_),
    .D(_04720_));
 sg13g2_buf_2 place10002 (.A(net9998),
    .X(net10002));
 sg13g2_nand3_1 _22537_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[2] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[1] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[3] ),
    .Y(_04724_));
 sg13g2_buf_16 clkbuf_leaf_372_clk (.X(clknet_leaf_372_clk),
    .A(clknet_8_121_0_clk));
 sg13g2_buf_2 place9968 (.A(net9967),
    .X(net9968));
 sg13g2_nand2_1 _22540_ (.Y(_04727_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[4] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[0] ));
 sg13g2_nor2_1 _22541_ (.A(_04724_),
    .B(_04727_),
    .Y(_04728_));
 sg13g2_nand2_2 _22542_ (.Y(_04729_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[5] ),
    .B(_04728_));
 sg13g2_buf_2 place9969 (.A(_10126_),
    .X(net9969));
 sg13g2_nand3_1 _22544_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[12] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[11] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[13] ),
    .Y(_04731_));
 sg13g2_nor3_2 _22545_ (.A(_04722_),
    .B(_04729_),
    .C(_04731_),
    .Y(_04732_));
 sg13g2_inv_2 _22546_ (.Y(_04733_),
    .A(_04732_));
 sg13g2_buf_2 place9967 (.A(net9965),
    .X(net9967));
 sg13g2_buf_2 place9971 (.A(net9970),
    .X(net9971));
 sg13g2_nand4_1 _22549_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[30] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[29] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[31] ),
    .Y(_04736_),
    .D(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[28] ));
 sg13g2_nor3_2 _22550_ (.A(_04718_),
    .B(_04733_),
    .C(_04736_),
    .Y(_04737_));
 sg13g2_and4_1 _22551_ (.A(net11049),
    .B(_00111_),
    .C(_04556_),
    .D(_04737_),
    .X(_00496_));
 sg13g2_nand2_1 _22552_ (.Y(_04738_),
    .A(net11052),
    .B(_11418_));
 sg13g2_a21oi_1 _22553_ (.A1(_08861_),
    .A2(_08304_),
    .Y(_01775_),
    .B1(_04738_));
 sg13g2_nand2_2 _22554_ (.Y(_04739_),
    .A(net10364),
    .B(net10661));
 sg13g2_nor2_2 _22555_ (.A(_08332_),
    .B(_04739_),
    .Y(_04740_));
 sg13g2_nor2b_1 _22556_ (.A(_04740_),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.mem_do_prefetch ),
    .Y(_04741_));
 sg13g2_a21oi_1 _22557_ (.A1(_00051_),
    .A2(_04740_),
    .Y(_04742_),
    .B1(_04741_));
 sg13g2_nor3_1 _22558_ (.A(net11014),
    .B(_08326_),
    .C(_04742_),
    .Y(_01821_));
 sg13g2_a22oi_1 _22559_ (.Y(_04743_),
    .B1(_07967_),
    .B2(_07964_),
    .A2(_07956_),
    .A1(net10610));
 sg13g2_nor2_1 _22560_ (.A(net11013),
    .B(_04743_),
    .Y(_01822_));
 sg13g2_nand2b_1 _22561_ (.Y(_04744_),
    .B(net10708),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.mem_do_prefetch ));
 sg13g2_o21ai_1 _22562_ (.B1(_04744_),
    .Y(_04745_),
    .A1(net10708),
    .A2(_04739_));
 sg13g2_nor2_1 _22563_ (.A(_08341_),
    .B(_08348_),
    .Y(_04746_));
 sg13g2_nor4_1 _22564_ (.A(_08390_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_do_prefetch ),
    .C(_08325_),
    .D(_04746_),
    .Y(_04747_));
 sg13g2_a21oi_1 _22565_ (.A1(_08390_),
    .A2(_04745_),
    .Y(_04748_),
    .B1(_04747_));
 sg13g2_nor2_1 _22566_ (.A(net10722),
    .B(net10714),
    .Y(_04749_));
 sg13g2_nor2_1 _22567_ (.A(\u_ac_controller_soc_inst.u_picorv32.is_lui_auipc_jal ),
    .B(\u_ac_controller_soc_inst.u_picorv32.is_jalr_addi_slti_sltiu_xori_ori_andi ),
    .Y(_04750_));
 sg13g2_nand4_1 _22568_ (.B(_00101_),
    .C(\u_ac_controller_soc_inst.u_picorv32.is_sll_srl_sra ),
    .A(net11052),
    .Y(_04751_),
    .D(_04750_));
 sg13g2_a21oi_1 _22569_ (.A1(_08343_),
    .A2(_04751_),
    .Y(_04752_),
    .B1(_08390_));
 sg13g2_a221oi_1 _22570_ (.B2(_00109_),
    .C1(_04752_),
    .B1(_04749_),
    .A1(net11051),
    .Y(_04753_),
    .A2(_11937_));
 sg13g2_mux2_1 _22571_ (.A0(\u_ac_controller_soc_inst.u_picorv32.mem_do_rinst ),
    .A1(_04748_),
    .S(_04753_),
    .X(_04754_));
 sg13g2_or4_1 _22572_ (.A(net10722),
    .B(net10714),
    .C(net10708),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpu_state[0] ),
    .X(_04755_));
 sg13g2_nor4_1 _22573_ (.A(_00102_),
    .B(_07972_),
    .C(_08865_),
    .D(_04755_),
    .Y(_04756_));
 sg13g2_a22oi_1 _22574_ (.Y(_04757_),
    .B1(_04756_),
    .B2(_08859_),
    .A2(_04754_),
    .A1(_07956_));
 sg13g2_nor2_1 _22575_ (.A(net11013),
    .B(_04757_),
    .Y(_01823_));
 sg13g2_nor4_1 _22576_ (.A(net10609),
    .B(net10695),
    .C(\u_ac_controller_soc_inst.u_picorv32.cpu_state[3] ),
    .D(_04755_),
    .Y(_04758_));
 sg13g2_a22oi_1 _22577_ (.Y(_04759_),
    .B1(_07967_),
    .B2(_04758_),
    .A2(_07956_),
    .A1(net10609));
 sg13g2_nor2_1 _22578_ (.A(net11013),
    .B(_04759_),
    .Y(_01824_));
 sg13g2_a21o_1 _22579_ (.A2(_08151_),
    .A1(_00098_),
    .B1(net10455),
    .X(_04760_));
 sg13g2_mux2_1 _22580_ (.A0(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[22] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_ddr ),
    .S(_08255_),
    .X(_04761_));
 sg13g2_nor2b_1 _22581_ (.A(_04760_),
    .B_N(_04761_),
    .Y(_02043_));
 sg13g2_buf_2 place9973 (.A(net9972),
    .X(net9973));
 sg13g2_nand2_1 _22583_ (.Y(_04763_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_qspi ),
    .B(_08255_));
 sg13g2_o21ai_1 _22584_ (.B1(_04763_),
    .Y(_04764_),
    .A1(_08264_),
    .A2(_08255_));
 sg13g2_nor2b_1 _22585_ (.A(_04760_),
    .B_N(_04764_),
    .Y(_02044_));
 sg13g2_a21oi_1 _22586_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[1] ),
    .A2(net9706),
    .Y(_04765_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_rd ));
 sg13g2_nor2_1 _22587_ (.A(net9653),
    .B(_04765_),
    .Y(_02045_));
 sg13g2_or2_1 _22588_ (.X(_04766_),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.state[8] ),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[11] ));
 sg13g2_or3_1 _22589_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[2] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.state[4] ),
    .C(_04766_),
    .X(_04767_));
 sg13g2_nor4_2 _22590_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[0] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.state[3] ),
    .C(_03746_),
    .Y(_04768_),
    .D(_04767_));
 sg13g2_nor2_1 _22591_ (.A(_00100_),
    .B(_08243_),
    .Y(_04769_));
 sg13g2_nor2_2 _22592_ (.A(_04768_),
    .B(_04769_),
    .Y(_04770_));
 sg13g2_nand3_1 _22593_ (.B(_04766_),
    .C(_04770_),
    .A(_03757_),
    .Y(_04771_));
 sg13g2_nand2_2 _22594_ (.Y(_04772_),
    .A(_03757_),
    .B(_04770_));
 sg13g2_nand2_1 _22595_ (.Y(_04773_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[0] ),
    .B(_04772_));
 sg13g2_a21oi_1 _22596_ (.A1(_04771_),
    .A2(_04773_),
    .Y(_02046_),
    .B1(net10455));
 sg13g2_a21oi_1 _22597_ (.A1(_03757_),
    .A2(_04770_),
    .Y(_04774_),
    .B1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[1] ));
 sg13g2_nor3_1 _22598_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[11] ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.state[5] ),
    .C(_04772_),
    .Y(_04775_));
 sg13g2_nor3_1 _22599_ (.A(net10455),
    .B(_04774_),
    .C(_04775_),
    .Y(_02047_));
 sg13g2_mux2_1 _22600_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.state[3] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[2] ),
    .S(_04772_),
    .X(_04776_));
 sg13g2_and2_1 _22601_ (.A(_08215_),
    .B(_04776_),
    .X(_02048_));
 sg13g2_nor3_1 _22602_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.state[0] ),
    .B(_03745_),
    .C(_04767_),
    .Y(_04777_));
 sg13g2_and3_1 _22603_ (.X(_04778_),
    .A(_07982_),
    .B(_08262_),
    .C(_04777_));
 sg13g2_nor4_1 _22604_ (.A(net10455),
    .B(net9705),
    .C(_04768_),
    .D(_04778_),
    .Y(_02049_));
 sg13g2_a21oi_1 _22605_ (.A1(_07742_),
    .A2(_03810_),
    .Y(_02073_),
    .B1(_08228_));
 sg13g2_nand2_2 _22606_ (.Y(_04779_),
    .A(_08171_),
    .B(_08571_));
 sg13g2_buf_2 place9972 (.A(net9969),
    .X(net9972));
 sg13g2_a22oi_1 _22608_ (.Y(_04781_),
    .B1(_08196_),
    .B2(_08197_),
    .A2(_08193_),
    .A1(net10465));
 sg13g2_o21ai_1 _22609_ (.B1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[0] ),
    .Y(_04782_),
    .A1(_04779_),
    .A2(net10260));
 sg13g2_o21ai_1 _22610_ (.B1(_04782_),
    .Y(_04783_),
    .A1(_04779_),
    .A2(_04781_));
 sg13g2_inv_1 _22611_ (.Y(_04784_),
    .A(_04783_));
 sg13g2_nor3_1 _22612_ (.A(_00095_),
    .B(_08222_),
    .C(_04784_),
    .Y(_02108_));
 sg13g2_a21oi_1 _22613_ (.A1(_08186_),
    .A2(_08197_),
    .Y(_04785_),
    .B1(net10465));
 sg13g2_or2_1 _22614_ (.X(_04786_),
    .B(_08199_),
    .A(_08186_));
 sg13g2_o21ai_1 _22615_ (.B1(_04786_),
    .Y(_04787_),
    .A1(_00091_),
    .A2(_04785_));
 sg13g2_a21oi_1 _22616_ (.A1(_08175_),
    .A2(net10260),
    .Y(_04788_),
    .B1(_04787_));
 sg13g2_nor2_1 _22617_ (.A(_04779_),
    .B(_04788_),
    .Y(_04789_));
 sg13g2_a21oi_1 _22618_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1] ),
    .A2(_04779_),
    .Y(_04790_),
    .B1(_04789_));
 sg13g2_nor3_1 _22619_ (.A(_00095_),
    .B(net9705),
    .C(_04790_),
    .Y(_02109_));
 sg13g2_xor2_1 _22620_ (.B(_08188_),
    .A(_00093_),
    .X(_04791_));
 sg13g2_nor2_1 _22621_ (.A(_08178_),
    .B(_08560_),
    .Y(_04792_));
 sg13g2_a21oi_1 _22622_ (.A1(_08560_),
    .A2(_04791_),
    .Y(_04793_),
    .B1(_04792_));
 sg13g2_nand2_1 _22623_ (.Y(_04794_),
    .A(net10464),
    .B(_08164_));
 sg13g2_o21ai_1 _22624_ (.B1(_04794_),
    .Y(_04795_),
    .A1(net10464),
    .A2(_04793_));
 sg13g2_nor2_1 _22625_ (.A(_04779_),
    .B(_04795_),
    .Y(_04796_));
 sg13g2_a21oi_1 _22626_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2] ),
    .A2(_04779_),
    .Y(_04797_),
    .B1(_04796_));
 sg13g2_nor3_1 _22627_ (.A(_00095_),
    .B(net9705),
    .C(_04797_),
    .Y(_02110_));
 sg13g2_nor2_2 _22628_ (.A(_08204_),
    .B(_08171_),
    .Y(_04798_));
 sg13g2_nor3_1 _22629_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk ),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_csb ),
    .C(_04798_),
    .Y(_04799_));
 sg13g2_a21oi_1 _22630_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk ),
    .A2(_04798_),
    .Y(_04800_),
    .B1(_04799_));
 sg13g2_nor3_1 _22631_ (.A(_00095_),
    .B(_08222_),
    .C(_04800_),
    .Y(_02117_));
 sg13g2_o21ai_1 _22632_ (.B1(_08240_),
    .Y(_04801_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.state[10] ),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.state[7] ));
 sg13g2_nor2b_1 _22633_ (.A(net9653),
    .B_N(_04801_),
    .Y(_02143_));
 sg13g2_nand2_2 _22634_ (.Y(_04802_),
    .A(_00106_),
    .B(_04553_));
 sg13g2_nand2_2 _22635_ (.Y(_04803_),
    .A(net10247),
    .B(_04802_));
 sg13g2_nor2_2 _22636_ (.A(net10606),
    .B(_04803_),
    .Y(_04804_));
 sg13g2_buf_2 place9965 (.A(_10126_),
    .X(net9965));
 sg13g2_nor3_1 _22638_ (.A(_00104_),
    .B(_00105_),
    .C(_07872_),
    .Y(_04806_));
 sg13g2_nand3_1 _22639_ (.B(_04550_),
    .C(_04806_),
    .A(net10246),
    .Y(_04807_));
 sg13g2_buf_2 place9970 (.A(net9969),
    .X(net9970));
 sg13g2_nand3b_1 _22641_ (.B(_08078_),
    .C(net10617),
    .Y(_04809_),
    .A_N(_04807_));
 sg13g2_buf_2 place9966 (.A(net9965),
    .X(net9966));
 sg13g2_nor3_2 _22643_ (.A(_08126_),
    .B(net10459),
    .C(_04809_),
    .Y(_04811_));
 sg13g2_buf_16 clkbuf_leaf_374_clk (.X(clknet_leaf_374_clk),
    .A(clknet_8_115_0_clk));
 sg13g2_nand2_2 _22645_ (.Y(_04813_),
    .A(_04804_),
    .B(_04811_));
 sg13g2_buf_2 place9957 (.A(net9955),
    .X(net9957));
 sg13g2_buf_2 place10026 (.A(net10025),
    .X(net10026));
 sg13g2_buf_2 place9955 (.A(_10213_),
    .X(net9955));
 sg13g2_nand2_2 _22649_ (.Y(_04817_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[0] ),
    .B(net10246));
 sg13g2_buf_2 place9963 (.A(net9962),
    .X(net9963));
 sg13g2_nor2_1 _22651_ (.A(net9786),
    .B(_04817_),
    .Y(_04819_));
 sg13g2_a21oi_1 _22652_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[0] ),
    .A2(net9786),
    .Y(_04820_),
    .B1(_04819_));
 sg13g2_nor2_1 _22653_ (.A(net10986),
    .B(_04820_),
    .Y(_00176_));
 sg13g2_buf_2 place9962 (.A(net9961),
    .X(net9962));
 sg13g2_nand2_2 _22655_ (.Y(_04822_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[10] ),
    .B(net10250));
 sg13g2_nor2_1 _22656_ (.A(net9790),
    .B(_04822_),
    .Y(_04823_));
 sg13g2_a21oi_1 _22657_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[10] ),
    .A2(net9790),
    .Y(_04824_),
    .B1(_04823_));
 sg13g2_nor2_1 _22658_ (.A(net10985),
    .B(_04824_),
    .Y(_00177_));
 sg13g2_nand2_2 _22659_ (.Y(_04825_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[11] ),
    .B(net10250));
 sg13g2_nor2_1 _22660_ (.A(net9790),
    .B(_04825_),
    .Y(_04826_));
 sg13g2_a21oi_1 _22661_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[11] ),
    .A2(net9790),
    .Y(_04827_),
    .B1(_04826_));
 sg13g2_nor2_1 _22662_ (.A(net11002),
    .B(_04827_),
    .Y(_00178_));
 sg13g2_nand2_2 _22663_ (.Y(_04828_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[12] ),
    .B(net10250));
 sg13g2_nor2_1 _22664_ (.A(net9788),
    .B(_04828_),
    .Y(_04829_));
 sg13g2_a21oi_1 _22665_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[12] ),
    .A2(net9788),
    .Y(_04830_),
    .B1(_04829_));
 sg13g2_nor2_1 _22666_ (.A(net10984),
    .B(_04830_),
    .Y(_00179_));
 sg13g2_buf_2 place9959 (.A(_10213_),
    .X(net9959));
 sg13g2_nand2_2 _22668_ (.Y(_04832_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[13] ),
    .B(net10250));
 sg13g2_nor2_1 _22669_ (.A(net9790),
    .B(_04832_),
    .Y(_04833_));
 sg13g2_a21oi_1 _22670_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[13] ),
    .A2(net9790),
    .Y(_04834_),
    .B1(_04833_));
 sg13g2_nor2_1 _22671_ (.A(net11002),
    .B(_04834_),
    .Y(_00180_));
 sg13g2_nand2_2 _22672_ (.Y(_04835_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[14] ),
    .B(net10248));
 sg13g2_nor2_1 _22673_ (.A(_04813_),
    .B(_04835_),
    .Y(_04836_));
 sg13g2_a21oi_1 _22674_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[14] ),
    .A2(_04813_),
    .Y(_04837_),
    .B1(_04836_));
 sg13g2_nor2_1 _22675_ (.A(net10991),
    .B(_04837_),
    .Y(_00181_));
 sg13g2_nand2_2 _22676_ (.Y(_04838_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[15] ),
    .B(net10250));
 sg13g2_nor2_1 _22677_ (.A(net9790),
    .B(_04838_),
    .Y(_04839_));
 sg13g2_a21oi_1 _22678_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[15] ),
    .A2(net9790),
    .Y(_04840_),
    .B1(_04839_));
 sg13g2_nor2_1 _22679_ (.A(net10991),
    .B(_04840_),
    .Y(_00182_));
 sg13g2_nand2_2 _22680_ (.Y(_04841_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[16] ),
    .B(net10248));
 sg13g2_nor2_1 _22681_ (.A(_04813_),
    .B(_04841_),
    .Y(_04842_));
 sg13g2_a21oi_1 _22682_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[16] ),
    .A2(_04813_),
    .Y(_04843_),
    .B1(_04842_));
 sg13g2_nor2_1 _22683_ (.A(net10994),
    .B(_04843_),
    .Y(_00183_));
 sg13g2_buf_2 place9961 (.A(net9959),
    .X(net9961));
 sg13g2_nand2_2 _22685_ (.Y(_04845_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[17] ),
    .B(net10248));
 sg13g2_nor2_1 _22686_ (.A(net9780),
    .B(_04845_),
    .Y(_04846_));
 sg13g2_a21oi_1 _22687_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[17] ),
    .A2(net9781),
    .Y(_04847_),
    .B1(_04846_));
 sg13g2_nor2_1 _22688_ (.A(net10994),
    .B(_04847_),
    .Y(_00184_));
 sg13g2_nand2_2 _22689_ (.Y(_04848_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[18] ),
    .B(net10248));
 sg13g2_nor2_1 _22690_ (.A(net9780),
    .B(_04848_),
    .Y(_04849_));
 sg13g2_a21oi_1 _22691_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[18] ),
    .A2(net9780),
    .Y(_04850_),
    .B1(_04849_));
 sg13g2_nor2_1 _22692_ (.A(net10994),
    .B(_04850_),
    .Y(_00185_));
 sg13g2_buf_2 place9956 (.A(net9955),
    .X(net9956));
 sg13g2_nand2_2 _22694_ (.Y(_04852_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[19] ),
    .B(net10248));
 sg13g2_nor2_1 _22695_ (.A(net9780),
    .B(_04852_),
    .Y(_04853_));
 sg13g2_a21oi_1 _22696_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[19] ),
    .A2(net9780),
    .Y(_04854_),
    .B1(_04853_));
 sg13g2_nor2_1 _22697_ (.A(net10994),
    .B(_04854_),
    .Y(_00186_));
 sg13g2_buf_2 place9958 (.A(net9957),
    .X(net9958));
 sg13g2_nand2_2 _22699_ (.Y(_04856_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[1] ),
    .B(net10249));
 sg13g2_nor2_1 _22700_ (.A(net9786),
    .B(_04856_),
    .Y(_04857_));
 sg13g2_a21oi_1 _22701_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[1] ),
    .A2(net9786),
    .Y(_04858_),
    .B1(_04857_));
 sg13g2_nor2_1 _22702_ (.A(net10981),
    .B(_04858_),
    .Y(_00187_));
 sg13g2_nand2_2 _22703_ (.Y(_04859_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[20] ),
    .B(net10251));
 sg13g2_nor2_1 _22704_ (.A(net9781),
    .B(_04859_),
    .Y(_04860_));
 sg13g2_a21oi_1 _22705_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[20] ),
    .A2(net9781),
    .Y(_04861_),
    .B1(_04860_));
 sg13g2_nor2_1 _22706_ (.A(net10993),
    .B(_04861_),
    .Y(_00188_));
 sg13g2_nand2_2 _22707_ (.Y(_04862_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[21] ),
    .B(net10251));
 sg13g2_nor2_1 _22708_ (.A(net9782),
    .B(_04862_),
    .Y(_04863_));
 sg13g2_a21oi_1 _22709_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[21] ),
    .A2(net9782),
    .Y(_04864_),
    .B1(_04863_));
 sg13g2_nor2_1 _22710_ (.A(net10996),
    .B(_04864_),
    .Y(_00189_));
 sg13g2_buf_2 place9960 (.A(net9959),
    .X(net9960));
 sg13g2_nand2_2 _22712_ (.Y(_04866_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[22] ),
    .B(net10251));
 sg13g2_nor2_1 _22713_ (.A(net9781),
    .B(_04866_),
    .Y(_04867_));
 sg13g2_a21oi_1 _22714_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[22] ),
    .A2(net9781),
    .Y(_04868_),
    .B1(_04867_));
 sg13g2_nor2_1 _22715_ (.A(net10996),
    .B(_04868_),
    .Y(_00190_));
 sg13g2_nand2_2 _22716_ (.Y(_04869_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[23] ),
    .B(net10251));
 sg13g2_nor2_1 _22717_ (.A(net9782),
    .B(_04869_),
    .Y(_04870_));
 sg13g2_a21oi_1 _22718_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[23] ),
    .A2(net9782),
    .Y(_04871_),
    .B1(_04870_));
 sg13g2_nor2_1 _22719_ (.A(net10996),
    .B(_04871_),
    .Y(_00191_));
 sg13g2_nand2_2 _22720_ (.Y(_04872_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[24] ),
    .B(net10246));
 sg13g2_nor2_1 _22721_ (.A(net9782),
    .B(_04872_),
    .Y(_04873_));
 sg13g2_a21oi_1 _22722_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[24] ),
    .A2(net9783),
    .Y(_04874_),
    .B1(_04873_));
 sg13g2_nor2_1 _22723_ (.A(net10998),
    .B(_04874_),
    .Y(_00192_));
 sg13g2_nand2_2 _22724_ (.Y(_04875_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[25] ),
    .B(net10246));
 sg13g2_nor2_1 _22725_ (.A(net9783),
    .B(_04875_),
    .Y(_04876_));
 sg13g2_a21oi_1 _22726_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[25] ),
    .A2(net9783),
    .Y(_04877_),
    .B1(_04876_));
 sg13g2_nor2_1 _22727_ (.A(net10998),
    .B(_04877_),
    .Y(_00193_));
 sg13g2_buf_16 clkbuf_leaf_375_clk (.X(clknet_leaf_375_clk),
    .A(clknet_8_120_0_clk));
 sg13g2_nand2_2 _22729_ (.Y(_04879_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[26] ),
    .B(net10251));
 sg13g2_nor2_1 _22730_ (.A(net9783),
    .B(_04879_),
    .Y(_04880_));
 sg13g2_a21oi_1 _22731_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[26] ),
    .A2(net9783),
    .Y(_04881_),
    .B1(_04880_));
 sg13g2_nor2_1 _22732_ (.A(net10998),
    .B(_04881_),
    .Y(_00194_));
 sg13g2_nand2_2 _22733_ (.Y(_04882_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[27] ),
    .B(net10251));
 sg13g2_nor2_1 _22734_ (.A(net9784),
    .B(_04882_),
    .Y(_04883_));
 sg13g2_a21oi_1 _22735_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[27] ),
    .A2(net9785),
    .Y(_04884_),
    .B1(_04883_));
 sg13g2_nor2_1 _22736_ (.A(net10997),
    .B(_04884_),
    .Y(_00195_));
 sg13g2_buf_2 place9951 (.A(net9950),
    .X(net9951));
 sg13g2_nand2_2 _22738_ (.Y(_04886_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[28] ),
    .B(net10251));
 sg13g2_nor2_1 _22739_ (.A(net9784),
    .B(_04886_),
    .Y(_04887_));
 sg13g2_a21oi_1 _22740_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[28] ),
    .A2(net9784),
    .Y(_04888_),
    .B1(_04887_));
 sg13g2_nor2_1 _22741_ (.A(net10997),
    .B(_04888_),
    .Y(_00196_));
 sg13g2_buf_2 place9950 (.A(net9949),
    .X(net9950));
 sg13g2_nand2_2 _22743_ (.Y(_04890_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[29] ),
    .B(net10246));
 sg13g2_nor2_1 _22744_ (.A(net9784),
    .B(_04890_),
    .Y(_04891_));
 sg13g2_a21oi_1 _22745_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[29] ),
    .A2(net9784),
    .Y(_04892_),
    .B1(_04891_));
 sg13g2_nor2_1 _22746_ (.A(net11000),
    .B(_04892_),
    .Y(_00197_));
 sg13g2_nand2_2 _22747_ (.Y(_04893_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[2] ),
    .B(net10249));
 sg13g2_nor2_1 _22748_ (.A(net9786),
    .B(_04893_),
    .Y(_04894_));
 sg13g2_a21oi_1 _22749_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[2] ),
    .A2(net9786),
    .Y(_04895_),
    .B1(_04894_));
 sg13g2_nor2_1 _22750_ (.A(net10981),
    .B(_04895_),
    .Y(_00198_));
 sg13g2_nand2_2 _22751_ (.Y(_04896_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[30] ),
    .B(net10246));
 sg13g2_nor2_1 _22752_ (.A(net9785),
    .B(_04896_),
    .Y(_04897_));
 sg13g2_a21oi_1 _22753_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[30] ),
    .A2(net9785),
    .Y(_04898_),
    .B1(_04897_));
 sg13g2_nor2_1 _22754_ (.A(net11000),
    .B(_04898_),
    .Y(_00199_));
 sg13g2_buf_2 place10023 (.A(_11043_),
    .X(net10023));
 sg13g2_buf_2 place9947 (.A(net9945),
    .X(net9947));
 sg13g2_nand2_2 _22757_ (.Y(_04901_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[31] ),
    .B(net10251));
 sg13g2_nor2_1 _22758_ (.A(net9785),
    .B(_04901_),
    .Y(_04902_));
 sg13g2_a21oi_1 _22759_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[31] ),
    .A2(net9785),
    .Y(_04903_),
    .B1(_04902_));
 sg13g2_nor2_1 _22760_ (.A(net11000),
    .B(_04903_),
    .Y(_00200_));
 sg13g2_nand2_2 _22761_ (.Y(_04904_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[3] ),
    .B(net10249));
 sg13g2_nor2_1 _22762_ (.A(net9786),
    .B(_04904_),
    .Y(_04905_));
 sg13g2_a21oi_1 _22763_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[3] ),
    .A2(net9787),
    .Y(_04906_),
    .B1(_04905_));
 sg13g2_nor2_1 _22764_ (.A(net10981),
    .B(_04906_),
    .Y(_00201_));
 sg13g2_nand2_2 _22765_ (.Y(_04907_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[4] ),
    .B(net10249));
 sg13g2_nor2_1 _22766_ (.A(net9787),
    .B(_04907_),
    .Y(_04908_));
 sg13g2_a21oi_1 _22767_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[4] ),
    .A2(net9787),
    .Y(_04909_),
    .B1(_04908_));
 sg13g2_nor2_1 _22768_ (.A(net10984),
    .B(_04909_),
    .Y(_00202_));
 sg13g2_nand2_2 _22769_ (.Y(_04910_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[5] ),
    .B(net10249));
 sg13g2_nor2_1 _22770_ (.A(net9789),
    .B(_04910_),
    .Y(_04911_));
 sg13g2_a21oi_1 _22771_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[5] ),
    .A2(net9787),
    .Y(_04912_),
    .B1(_04911_));
 sg13g2_nor2_1 _22772_ (.A(net10984),
    .B(_04912_),
    .Y(_00203_));
 sg13g2_nand2_2 _22773_ (.Y(_04913_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[6] ),
    .B(net10249));
 sg13g2_nor2_1 _22774_ (.A(net9789),
    .B(_04913_),
    .Y(_04914_));
 sg13g2_a21oi_1 _22775_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[6] ),
    .A2(net9789),
    .Y(_04915_),
    .B1(_04914_));
 sg13g2_nor2_1 _22776_ (.A(net10984),
    .B(_04915_),
    .Y(_00204_));
 sg13g2_nand2_2 _22777_ (.Y(_04916_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[7] ),
    .B(net10250));
 sg13g2_nor2_1 _22778_ (.A(net9789),
    .B(_04916_),
    .Y(_04917_));
 sg13g2_a21oi_1 _22779_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[7] ),
    .A2(net9789),
    .Y(_04918_),
    .B1(_04917_));
 sg13g2_nor2_1 _22780_ (.A(net10984),
    .B(_04918_),
    .Y(_00205_));
 sg13g2_nand2_2 _22781_ (.Y(_04919_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[8] ),
    .B(net10250));
 sg13g2_nor2_1 _22782_ (.A(net9789),
    .B(_04919_),
    .Y(_04920_));
 sg13g2_a21oi_1 _22783_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[8] ),
    .A2(net9789),
    .Y(_04921_),
    .B1(_04920_));
 sg13g2_nor2_1 _22784_ (.A(net10984),
    .B(_04921_),
    .Y(_00206_));
 sg13g2_nand2_2 _22785_ (.Y(_04922_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[9] ),
    .B(net10250));
 sg13g2_nor2_1 _22786_ (.A(net9789),
    .B(_04922_),
    .Y(_04923_));
 sg13g2_a21oi_1 _22787_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[9] ),
    .A2(net9788),
    .Y(_04924_),
    .B1(_04923_));
 sg13g2_nor2_1 _22788_ (.A(net10985),
    .B(_04924_),
    .Y(_00207_));
 sg13g2_and2_1 _22789_ (.A(resetn),
    .B(gpio_in1),
    .X(_00208_));
 sg13g2_and2_1 _22790_ (.A(resetn),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in1_sync1 ),
    .X(_00209_));
 sg13g2_buf_2 place9946 (.A(net9945),
    .X(net9946));
 sg13g2_and2_1 _22792_ (.A(resetn),
    .B(gpio_in2),
    .X(_00210_));
 sg13g2_and2_1 _22793_ (.A(resetn),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in2_sync1 ),
    .X(_00211_));
 sg13g2_nor3_2 _22794_ (.A(net10615),
    .B(net10617),
    .C(_04807_),
    .Y(_04926_));
 sg13g2_buf_2 place9953 (.A(net9949),
    .X(net9953));
 sg13g2_nand3_1 _22796_ (.B(_04803_),
    .C(_04926_),
    .A(net10620),
    .Y(_04928_));
 sg13g2_o21ai_1 _22797_ (.B1(_04928_),
    .Y(_04929_),
    .A1(gpio_io1_oe),
    .A2(_04926_));
 sg13g2_nor2_1 _22798_ (.A(_04803_),
    .B(_04809_),
    .Y(_04930_));
 sg13g2_nand3b_1 _22799_ (.B(_04930_),
    .C(net10620),
    .Y(_04931_),
    .A_N(\u_ac_controller_soc_inst.cbus_wdata[0] ));
 sg13g2_o21ai_1 _22800_ (.B1(_04931_),
    .Y(_04932_),
    .A1(gpio_io1_oe),
    .A2(_04930_));
 sg13g2_mux2_1 _22801_ (.A0(_04929_),
    .A1(_04932_),
    .S(_08126_),
    .X(_04933_));
 sg13g2_nor2_2 _22802_ (.A(net10987),
    .B(net10186),
    .Y(_00248_));
 sg13g2_o21ai_1 _22803_ (.B1(_00248_),
    .Y(_04934_),
    .A1(net10620),
    .A2(gpio_io1_oe));
 sg13g2_nor2_1 _22804_ (.A(_04933_),
    .B(_04934_),
    .Y(_00212_));
 sg13g2_nand2_1 _22805_ (.Y(_04935_),
    .A(_08126_),
    .B(net10459));
 sg13g2_a21oi_2 _22806_ (.B1(_04809_),
    .Y(_04936_),
    .A2(net10247),
    .A1(_04935_));
 sg13g2_nand2_1 _22807_ (.Y(_04937_),
    .A(_04803_),
    .B(_04936_));
 sg13g2_or2_1 _22808_ (.X(_04938_),
    .B(_04936_),
    .A(gpio_io2_oe));
 sg13g2_nand3_1 _22809_ (.B(net10459),
    .C(_04930_),
    .A(net10618),
    .Y(_04939_));
 sg13g2_mux2_1 _22810_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[0] ),
    .A1(_04938_),
    .S(_04939_),
    .X(_04940_));
 sg13g2_and3_1 _22811_ (.X(_00213_),
    .A(_00248_),
    .B(_04937_),
    .C(_04940_));
 sg13g2_nand4_1 _22812_ (.B(net10620),
    .C(_04804_),
    .A(net10618),
    .Y(_04941_),
    .D(_04926_));
 sg13g2_nand2_1 _22813_ (.Y(_04942_),
    .A(gpio_out1),
    .B(_04941_));
 sg13g2_or2_1 _22814_ (.X(_04943_),
    .B(_04941_),
    .A(_04817_));
 sg13g2_buf_2 place10217 (.A(_11408_),
    .X(net10217));
 sg13g2_a21oi_1 _22816_ (.A1(_04942_),
    .A2(_04943_),
    .Y(_00214_),
    .B1(net11035));
 sg13g2_nand2_2 _22817_ (.Y(_04945_),
    .A(_04804_),
    .B(_04936_));
 sg13g2_nand2_1 _22818_ (.Y(_04946_),
    .A(gpio_out2),
    .B(_04945_));
 sg13g2_o21ai_1 _22819_ (.B1(_04946_),
    .Y(_04947_),
    .A1(_04817_),
    .A2(_04945_));
 sg13g2_and2_1 _22820_ (.A(resetn),
    .B(_04947_),
    .X(_00215_));
 sg13g2_nand2_1 _22821_ (.Y(_04948_),
    .A(net10459),
    .B(_07707_));
 sg13g2_nand3_1 _22822_ (.B(net10617),
    .C(net10247),
    .A(net10620),
    .Y(_04949_));
 sg13g2_a21oi_1 _22823_ (.A1(_04948_),
    .A2(_04949_),
    .Y(_04950_),
    .B1(net10618));
 sg13g2_and4_1 _22824_ (.A(net10618),
    .B(net10459),
    .C(net10617),
    .D(net10247),
    .X(_04951_));
 sg13g2_nor4_1 _22825_ (.A(net10615),
    .B(_04807_),
    .C(_04950_),
    .D(_04951_),
    .Y(_04952_));
 sg13g2_nor4_2 _22826_ (.A(net10615),
    .B(net10617),
    .C(_04935_),
    .Y(_04953_),
    .D(_04807_));
 sg13g2_nor2_1 _22827_ (.A(net10186),
    .B(_04802_),
    .Y(_04954_));
 sg13g2_o21ai_1 _22828_ (.B1(_04954_),
    .Y(_04955_),
    .A1(_04952_),
    .A2(_04953_));
 sg13g2_buf_2 place9945 (.A(_10293_),
    .X(net9945));
 sg13g2_buf_2 place9949 (.A(_10293_),
    .X(net9949));
 sg13g2_buf_2 place9948 (.A(net9947),
    .X(net9948));
 sg13g2_nand2b_1 _22832_ (.Y(_04959_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_enable ),
    .A_N(_04952_));
 sg13g2_buf_2 place9940 (.A(_10375_),
    .X(net9940));
 sg13g2_mux2_1 _22834_ (.A0(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[0] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in1_sync ),
    .S(net10620),
    .X(_04961_));
 sg13g2_a22oi_1 _22835_ (.Y(_04962_),
    .B1(_04961_),
    .B2(net10618),
    .A2(_04562_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[0] ));
 sg13g2_nor2b_1 _22836_ (.A(_04962_),
    .B_N(_04926_),
    .Y(_04963_));
 sg13g2_a221oi_1 _22837_ (.B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in2_sync ),
    .C1(_04963_),
    .B1(_04936_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[0] ),
    .Y(_04964_),
    .A2(_04811_));
 sg13g2_buf_2 place9939 (.A(net9936),
    .X(net9939));
 sg13g2_a21oi_1 _22839_ (.A1(_04959_),
    .A2(_04964_),
    .Y(_04966_),
    .B1(_04955_));
 sg13g2_a21oi_1 _22840_ (.A1(\u_ac_controller_soc_inst.io_rdata[0] ),
    .A2(_04955_),
    .Y(_04967_),
    .B1(_04966_));
 sg13g2_nor2_1 _22841_ (.A(net10987),
    .B(_04967_),
    .Y(_00216_));
 sg13g2_buf_2 place10033 (.A(net10032),
    .X(net10033));
 sg13g2_nand2_1 _22843_ (.Y(_04969_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[10] ),
    .B(net9824));
 sg13g2_buf_2 place9944 (.A(net9942),
    .X(net9944));
 sg13g2_and3_2 _22845_ (.X(_04971_),
    .A(net10618),
    .B(net10459),
    .C(_04926_));
 sg13g2_buf_2 place9952 (.A(net9951),
    .X(net9952));
 sg13g2_buf_2 place9964 (.A(net9962),
    .X(net9964));
 sg13g2_and2_1 _22848_ (.A(_04562_),
    .B(_04926_),
    .X(_04974_));
 sg13g2_buf_2 place9942 (.A(_10375_),
    .X(net9942));
 sg13g2_buf_2 place9954 (.A(net9953),
    .X(net9954));
 sg13g2_a22oi_1 _22851_ (.Y(_04977_),
    .B1(net9815),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[10] ),
    .A2(net9817),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[10] ));
 sg13g2_a21oi_2 _22852_ (.B1(net9771),
    .Y(_04978_),
    .A2(_04977_),
    .A1(_04969_));
 sg13g2_a21oi_1 _22853_ (.A1(\u_ac_controller_soc_inst.io_rdata[10] ),
    .A2(net9772),
    .Y(_04979_),
    .B1(_04978_));
 sg13g2_nor2_1 _22854_ (.A(net10990),
    .B(_04979_),
    .Y(_00217_));
 sg13g2_buf_2 place9943 (.A(net9942),
    .X(net9943));
 sg13g2_nand2_1 _22856_ (.Y(_04981_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[11] ),
    .B(net9825));
 sg13g2_buf_2 place9941 (.A(_10375_),
    .X(net9941));
 sg13g2_a22oi_1 _22858_ (.Y(_04983_),
    .B1(net9815),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[11] ),
    .A2(net9817),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[11] ));
 sg13g2_a21oi_2 _22859_ (.B1(net9774),
    .Y(_04984_),
    .A2(_04983_),
    .A1(_04981_));
 sg13g2_a21oi_1 _22860_ (.A1(\u_ac_controller_soc_inst.io_rdata[11] ),
    .A2(net9775),
    .Y(_04985_),
    .B1(_04984_));
 sg13g2_nor2_1 _22861_ (.A(net10993),
    .B(_04985_),
    .Y(_00218_));
 sg13g2_nand2_1 _22862_ (.Y(_04986_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[12] ),
    .B(net9825));
 sg13g2_buf_16 clkbuf_leaf_376_clk (.X(clknet_leaf_376_clk),
    .A(clknet_8_108_0_clk));
 sg13g2_a22oi_1 _22864_ (.Y(_04988_),
    .B1(net9815),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[12] ),
    .A2(net9817),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[12] ));
 sg13g2_a21oi_1 _22865_ (.A1(_04986_),
    .A2(_04988_),
    .Y(_04989_),
    .B1(net9774));
 sg13g2_a21oi_1 _22866_ (.A1(\u_ac_controller_soc_inst.io_rdata[12] ),
    .A2(net9773),
    .Y(_04990_),
    .B1(_04989_));
 sg13g2_nor2_1 _22867_ (.A(net10990),
    .B(_04990_),
    .Y(_00219_));
 sg13g2_nand2_1 _22868_ (.Y(_04991_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[13] ),
    .B(net9825));
 sg13g2_buf_2 place9927 (.A(net9926),
    .X(net9927));
 sg13g2_a22oi_1 _22870_ (.Y(_04993_),
    .B1(net9815),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[13] ),
    .A2(net9817),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[13] ));
 sg13g2_a21oi_1 _22871_ (.A1(_04991_),
    .A2(_04993_),
    .Y(_04994_),
    .B1(net9774));
 sg13g2_a21oi_1 _22872_ (.A1(\u_ac_controller_soc_inst.io_rdata[13] ),
    .A2(net9775),
    .Y(_04995_),
    .B1(_04994_));
 sg13g2_nor2_1 _22873_ (.A(net10993),
    .B(_04995_),
    .Y(_00220_));
 sg13g2_nand2_1 _22874_ (.Y(_04996_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[14] ),
    .B(_04811_));
 sg13g2_buf_2 place9926 (.A(_10455_),
    .X(net9926));
 sg13g2_a22oi_1 _22876_ (.Y(_04998_),
    .B1(net9812),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[14] ),
    .A2(net9818),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[14] ));
 sg13g2_a21oi_2 _22877_ (.B1(net9773),
    .Y(_04999_),
    .A2(_04998_),
    .A1(_04996_));
 sg13g2_a21oi_1 _22878_ (.A1(\u_ac_controller_soc_inst.io_rdata[14] ),
    .A2(net9776),
    .Y(_05000_),
    .B1(_04999_));
 sg13g2_nor2_1 _22879_ (.A(net10996),
    .B(_05000_),
    .Y(_00221_));
 sg13g2_nand2_1 _22880_ (.Y(_05001_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[15] ),
    .B(net9825));
 sg13g2_buf_2 place9938 (.A(net9937),
    .X(net9938));
 sg13g2_a22oi_1 _22882_ (.Y(_05003_),
    .B1(net9812),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[15] ),
    .A2(net9817),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[15] ));
 sg13g2_a21oi_1 _22883_ (.A1(_05001_),
    .A2(_05003_),
    .Y(_05004_),
    .B1(net9774));
 sg13g2_a21oi_1 _22884_ (.A1(\u_ac_controller_soc_inst.io_rdata[15] ),
    .A2(net9773),
    .Y(_05005_),
    .B1(_05004_));
 sg13g2_nor2_1 _22885_ (.A(net10993),
    .B(_05005_),
    .Y(_00222_));
 sg13g2_nand2_1 _22886_ (.Y(_05006_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[16] ),
    .B(_04811_));
 sg13g2_buf_2 place9933 (.A(net9931),
    .X(net9933));
 sg13g2_a22oi_1 _22888_ (.Y(_05008_),
    .B1(net9812),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[16] ),
    .A2(net9818),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[16] ));
 sg13g2_a21oi_1 _22889_ (.A1(_05006_),
    .A2(_05008_),
    .Y(_05009_),
    .B1(net9775));
 sg13g2_a21oi_1 _22890_ (.A1(\u_ac_controller_soc_inst.io_rdata[16] ),
    .A2(net9776),
    .Y(_05010_),
    .B1(_05009_));
 sg13g2_nor2_1 _22891_ (.A(net10993),
    .B(_05010_),
    .Y(_00223_));
 sg13g2_nand2_1 _22892_ (.Y(_05011_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[17] ),
    .B(net9821));
 sg13g2_buf_2 place9929 (.A(net9926),
    .X(net9929));
 sg13g2_a22oi_1 _22894_ (.Y(_05013_),
    .B1(net9813),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[17] ),
    .A2(net9818),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[17] ));
 sg13g2_buf_2 place9932 (.A(net9931),
    .X(net9932));
 sg13g2_a21oi_1 _22896_ (.A1(_05011_),
    .A2(_05013_),
    .Y(_05015_),
    .B1(net9775));
 sg13g2_a21oi_1 _22897_ (.A1(\u_ac_controller_soc_inst.io_rdata[17] ),
    .A2(net9776),
    .Y(_05016_),
    .B1(_05015_));
 sg13g2_nor2_1 _22898_ (.A(net10997),
    .B(_05016_),
    .Y(_00224_));
 sg13g2_nand2_1 _22899_ (.Y(_05017_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[18] ),
    .B(net9821));
 sg13g2_buf_2 place9928 (.A(net9927),
    .X(net9928));
 sg13g2_a22oi_1 _22901_ (.Y(_05019_),
    .B1(net9813),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[18] ),
    .A2(net9818),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[18] ));
 sg13g2_a21oi_2 _22902_ (.B1(net9775),
    .Y(_05020_),
    .A2(_05019_),
    .A1(_05017_));
 sg13g2_a21oi_1 _22903_ (.A1(\u_ac_controller_soc_inst.io_rdata[18] ),
    .A2(net9779),
    .Y(_05021_),
    .B1(_05020_));
 sg13g2_nor2_1 _22904_ (.A(net11001),
    .B(_05021_),
    .Y(_00225_));
 sg13g2_buf_2 place9930 (.A(_10455_),
    .X(net9930));
 sg13g2_nand2_1 _22906_ (.Y(_05023_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[19] ),
    .B(net9821));
 sg13g2_buf_2 place9931 (.A(net9930),
    .X(net9931));
 sg13g2_a22oi_1 _22908_ (.Y(_05025_),
    .B1(net9813),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[19] ),
    .A2(net9818),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[19] ));
 sg13g2_a21oi_2 _22909_ (.B1(net9775),
    .Y(_05026_),
    .A2(_05025_),
    .A1(_05023_));
 sg13g2_a21oi_1 _22910_ (.A1(\u_ac_controller_soc_inst.io_rdata[19] ),
    .A2(net9779),
    .Y(_05027_),
    .B1(_05026_));
 sg13g2_nor2_1 _22911_ (.A(net11001),
    .B(_05027_),
    .Y(_00226_));
 sg13g2_buf_16 clkbuf_leaf_377_clk (.X(clknet_leaf_377_clk),
    .A(clknet_8_109_0_clk));
 sg13g2_nand2_1 _22913_ (.Y(_05029_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[1] ),
    .B(net9823));
 sg13g2_buf_2 place9924 (.A(net9923),
    .X(net9924));
 sg13g2_buf_2 place9918 (.A(net9917),
    .X(net9918));
 sg13g2_buf_2 place9922 (.A(_10496_),
    .X(net9922));
 sg13g2_a22oi_1 _22917_ (.Y(_05033_),
    .B1(net9812),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[1] ),
    .A2(net9816),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[1] ));
 sg13g2_a21oi_1 _22918_ (.A1(_05029_),
    .A2(_05033_),
    .Y(_05034_),
    .B1(_04955_));
 sg13g2_a21oi_1 _22919_ (.A1(\u_ac_controller_soc_inst.io_rdata[1] ),
    .A2(net9772),
    .Y(_05035_),
    .B1(_05034_));
 sg13g2_nor2_1 _22920_ (.A(net10989),
    .B(_05035_),
    .Y(_00227_));
 sg13g2_buf_2 place9921 (.A(_10496_),
    .X(net9921));
 sg13g2_nand2_1 _22922_ (.Y(_05037_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[20] ),
    .B(net9821));
 sg13g2_buf_2 place9937 (.A(net9936),
    .X(net9937));
 sg13g2_a22oi_1 _22924_ (.Y(_05039_),
    .B1(net9813),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[20] ),
    .A2(net9819),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[20] ));
 sg13g2_a21oi_1 _22925_ (.A1(_05037_),
    .A2(_05039_),
    .Y(_05040_),
    .B1(net9775));
 sg13g2_a21oi_1 _22926_ (.A1(\u_ac_controller_soc_inst.io_rdata[20] ),
    .A2(net9776),
    .Y(_05041_),
    .B1(_05040_));
 sg13g2_nor2_1 _22927_ (.A(net10996),
    .B(_05041_),
    .Y(_00228_));
 sg13g2_nand2_1 _22928_ (.Y(_05042_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[21] ),
    .B(net9821));
 sg13g2_buf_2 place9917 (.A(net9916),
    .X(net9917));
 sg13g2_a22oi_1 _22930_ (.Y(_05044_),
    .B1(net9813),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[21] ),
    .A2(net9819),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[21] ));
 sg13g2_a21oi_1 _22931_ (.A1(_05042_),
    .A2(_05044_),
    .Y(_05045_),
    .B1(net9776));
 sg13g2_a21oi_1 _22932_ (.A1(\u_ac_controller_soc_inst.io_rdata[21] ),
    .A2(net9776),
    .Y(_05046_),
    .B1(_05045_));
 sg13g2_nor2_1 _22933_ (.A(net10996),
    .B(_05046_),
    .Y(_00229_));
 sg13g2_nand2_1 _22934_ (.Y(_05047_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[22] ),
    .B(net9821));
 sg13g2_buf_2 place9916 (.A(_10496_),
    .X(net9916));
 sg13g2_a22oi_1 _22936_ (.Y(_05049_),
    .B1(net9813),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[22] ),
    .A2(net9819),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[22] ));
 sg13g2_a21oi_1 _22937_ (.A1(_05047_),
    .A2(_05049_),
    .Y(_05050_),
    .B1(net9776));
 sg13g2_a21oi_1 _22938_ (.A1(\u_ac_controller_soc_inst.io_rdata[22] ),
    .A2(net9777),
    .Y(_05051_),
    .B1(_05050_));
 sg13g2_nor2_1 _22939_ (.A(net10996),
    .B(_05051_),
    .Y(_00230_));
 sg13g2_nand2_1 _22940_ (.Y(_05052_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[23] ),
    .B(net9821));
 sg13g2_buf_2 place9923 (.A(net9922),
    .X(net9923));
 sg13g2_a22oi_1 _22942_ (.Y(_05054_),
    .B1(net9813),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[23] ),
    .A2(net9819),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[23] ));
 sg13g2_a21oi_1 _22943_ (.A1(_05052_),
    .A2(_05054_),
    .Y(_05055_),
    .B1(net9776));
 sg13g2_a21oi_1 _22944_ (.A1(\u_ac_controller_soc_inst.io_rdata[23] ),
    .A2(net9777),
    .Y(_05056_),
    .B1(_05055_));
 sg13g2_nor2_1 _22945_ (.A(net10997),
    .B(_05056_),
    .Y(_00231_));
 sg13g2_nand2_1 _22946_ (.Y(_05057_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[24] ),
    .B(net9822));
 sg13g2_a22oi_1 _22947_ (.Y(_05058_),
    .B1(net9814),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[24] ),
    .A2(net9820),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[24] ));
 sg13g2_a21oi_1 _22948_ (.A1(_05057_),
    .A2(_05058_),
    .Y(_05059_),
    .B1(net9777));
 sg13g2_a21oi_1 _22949_ (.A1(\u_ac_controller_soc_inst.io_rdata[24] ),
    .A2(net9778),
    .Y(_05060_),
    .B1(_05059_));
 sg13g2_nor2_1 _22950_ (.A(net10997),
    .B(_05060_),
    .Y(_00232_));
 sg13g2_nand2_1 _22951_ (.Y(_05061_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[25] ),
    .B(net9822));
 sg13g2_buf_2 place9919 (.A(net9917),
    .X(net9919));
 sg13g2_a22oi_1 _22953_ (.Y(_05063_),
    .B1(net9814),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[25] ),
    .A2(net9820),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[25] ));
 sg13g2_a21oi_1 _22954_ (.A1(_05061_),
    .A2(_05063_),
    .Y(_05064_),
    .B1(net9777));
 sg13g2_a21oi_1 _22955_ (.A1(\u_ac_controller_soc_inst.io_rdata[25] ),
    .A2(net9778),
    .Y(_05065_),
    .B1(_05064_));
 sg13g2_nor2_1 _22956_ (.A(net10997),
    .B(_05065_),
    .Y(_00233_));
 sg13g2_nand2_1 _22957_ (.Y(_05066_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[26] ),
    .B(net9822));
 sg13g2_buf_2 place9913 (.A(net9912),
    .X(net9913));
 sg13g2_a22oi_1 _22959_ (.Y(_05068_),
    .B1(net9814),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[26] ),
    .A2(net9820),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[26] ));
 sg13g2_buf_2 place9907 (.A(_10608_),
    .X(net9907));
 sg13g2_a21oi_1 _22961_ (.A1(_05066_),
    .A2(_05068_),
    .Y(_05070_),
    .B1(net9777));
 sg13g2_a21oi_1 _22962_ (.A1(\u_ac_controller_soc_inst.io_rdata[26] ),
    .A2(net9779),
    .Y(_05071_),
    .B1(_05070_));
 sg13g2_nor2_1 _22963_ (.A(net11001),
    .B(_05071_),
    .Y(_00234_));
 sg13g2_nand2_1 _22964_ (.Y(_05072_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[27] ),
    .B(net9822));
 sg13g2_buf_2 place10888 (.A(net10885),
    .X(net10888));
 sg13g2_a22oi_1 _22966_ (.Y(_05074_),
    .B1(net9814),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[27] ),
    .A2(net9820),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[27] ));
 sg13g2_a21oi_1 _22967_ (.A1(_05072_),
    .A2(_05074_),
    .Y(_05075_),
    .B1(net9778));
 sg13g2_a21oi_1 _22968_ (.A1(\u_ac_controller_soc_inst.io_rdata[27] ),
    .A2(net9779),
    .Y(_05076_),
    .B1(_05075_));
 sg13g2_nor2_1 _22969_ (.A(net11001),
    .B(_05076_),
    .Y(_00235_));
 sg13g2_buf_2 place9915 (.A(net9914),
    .X(net9915));
 sg13g2_nand2_1 _22971_ (.Y(_05078_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[28] ),
    .B(net9822));
 sg13g2_buf_2 place9911 (.A(_10608_),
    .X(net9911));
 sg13g2_a22oi_1 _22973_ (.Y(_05080_),
    .B1(net9814),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[28] ),
    .A2(net9820),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[28] ));
 sg13g2_a21oi_1 _22974_ (.A1(_05078_),
    .A2(_05080_),
    .Y(_05081_),
    .B1(net9778));
 sg13g2_a21oi_1 _22975_ (.A1(\u_ac_controller_soc_inst.io_rdata[28] ),
    .A2(net9778),
    .Y(_05082_),
    .B1(_05081_));
 sg13g2_nor2_1 _22976_ (.A(net11001),
    .B(_05082_),
    .Y(_00236_));
 sg13g2_buf_2 place9909 (.A(_10608_),
    .X(net9909));
 sg13g2_nand2_1 _22978_ (.Y(_05084_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[29] ),
    .B(net9822));
 sg13g2_buf_2 place9912 (.A(net9911),
    .X(net9912));
 sg13g2_buf_2 place9914 (.A(_10608_),
    .X(net9914));
 sg13g2_buf_2 place9908 (.A(net9907),
    .X(net9908));
 sg13g2_a22oi_1 _22982_ (.Y(_05088_),
    .B1(net9814),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[29] ),
    .A2(net9820),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[29] ));
 sg13g2_a21oi_1 _22983_ (.A1(_05084_),
    .A2(_05088_),
    .Y(_05089_),
    .B1(net9778));
 sg13g2_a21oi_1 _22984_ (.A1(\u_ac_controller_soc_inst.io_rdata[29] ),
    .A2(net9778),
    .Y(_05090_),
    .B1(_05089_));
 sg13g2_nor2_1 _22985_ (.A(net11001),
    .B(_05090_),
    .Y(_00237_));
 sg13g2_buf_2 place9910 (.A(net9909),
    .X(net9910));
 sg13g2_nand2_1 _22987_ (.Y(_05092_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[2] ),
    .B(net9823));
 sg13g2_buf_2 place9906 (.A(net9905),
    .X(net9906));
 sg13g2_a22oi_1 _22989_ (.Y(_05094_),
    .B1(net9812),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[2] ),
    .A2(net9816),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[2] ));
 sg13g2_a21oi_1 _22990_ (.A1(_05092_),
    .A2(_05094_),
    .Y(_05095_),
    .B1(_04955_));
 sg13g2_a21oi_1 _22991_ (.A1(\u_ac_controller_soc_inst.io_rdata[2] ),
    .A2(_04955_),
    .Y(_05096_),
    .B1(_05095_));
 sg13g2_nor2_1 _22992_ (.A(net10989),
    .B(_05096_),
    .Y(_00238_));
 sg13g2_nand2_1 _22993_ (.Y(_05097_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[30] ),
    .B(net9822));
 sg13g2_buf_2 place9920 (.A(net9919),
    .X(net9920));
 sg13g2_a22oi_1 _22995_ (.Y(_05099_),
    .B1(net9814),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[30] ),
    .A2(net9820),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[30] ));
 sg13g2_a21oi_1 _22996_ (.A1(_05097_),
    .A2(_05099_),
    .Y(_05100_),
    .B1(net9779));
 sg13g2_a21oi_1 _22997_ (.A1(\u_ac_controller_soc_inst.io_rdata[30] ),
    .A2(net9779),
    .Y(_05101_),
    .B1(_05100_));
 sg13g2_nor2_1 _22998_ (.A(net11001),
    .B(_05101_),
    .Y(_00239_));
 sg13g2_nand2_1 _22999_ (.Y(_05102_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[31] ),
    .B(net9822));
 sg13g2_buf_2 place9903 (.A(net9902),
    .X(net9903));
 sg13g2_a22oi_1 _23001_ (.Y(_05104_),
    .B1(net9814),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[31] ),
    .A2(net9820),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[31] ));
 sg13g2_a21oi_1 _23002_ (.A1(_05102_),
    .A2(_05104_),
    .Y(_05105_),
    .B1(net9779));
 sg13g2_a21oi_1 _23003_ (.A1(\u_ac_controller_soc_inst.io_rdata[31] ),
    .A2(net9779),
    .Y(_05106_),
    .B1(_05105_));
 sg13g2_nor2_1 _23004_ (.A(net11001),
    .B(_05106_),
    .Y(_00240_));
 sg13g2_nand2_1 _23005_ (.Y(_05107_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[3] ),
    .B(net9823));
 sg13g2_buf_2 place9901 (.A(net9898),
    .X(net9901));
 sg13g2_a22oi_1 _23007_ (.Y(_05109_),
    .B1(_04974_),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[3] ),
    .A2(net9816),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[3] ));
 sg13g2_a21oi_1 _23008_ (.A1(_05107_),
    .A2(_05109_),
    .Y(_05110_),
    .B1(net9771));
 sg13g2_a21oi_1 _23009_ (.A1(\u_ac_controller_soc_inst.io_rdata[3] ),
    .A2(net9772),
    .Y(_05111_),
    .B1(_05110_));
 sg13g2_nor2_1 _23010_ (.A(net10989),
    .B(_05111_),
    .Y(_00241_));
 sg13g2_nand2_1 _23011_ (.Y(_05112_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[4] ),
    .B(net9823));
 sg13g2_buf_2 place9905 (.A(net9904),
    .X(net9905));
 sg13g2_a22oi_1 _23013_ (.Y(_05114_),
    .B1(_04974_),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[4] ),
    .A2(net9816),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[4] ));
 sg13g2_a21oi_1 _23014_ (.A1(_05112_),
    .A2(_05114_),
    .Y(_05115_),
    .B1(net9771));
 sg13g2_a21oi_1 _23015_ (.A1(\u_ac_controller_soc_inst.io_rdata[4] ),
    .A2(net9772),
    .Y(_05116_),
    .B1(_05115_));
 sg13g2_nor2_1 _23016_ (.A(net10990),
    .B(_05116_),
    .Y(_00242_));
 sg13g2_nand2_1 _23017_ (.Y(_05117_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[5] ),
    .B(net9824));
 sg13g2_buf_2 place9900 (.A(net9898),
    .X(net9900));
 sg13g2_a22oi_1 _23019_ (.Y(_05119_),
    .B1(_04974_),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[5] ),
    .A2(net9816),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[5] ));
 sg13g2_a21oi_1 _23020_ (.A1(_05117_),
    .A2(_05119_),
    .Y(_05120_),
    .B1(net9771));
 sg13g2_a21oi_1 _23021_ (.A1(\u_ac_controller_soc_inst.io_rdata[5] ),
    .A2(net9774),
    .Y(_05121_),
    .B1(_05120_));
 sg13g2_nor2_1 _23022_ (.A(net11002),
    .B(_05121_),
    .Y(_00243_));
 sg13g2_nand2_1 _23023_ (.Y(_05122_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[6] ),
    .B(net9824));
 sg13g2_buf_2 place9898 (.A(_10688_),
    .X(net9898));
 sg13g2_a22oi_1 _23025_ (.Y(_05124_),
    .B1(net9815),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[6] ),
    .A2(net9816),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[6] ));
 sg13g2_a21oi_2 _23026_ (.B1(net9771),
    .Y(_05125_),
    .A2(_05124_),
    .A1(_05122_));
 sg13g2_a21oi_1 _23027_ (.A1(\u_ac_controller_soc_inst.io_rdata[6] ),
    .A2(net9773),
    .Y(_05126_),
    .B1(_05125_));
 sg13g2_nor2_1 _23028_ (.A(net10990),
    .B(_05126_),
    .Y(_00244_));
 sg13g2_nand2_1 _23029_ (.Y(_05127_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[7] ),
    .B(net9824));
 sg13g2_buf_2 place9899 (.A(net9898),
    .X(net9899));
 sg13g2_a22oi_1 _23031_ (.Y(_05129_),
    .B1(net9815),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[7] ),
    .A2(net9817),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[7] ));
 sg13g2_a21oi_2 _23032_ (.B1(net9771),
    .Y(_05130_),
    .A2(_05129_),
    .A1(_05127_));
 sg13g2_a21oi_1 _23033_ (.A1(\u_ac_controller_soc_inst.io_rdata[7] ),
    .A2(_04955_),
    .Y(_05131_),
    .B1(_05130_));
 sg13g2_nor2_1 _23034_ (.A(net10989),
    .B(_05131_),
    .Y(_00245_));
 sg13g2_nand2_1 _23035_ (.Y(_05132_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[8] ),
    .B(net9824));
 sg13g2_buf_2 place9902 (.A(_10688_),
    .X(net9902));
 sg13g2_a22oi_1 _23037_ (.Y(_05134_),
    .B1(net9815),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[8] ),
    .A2(net9817),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[8] ));
 sg13g2_a21oi_2 _23038_ (.B1(net9771),
    .Y(_05135_),
    .A2(_05134_),
    .A1(_05132_));
 sg13g2_a21oi_1 _23039_ (.A1(\u_ac_controller_soc_inst.io_rdata[8] ),
    .A2(net9773),
    .Y(_05136_),
    .B1(_05135_));
 sg13g2_nor2_1 _23040_ (.A(net10990),
    .B(_05136_),
    .Y(_00246_));
 sg13g2_nand2_1 _23041_ (.Y(_05137_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[9] ),
    .B(net9825));
 sg13g2_buf_2 place9904 (.A(_10688_),
    .X(net9904));
 sg13g2_a22oi_1 _23043_ (.Y(_05139_),
    .B1(net9815),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[9] ),
    .A2(net9817),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[9] ));
 sg13g2_a21oi_1 _23044_ (.A1(_05137_),
    .A2(_05139_),
    .Y(_05140_),
    .B1(net9771));
 sg13g2_a21oi_1 _23045_ (.A1(\u_ac_controller_soc_inst.io_rdata[9] ),
    .A2(net9774),
    .Y(_05141_),
    .B1(_05140_));
 sg13g2_nor2_1 _23046_ (.A(net11002),
    .B(_05141_),
    .Y(_00247_));
 sg13g2_buf_16 clkbuf_leaf_378_clk (.X(clknet_leaf_378_clk),
    .A(clknet_8_120_0_clk));
 sg13g2_nand2_1 _23048_ (.Y(_05143_),
    .A(_04804_),
    .B(_04971_));
 sg13g2_buf_2 place9891 (.A(net9889),
    .X(net9891));
 sg13g2_buf_2 place10946 (.A(net10945),
    .X(net10946));
 sg13g2_buf_2 place9895 (.A(net9894),
    .X(net9895));
 sg13g2_nor2_1 _23052_ (.A(_04817_),
    .B(_05143_),
    .Y(_05147_));
 sg13g2_a21oi_1 _23053_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[0] ),
    .A2(net9761),
    .Y(_05148_),
    .B1(_05147_));
 sg13g2_nor2_1 _23054_ (.A(net10989),
    .B(_05148_),
    .Y(_00249_));
 sg13g2_nor2_1 _23055_ (.A(_04822_),
    .B(net9764),
    .Y(_05149_));
 sg13g2_a21oi_1 _23056_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[10] ),
    .A2(net9764),
    .Y(_05150_),
    .B1(_05149_));
 sg13g2_nor2_1 _23057_ (.A(net10985),
    .B(_05150_),
    .Y(_00250_));
 sg13g2_nor2_1 _23058_ (.A(_04825_),
    .B(net9764),
    .Y(_05151_));
 sg13g2_a21oi_1 _23059_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[11] ),
    .A2(net9764),
    .Y(_05152_),
    .B1(_05151_));
 sg13g2_nor2_1 _23060_ (.A(net10985),
    .B(_05152_),
    .Y(_00251_));
 sg13g2_nor2_1 _23061_ (.A(_04828_),
    .B(net9764),
    .Y(_05153_));
 sg13g2_a21oi_1 _23062_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[12] ),
    .A2(net9764),
    .Y(_05154_),
    .B1(_05153_));
 sg13g2_nor2_1 _23063_ (.A(net10985),
    .B(_05154_),
    .Y(_00252_));
 sg13g2_nor2_1 _23064_ (.A(_04832_),
    .B(net9764),
    .Y(_05155_));
 sg13g2_a21oi_1 _23065_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[13] ),
    .A2(net9765),
    .Y(_05156_),
    .B1(_05155_));
 sg13g2_nor2_1 _23066_ (.A(net10991),
    .B(_05156_),
    .Y(_00253_));
 sg13g2_nor2_1 _23067_ (.A(_04835_),
    .B(net9765),
    .Y(_05157_));
 sg13g2_a21oi_1 _23068_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[14] ),
    .A2(net9765),
    .Y(_05158_),
    .B1(_05157_));
 sg13g2_nor2_1 _23069_ (.A(net10992),
    .B(_05158_),
    .Y(_00254_));
 sg13g2_nor2_1 _23070_ (.A(_04838_),
    .B(net9765),
    .Y(_05159_));
 sg13g2_a21oi_1 _23071_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[15] ),
    .A2(net9765),
    .Y(_05160_),
    .B1(_05159_));
 sg13g2_nor2_1 _23072_ (.A(net10991),
    .B(_05160_),
    .Y(_00255_));
 sg13g2_nor2_1 _23073_ (.A(_04841_),
    .B(net9765),
    .Y(_05161_));
 sg13g2_a21oi_1 _23074_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[16] ),
    .A2(net9767),
    .Y(_05162_),
    .B1(_05161_));
 sg13g2_nor2_1 _23075_ (.A(net10994),
    .B(_05162_),
    .Y(_00256_));
 sg13g2_buf_2 place9897 (.A(_10770_),
    .X(net9897));
 sg13g2_nor2_1 _23077_ (.A(_04845_),
    .B(net9767),
    .Y(_05164_));
 sg13g2_a21oi_1 _23078_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[17] ),
    .A2(net9767),
    .Y(_05165_),
    .B1(_05164_));
 sg13g2_nor2_1 _23079_ (.A(net10992),
    .B(_05165_),
    .Y(_00257_));
 sg13g2_nor2_1 _23080_ (.A(_04848_),
    .B(net9767),
    .Y(_05166_));
 sg13g2_a21oi_1 _23081_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[18] ),
    .A2(net9767),
    .Y(_05167_),
    .B1(_05166_));
 sg13g2_nor2_1 _23082_ (.A(net10992),
    .B(_05167_),
    .Y(_00258_));
 sg13g2_buf_2 place9896 (.A(net9894),
    .X(net9896));
 sg13g2_buf_2 place9892 (.A(net9891),
    .X(net9892));
 sg13g2_nor2_1 _23085_ (.A(_04852_),
    .B(net9767),
    .Y(_05170_));
 sg13g2_a21oi_1 _23086_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[19] ),
    .A2(net9767),
    .Y(_05171_),
    .B1(_05170_));
 sg13g2_nor2_1 _23087_ (.A(net10992),
    .B(_05171_),
    .Y(_00259_));
 sg13g2_nor2_1 _23088_ (.A(_04856_),
    .B(net9761),
    .Y(_05172_));
 sg13g2_a21oi_1 _23089_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[1] ),
    .A2(net9762),
    .Y(_05173_),
    .B1(_05172_));
 sg13g2_nor2_1 _23090_ (.A(net10984),
    .B(_05173_),
    .Y(_00260_));
 sg13g2_nor2_1 _23091_ (.A(_04859_),
    .B(net9768),
    .Y(_05174_));
 sg13g2_a21oi_1 _23092_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[20] ),
    .A2(net9768),
    .Y(_05175_),
    .B1(_05174_));
 sg13g2_nor2_1 _23093_ (.A(net10995),
    .B(_05175_),
    .Y(_00261_));
 sg13g2_nor2_1 _23094_ (.A(_04862_),
    .B(net9768),
    .Y(_05176_));
 sg13g2_a21oi_1 _23095_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[21] ),
    .A2(net9768),
    .Y(_05177_),
    .B1(_05176_));
 sg13g2_nor2_1 _23096_ (.A(net10995),
    .B(_05177_),
    .Y(_00262_));
 sg13g2_nor2_1 _23097_ (.A(_04866_),
    .B(net9768),
    .Y(_05178_));
 sg13g2_a21oi_1 _23098_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[22] ),
    .A2(net9768),
    .Y(_05179_),
    .B1(_05178_));
 sg13g2_nor2_1 _23099_ (.A(net10995),
    .B(_05179_),
    .Y(_00263_));
 sg13g2_nor2_1 _23100_ (.A(_04869_),
    .B(net9768),
    .Y(_05180_));
 sg13g2_a21oi_1 _23101_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[23] ),
    .A2(net9768),
    .Y(_05181_),
    .B1(_05180_));
 sg13g2_nor2_1 _23102_ (.A(net10995),
    .B(_05181_),
    .Y(_00264_));
 sg13g2_nor2_1 _23103_ (.A(_04872_),
    .B(net9769),
    .Y(_05182_));
 sg13g2_a21oi_1 _23104_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[24] ),
    .A2(net9766),
    .Y(_05183_),
    .B1(_05182_));
 sg13g2_nor2_1 _23105_ (.A(net10998),
    .B(_05183_),
    .Y(_00265_));
 sg13g2_nor2_1 _23106_ (.A(_04875_),
    .B(net9769),
    .Y(_05184_));
 sg13g2_a21oi_1 _23107_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[25] ),
    .A2(net9769),
    .Y(_05185_),
    .B1(_05184_));
 sg13g2_nor2_1 _23108_ (.A(net10999),
    .B(_05185_),
    .Y(_00266_));
 sg13g2_buf_2 place9894 (.A(_10770_),
    .X(net9894));
 sg13g2_nor2_1 _23110_ (.A(_04879_),
    .B(net9769),
    .Y(_05187_));
 sg13g2_a21oi_1 _23111_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[26] ),
    .A2(net9769),
    .Y(_05188_),
    .B1(_05187_));
 sg13g2_nor2_1 _23112_ (.A(net10999),
    .B(_05188_),
    .Y(_00267_));
 sg13g2_nor2_1 _23113_ (.A(_04882_),
    .B(net9770),
    .Y(_05189_));
 sg13g2_a21oi_1 _23114_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[27] ),
    .A2(net9770),
    .Y(_05190_),
    .B1(_05189_));
 sg13g2_nor2_1 _23115_ (.A(net10998),
    .B(_05190_),
    .Y(_00268_));
 sg13g2_buf_2 place9890 (.A(net9889),
    .X(net9890));
 sg13g2_buf_2 place9889 (.A(_10770_),
    .X(net9889));
 sg13g2_nor2_1 _23118_ (.A(_04886_),
    .B(net9769),
    .Y(_05193_));
 sg13g2_a21oi_1 _23119_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[28] ),
    .A2(net9769),
    .Y(_05194_),
    .B1(_05193_));
 sg13g2_nor2_1 _23120_ (.A(net10999),
    .B(_05194_),
    .Y(_00269_));
 sg13g2_nor2_1 _23121_ (.A(_04890_),
    .B(net9770),
    .Y(_05195_));
 sg13g2_a21oi_1 _23122_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[29] ),
    .A2(net9770),
    .Y(_05196_),
    .B1(_05195_));
 sg13g2_nor2_1 _23123_ (.A(net10998),
    .B(_05196_),
    .Y(_00270_));
 sg13g2_nor2_1 _23124_ (.A(_04893_),
    .B(net9761),
    .Y(_05197_));
 sg13g2_a21oi_1 _23125_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[2] ),
    .A2(net9761),
    .Y(_05198_),
    .B1(_05197_));
 sg13g2_nor2_1 _23126_ (.A(net10982),
    .B(_05198_),
    .Y(_00271_));
 sg13g2_nor2_1 _23127_ (.A(_04896_),
    .B(net9770),
    .Y(_05199_));
 sg13g2_a21oi_1 _23128_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[30] ),
    .A2(net9770),
    .Y(_05200_),
    .B1(_05199_));
 sg13g2_nor2_1 _23129_ (.A(net11000),
    .B(_05200_),
    .Y(_00272_));
 sg13g2_nor2_1 _23130_ (.A(_04901_),
    .B(net9770),
    .Y(_05201_));
 sg13g2_a21oi_1 _23131_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[31] ),
    .A2(net9770),
    .Y(_05202_),
    .B1(_05201_));
 sg13g2_nor2_1 _23132_ (.A(net11000),
    .B(_05202_),
    .Y(_00273_));
 sg13g2_nor2_1 _23133_ (.A(_04904_),
    .B(net9761),
    .Y(_05203_));
 sg13g2_a21oi_1 _23134_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[3] ),
    .A2(net9761),
    .Y(_05204_),
    .B1(_05203_));
 sg13g2_nor2_1 _23135_ (.A(net10982),
    .B(_05204_),
    .Y(_00274_));
 sg13g2_nor2_1 _23136_ (.A(_04907_),
    .B(net9762),
    .Y(_05205_));
 sg13g2_a21oi_1 _23137_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[4] ),
    .A2(net9762),
    .Y(_05206_),
    .B1(_05205_));
 sg13g2_nor2_1 _23138_ (.A(net10982),
    .B(_05206_),
    .Y(_00275_));
 sg13g2_nor2_1 _23139_ (.A(_04910_),
    .B(net9762),
    .Y(_05207_));
 sg13g2_a21oi_1 _23140_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[5] ),
    .A2(net9762),
    .Y(_05208_),
    .B1(_05207_));
 sg13g2_nor2_1 _23141_ (.A(net10983),
    .B(_05208_),
    .Y(_00276_));
 sg13g2_nor2_1 _23142_ (.A(_04913_),
    .B(net9762),
    .Y(_05209_));
 sg13g2_a21oi_1 _23143_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[6] ),
    .A2(net9762),
    .Y(_05210_),
    .B1(_05209_));
 sg13g2_nor2_1 _23144_ (.A(net10983),
    .B(_05210_),
    .Y(_00277_));
 sg13g2_nor2_1 _23145_ (.A(_04916_),
    .B(net9763),
    .Y(_05211_));
 sg13g2_a21oi_1 _23146_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[7] ),
    .A2(net9763),
    .Y(_05212_),
    .B1(_05211_));
 sg13g2_nor2_1 _23147_ (.A(net10983),
    .B(_05212_),
    .Y(_00278_));
 sg13g2_buf_2 place9893 (.A(net9891),
    .X(net9893));
 sg13g2_buf_16 clkbuf_leaf_379_clk (.X(clknet_leaf_379_clk),
    .A(clknet_8_120_0_clk));
 sg13g2_nor2_1 _23150_ (.A(_04919_),
    .B(net9763),
    .Y(_05215_));
 sg13g2_a21oi_1 _23151_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[8] ),
    .A2(net9763),
    .Y(_05216_),
    .B1(_05215_));
 sg13g2_nor2_1 _23152_ (.A(net10983),
    .B(_05216_),
    .Y(_00279_));
 sg13g2_nor2_1 _23153_ (.A(_04922_),
    .B(net9763),
    .Y(_05217_));
 sg13g2_a21oi_1 _23154_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[9] ),
    .A2(net9763),
    .Y(_05218_),
    .B1(_05217_));
 sg13g2_nor2_1 _23155_ (.A(net10983),
    .B(_05218_),
    .Y(_00280_));
 sg13g2_and3_1 _23156_ (.X(_05219_),
    .A(_04804_),
    .B(_04817_),
    .C(_04953_));
 sg13g2_a21oi_1 _23157_ (.A1(_04804_),
    .A2(_04953_),
    .Y(_05220_),
    .B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_enable ));
 sg13g2_o21ai_1 _23158_ (.B1(net11038),
    .Y(_00281_),
    .A1(_05219_),
    .A2(_05220_));
 sg13g2_xor2_1 _23159_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[30] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[30] ),
    .X(_05221_));
 sg13g2_nor2b_1 _23160_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[29] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[29] ),
    .Y(_05222_));
 sg13g2_xor2_1 _23161_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[31] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[31] ),
    .X(_05223_));
 sg13g2_nor3_1 _23162_ (.A(_05221_),
    .B(_05222_),
    .C(_05223_),
    .Y(_05224_));
 sg13g2_xor2_1 _23163_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[26] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26] ),
    .X(_05225_));
 sg13g2_nor2b_1 _23164_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[25] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[25] ),
    .Y(_05226_));
 sg13g2_xor2_1 _23165_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[27] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[27] ),
    .X(_05227_));
 sg13g2_nor3_1 _23166_ (.A(_05225_),
    .B(_05226_),
    .C(_05227_),
    .Y(_05228_));
 sg13g2_nor2_1 _23167_ (.A(_04183_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[28] ),
    .Y(_05229_));
 sg13g2_inv_1 _23168_ (.Y(_05230_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[24] ));
 sg13g2_nor2b_1 _23169_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[25] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[25] ),
    .Y(_05231_));
 sg13g2_a21o_1 _23170_ (.A2(_05230_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24] ),
    .B1(_05231_),
    .X(_05232_));
 sg13g2_nor2b_1 _23171_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[28] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[28] ),
    .Y(_05233_));
 sg13g2_nand2b_1 _23172_ (.Y(_05234_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[29] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[29] ));
 sg13g2_o21ai_1 _23173_ (.B1(_05234_),
    .Y(_05235_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24] ),
    .A2(_05230_));
 sg13g2_nor4_1 _23174_ (.A(_05229_),
    .B(_05232_),
    .C(_05233_),
    .D(_05235_),
    .Y(_05236_));
 sg13g2_nand3_1 _23175_ (.B(_05228_),
    .C(_05236_),
    .A(_05224_),
    .Y(_05237_));
 sg13g2_xor2_1 _23176_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[22] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22] ),
    .X(_05238_));
 sg13g2_nor2b_1 _23177_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[21] ),
    .Y(_05239_));
 sg13g2_xor2_1 _23178_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[23] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[23] ),
    .X(_05240_));
 sg13g2_nor3_1 _23179_ (.A(_05238_),
    .B(_05239_),
    .C(_05240_),
    .Y(_05241_));
 sg13g2_o21ai_1 _23180_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[19] ),
    .Y(_05242_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[18] ),
    .A2(_04201_));
 sg13g2_o21ai_1 _23181_ (.B1(_04199_),
    .Y(_05243_),
    .A1(_04198_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[18] ));
 sg13g2_or2_1 _23182_ (.X(_05244_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[18] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[18] ));
 sg13g2_nand2_1 _23183_ (.Y(_05245_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[18] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[18] ));
 sg13g2_xor2_1 _23184_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[19] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[19] ),
    .X(_05246_));
 sg13g2_a221oi_1 _23185_ (.B2(_05245_),
    .C1(_05246_),
    .B1(_05244_),
    .A1(_04159_),
    .Y(_05247_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[17] ));
 sg13g2_nand2b_1 _23186_ (.Y(_05248_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[17] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[17] ));
 sg13g2_o21ai_1 _23187_ (.B1(_05248_),
    .Y(_05249_),
    .A1(_04152_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[16] ));
 sg13g2_nor2_1 _23188_ (.A(_04197_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[20] ),
    .Y(_05250_));
 sg13g2_a221oi_1 _23189_ (.B2(_05249_),
    .C1(_05250_),
    .B1(_05247_),
    .A1(_05242_),
    .Y(_05251_),
    .A2(_05243_));
 sg13g2_nor2b_1 _23190_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[20] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[20] ),
    .Y(_05252_));
 sg13g2_nand2b_1 _23191_ (.Y(_05253_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[21] ));
 sg13g2_o21ai_1 _23192_ (.B1(_05253_),
    .Y(_05254_),
    .A1(_05251_),
    .A2(_05252_));
 sg13g2_nand2b_1 _23193_ (.Y(_05255_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[22] ));
 sg13g2_o21ai_1 _23194_ (.B1(_04262_),
    .Y(_05256_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[23] ),
    .A2(_05255_));
 sg13g2_nand2_1 _23195_ (.Y(_05257_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[23] ),
    .B(_05255_));
 sg13g2_xor2_1 _23196_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[14] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14] ),
    .X(_05258_));
 sg13g2_nor2b_1 _23197_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[13] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[13] ),
    .Y(_05259_));
 sg13g2_xor2_1 _23198_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[15] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[15] ),
    .X(_05260_));
 sg13g2_nor3_2 _23199_ (.A(_05258_),
    .B(_05259_),
    .C(_05260_),
    .Y(_05261_));
 sg13g2_nor2b_1 _23200_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[12] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[12] ),
    .Y(_05262_));
 sg13g2_nand2b_1 _23201_ (.Y(_05263_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[10] ));
 sg13g2_nand2b_1 _23202_ (.Y(_05264_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[10] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10] ));
 sg13g2_xor2_1 _23203_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[11] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[11] ),
    .X(_05265_));
 sg13g2_a21oi_1 _23204_ (.A1(_04102_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[9] ),
    .Y(_05266_),
    .B1(_05265_));
 sg13g2_nand3_1 _23205_ (.B(_05264_),
    .C(_05266_),
    .A(_05263_),
    .Y(_05267_));
 sg13g2_inv_1 _23206_ (.Y(_05268_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[8] ));
 sg13g2_inv_1 _23207_ (.Y(_05269_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[9] ));
 sg13g2_a22oi_1 _23208_ (.Y(_05270_),
    .B1(_05269_),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9] ),
    .A2(_05268_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[8] ));
 sg13g2_nor2_1 _23209_ (.A(_05267_),
    .B(_05270_),
    .Y(_05271_));
 sg13g2_o21ai_1 _23210_ (.B1(_04090_),
    .Y(_05272_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[11] ),
    .A2(_05263_));
 sg13g2_nand2_1 _23211_ (.Y(_05273_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[11] ),
    .B(_05263_));
 sg13g2_and2_1 _23212_ (.A(_05272_),
    .B(_05273_),
    .X(_05274_));
 sg13g2_nor2_1 _23213_ (.A(_04094_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[12] ),
    .Y(_05275_));
 sg13g2_nor3_1 _23214_ (.A(_05271_),
    .B(_05274_),
    .C(_05275_),
    .Y(_05276_));
 sg13g2_nand2b_1 _23215_ (.Y(_05277_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[13] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[13] ));
 sg13g2_o21ai_1 _23216_ (.B1(_05277_),
    .Y(_05278_),
    .A1(_05262_),
    .A2(_05276_));
 sg13g2_nand2b_1 _23217_ (.Y(_05279_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[14] ));
 sg13g2_o21ai_1 _23218_ (.B1(_04242_),
    .Y(_05280_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[15] ),
    .A2(_05279_));
 sg13g2_nand2_1 _23219_ (.Y(_05281_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[15] ),
    .B(_05279_));
 sg13g2_a22oi_1 _23220_ (.Y(_05282_),
    .B1(_05280_),
    .B2(_05281_),
    .A2(_05278_),
    .A1(_05261_));
 sg13g2_nand2b_1 _23221_ (.Y(_05283_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[6] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[6] ));
 sg13g2_nand2b_1 _23222_ (.Y(_05284_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[6] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[6] ));
 sg13g2_xor2_1 _23223_ (.B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[7] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[7] ),
    .X(_05285_));
 sg13g2_a21oi_1 _23224_ (.A1(_04053_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[5] ),
    .Y(_05286_),
    .B1(_05285_));
 sg13g2_and3_2 _23225_ (.X(_05287_),
    .A(_05283_),
    .B(_05284_),
    .C(_05286_));
 sg13g2_inv_1 _23226_ (.Y(_05288_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[3] ));
 sg13g2_nand2b_1 _23227_ (.Y(_05289_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[2] ));
 sg13g2_nor2b_2 _23228_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[0] ),
    .Y(_05290_));
 sg13g2_nor2_1 _23229_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[1] ),
    .B(_05290_),
    .Y(_05291_));
 sg13g2_a21oi_1 _23230_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[1] ),
    .A2(_05290_),
    .Y(_05292_),
    .B1(_04063_));
 sg13g2_nor2_1 _23231_ (.A(_05291_),
    .B(_05292_),
    .Y(_05293_));
 sg13g2_nor2b_1 _23232_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[2] ),
    .Y(_05294_));
 sg13g2_a221oi_1 _23233_ (.B2(_05293_),
    .C1(_05294_),
    .B1(_05289_),
    .A1(_04070_),
    .Y(_05295_),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[3] ));
 sg13g2_a21oi_1 _23234_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[3] ),
    .A2(_05288_),
    .Y(_05296_),
    .B1(_05295_));
 sg13g2_inv_1 _23235_ (.Y(_05297_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[4] ));
 sg13g2_nor2_1 _23236_ (.A(net10761),
    .B(_05297_),
    .Y(_05298_));
 sg13g2_nor2_1 _23237_ (.A(_04053_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[5] ),
    .Y(_05299_));
 sg13g2_a21oi_1 _23238_ (.A1(net10761),
    .A2(_05297_),
    .Y(_05300_),
    .B1(_05299_));
 sg13g2_o21ai_1 _23239_ (.B1(_05300_),
    .Y(_05301_),
    .A1(_05296_),
    .A2(_05298_));
 sg13g2_nand2_1 _23240_ (.Y(_05302_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[7] ),
    .B(_05283_));
 sg13g2_o21ai_1 _23241_ (.B1(_04051_),
    .Y(_05303_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[7] ),
    .A2(_05283_));
 sg13g2_a22oi_1 _23242_ (.Y(_05304_),
    .B1(_05302_),
    .B2(_05303_),
    .A2(_05301_),
    .A1(_05287_));
 sg13g2_nand2_1 _23243_ (.Y(_05305_),
    .A(_04082_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[8] ));
 sg13g2_nand3_1 _23244_ (.B(_05270_),
    .C(_05305_),
    .A(_05277_),
    .Y(_05306_));
 sg13g2_nor4_1 _23245_ (.A(_05267_),
    .B(_05262_),
    .C(_05275_),
    .D(_05306_),
    .Y(_05307_));
 sg13g2_nand3b_1 _23246_ (.B(_05307_),
    .C(_05261_),
    .Y(_05308_),
    .A_N(_05304_));
 sg13g2_xnor2_1 _23247_ (.Y(_05309_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[16] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[16] ));
 sg13g2_nand3_1 _23248_ (.B(_05248_),
    .C(_05309_),
    .A(_05253_),
    .Y(_05310_));
 sg13g2_nor3_1 _23249_ (.A(_05250_),
    .B(_05252_),
    .C(_05310_),
    .Y(_05311_));
 sg13g2_nand3_1 _23250_ (.B(_05247_),
    .C(_05311_),
    .A(_05241_),
    .Y(_05312_));
 sg13g2_a21oi_2 _23251_ (.B1(_05312_),
    .Y(_05313_),
    .A2(_05308_),
    .A1(_05282_));
 sg13g2_a221oi_1 _23252_ (.B2(_05257_),
    .C1(_05313_),
    .B1(_05256_),
    .A1(_05241_),
    .Y(_05314_),
    .A2(_05254_));
 sg13g2_nand2b_1 _23253_ (.Y(_05315_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[26] ));
 sg13g2_o21ai_1 _23254_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[27] ),
    .Y(_05316_),
    .A1(_04184_),
    .A2(_05315_));
 sg13g2_nand2_1 _23255_ (.Y(_05317_),
    .A(_04184_),
    .B(_05315_));
 sg13g2_a221oi_1 _23256_ (.B2(_05232_),
    .C1(_05229_),
    .B1(_05228_),
    .A1(_05316_),
    .Y(_05318_),
    .A2(_05317_));
 sg13g2_o21ai_1 _23257_ (.B1(_05234_),
    .Y(_05319_),
    .A1(_05318_),
    .A2(_05233_));
 sg13g2_nand2b_1 _23258_ (.Y(_05320_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[30] ),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[30] ));
 sg13g2_o21ai_1 _23259_ (.B1(_04111_),
    .Y(_05321_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[31] ),
    .A2(_05320_));
 sg13g2_nand2_1 _23260_ (.Y(_05322_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[31] ),
    .B(_05320_));
 sg13g2_a22oi_1 _23261_ (.Y(_05323_),
    .B1(_05321_),
    .B2(_05322_),
    .A2(_05319_),
    .A1(_05224_));
 sg13g2_o21ai_1 _23262_ (.B1(_05323_),
    .Y(_05324_),
    .A1(_05237_),
    .A2(_05314_));
 sg13g2_nor2b_1 _23263_ (.A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[0] ),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0] ),
    .Y(_05325_));
 sg13g2_xnor2_1 _23264_ (.Y(_05326_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[3] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[3] ));
 sg13g2_xnor2_1 _23265_ (.Y(_05327_),
    .A(net10761),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[4] ));
 sg13g2_xnor2_1 _23266_ (.Y(_05328_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[1] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[1] ));
 sg13g2_xnor2_1 _23267_ (.Y(_05329_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[2] ));
 sg13g2_nand4_1 _23268_ (.B(_05327_),
    .C(_05328_),
    .A(_05326_),
    .Y(_05330_),
    .D(_05329_));
 sg13g2_nor4_2 _23269_ (.A(_05299_),
    .B(_05290_),
    .C(_05325_),
    .Y(_05331_),
    .D(_05330_));
 sg13g2_nand4_1 _23270_ (.B(_05307_),
    .C(_05287_),
    .A(_05261_),
    .Y(_05332_),
    .D(_05331_));
 sg13g2_or3_1 _23271_ (.A(_05237_),
    .B(_05312_),
    .C(_05332_),
    .X(_05333_));
 sg13g2_a21oi_2 _23272_ (.B1(_04218_),
    .Y(_00282_),
    .A2(_05333_),
    .A1(_05324_));
 sg13g2_nand2_2 _23273_ (.Y(_05334_),
    .A(_04804_),
    .B(_04974_));
 sg13g2_buf_2 place9883 (.A(net9881),
    .X(net9883));
 sg13g2_buf_2 place9881 (.A(_10850_),
    .X(net9881));
 sg13g2_buf_2 place10939 (.A(net10935),
    .X(net10939));
 sg13g2_nor2_1 _23277_ (.A(_04817_),
    .B(_05334_),
    .Y(_05338_));
 sg13g2_a21oi_1 _23278_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[0] ),
    .A2(_05334_),
    .Y(_05339_),
    .B1(_05338_));
 sg13g2_nor2_1 _23279_ (.A(net10989),
    .B(_05339_),
    .Y(_00283_));
 sg13g2_nor2_1 _23280_ (.A(_04822_),
    .B(net9754),
    .Y(_05340_));
 sg13g2_a21oi_1 _23281_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[10] ),
    .A2(net9754),
    .Y(_05341_),
    .B1(_05340_));
 sg13g2_nor2_1 _23282_ (.A(net10985),
    .B(_05341_),
    .Y(_00284_));
 sg13g2_nor2_1 _23283_ (.A(_04825_),
    .B(net9754),
    .Y(_05342_));
 sg13g2_a21oi_1 _23284_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[11] ),
    .A2(net9754),
    .Y(_05343_),
    .B1(_05342_));
 sg13g2_nor2_1 _23285_ (.A(net10985),
    .B(_05343_),
    .Y(_00285_));
 sg13g2_nor2_1 _23286_ (.A(_04828_),
    .B(net9754),
    .Y(_05344_));
 sg13g2_a21oi_1 _23287_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[12] ),
    .A2(net9754),
    .Y(_05345_),
    .B1(_05344_));
 sg13g2_nor2_1 _23288_ (.A(net11002),
    .B(_05345_),
    .Y(_00286_));
 sg13g2_nor2_1 _23289_ (.A(_04832_),
    .B(net9755),
    .Y(_05346_));
 sg13g2_a21oi_1 _23290_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[13] ),
    .A2(net9755),
    .Y(_05347_),
    .B1(_05346_));
 sg13g2_nor2_1 _23291_ (.A(net10991),
    .B(_05347_),
    .Y(_00287_));
 sg13g2_nor2_1 _23292_ (.A(_04835_),
    .B(net9755),
    .Y(_05348_));
 sg13g2_a21oi_1 _23293_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[14] ),
    .A2(net9755),
    .Y(_05349_),
    .B1(_05348_));
 sg13g2_nor2_1 _23294_ (.A(net10991),
    .B(_05349_),
    .Y(_00288_));
 sg13g2_nor2_1 _23295_ (.A(_04838_),
    .B(net9755),
    .Y(_05350_));
 sg13g2_a21oi_1 _23296_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[15] ),
    .A2(net9755),
    .Y(_05351_),
    .B1(_05350_));
 sg13g2_nor2_1 _23297_ (.A(net10991),
    .B(_05351_),
    .Y(_00289_));
 sg13g2_nor2_1 _23298_ (.A(_04841_),
    .B(net9756),
    .Y(_05352_));
 sg13g2_a21oi_1 _23299_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[16] ),
    .A2(net9757),
    .Y(_05353_),
    .B1(_05352_));
 sg13g2_nor2_1 _23300_ (.A(net10994),
    .B(_05353_),
    .Y(_00290_));
 sg13g2_buf_2 place9886 (.A(_10850_),
    .X(net9886));
 sg13g2_buf_2 place9925 (.A(net9922),
    .X(net9925));
 sg13g2_nor2_1 _23303_ (.A(_04845_),
    .B(net9756),
    .Y(_05356_));
 sg13g2_a21oi_1 _23304_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[17] ),
    .A2(net9756),
    .Y(_05357_),
    .B1(_05356_));
 sg13g2_nor2_1 _23305_ (.A(net10994),
    .B(_05357_),
    .Y(_00291_));
 sg13g2_nor2_1 _23306_ (.A(_04848_),
    .B(net9756),
    .Y(_05358_));
 sg13g2_a21oi_1 _23307_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[18] ),
    .A2(net9756),
    .Y(_05359_),
    .B1(_05358_));
 sg13g2_nor2_1 _23308_ (.A(net10992),
    .B(_05359_),
    .Y(_00292_));
 sg13g2_buf_2 place9885 (.A(_10850_),
    .X(net9885));
 sg13g2_nor2_1 _23310_ (.A(_04852_),
    .B(net9756),
    .Y(_05361_));
 sg13g2_a21oi_1 _23311_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[19] ),
    .A2(net9756),
    .Y(_05362_),
    .B1(_05361_));
 sg13g2_nor2_1 _23312_ (.A(net10992),
    .B(_05362_),
    .Y(_00293_));
 sg13g2_nor2_1 _23313_ (.A(_04856_),
    .B(_05334_),
    .Y(_05363_));
 sg13g2_a21oi_1 _23314_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[1] ),
    .A2(_05334_),
    .Y(_05364_),
    .B1(_05363_));
 sg13g2_nor2_1 _23315_ (.A(net10981),
    .B(_05364_),
    .Y(_00294_));
 sg13g2_nor2_1 _23316_ (.A(_04859_),
    .B(net9757),
    .Y(_05365_));
 sg13g2_a21oi_1 _23317_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[20] ),
    .A2(net9757),
    .Y(_05366_),
    .B1(_05365_));
 sg13g2_nor2_1 _23318_ (.A(net10995),
    .B(_05366_),
    .Y(_00295_));
 sg13g2_nor2_1 _23319_ (.A(_04862_),
    .B(net9758),
    .Y(_05367_));
 sg13g2_a21oi_1 _23320_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[21] ),
    .A2(net9758),
    .Y(_05368_),
    .B1(_05367_));
 sg13g2_nor2_1 _23321_ (.A(net10995),
    .B(_05368_),
    .Y(_00296_));
 sg13g2_nor2_1 _23322_ (.A(_04866_),
    .B(net9757),
    .Y(_05369_));
 sg13g2_a21oi_1 _23323_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[22] ),
    .A2(net9757),
    .Y(_05370_),
    .B1(_05369_));
 sg13g2_nor2_1 _23324_ (.A(net10995),
    .B(_05370_),
    .Y(_00297_));
 sg13g2_nor2_1 _23325_ (.A(_04869_),
    .B(net9757),
    .Y(_05371_));
 sg13g2_a21oi_1 _23326_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[23] ),
    .A2(net9757),
    .Y(_05372_),
    .B1(_05371_));
 sg13g2_nor2_1 _23327_ (.A(net10995),
    .B(_05372_),
    .Y(_00298_));
 sg13g2_nor2_1 _23328_ (.A(_04872_),
    .B(net9758),
    .Y(_05373_));
 sg13g2_a21oi_1 _23329_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[24] ),
    .A2(net9759),
    .Y(_05374_),
    .B1(_05373_));
 sg13g2_nor2_1 _23330_ (.A(net10998),
    .B(_05374_),
    .Y(_00299_));
 sg13g2_nor2_1 _23331_ (.A(_04875_),
    .B(net9758),
    .Y(_05375_));
 sg13g2_a21oi_1 _23332_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[25] ),
    .A2(net9758),
    .Y(_05376_),
    .B1(_05375_));
 sg13g2_nor2_1 _23333_ (.A(net10999),
    .B(_05376_),
    .Y(_00300_));
 sg13g2_buf_2 place9884 (.A(_10850_),
    .X(net9884));
 sg13g2_buf_2 place9888 (.A(net9886),
    .X(net9888));
 sg13g2_nor2_1 _23336_ (.A(_04879_),
    .B(net9759),
    .Y(_05379_));
 sg13g2_a21oi_1 _23337_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[26] ),
    .A2(net9759),
    .Y(_05380_),
    .B1(_05379_));
 sg13g2_nor2_1 _23338_ (.A(net10999),
    .B(_05380_),
    .Y(_00301_));
 sg13g2_nor2_1 _23339_ (.A(_04882_),
    .B(net9759),
    .Y(_05381_));
 sg13g2_a21oi_1 _23340_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[27] ),
    .A2(net9759),
    .Y(_05382_),
    .B1(_05381_));
 sg13g2_nor2_1 _23341_ (.A(net10999),
    .B(_05382_),
    .Y(_00302_));
 sg13g2_buf_2 place9887 (.A(net9886),
    .X(net9887));
 sg13g2_nor2_1 _23343_ (.A(_04886_),
    .B(net9759),
    .Y(_05384_));
 sg13g2_a21oi_1 _23344_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[28] ),
    .A2(net9760),
    .Y(_05385_),
    .B1(_05384_));
 sg13g2_nor2_1 _23345_ (.A(net10999),
    .B(_05385_),
    .Y(_00303_));
 sg13g2_nor2_1 _23346_ (.A(_04890_),
    .B(net9760),
    .Y(_05386_));
 sg13g2_a21oi_1 _23347_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[29] ),
    .A2(net9760),
    .Y(_05387_),
    .B1(_05386_));
 sg13g2_nor2_1 _23348_ (.A(net10999),
    .B(_05387_),
    .Y(_00304_));
 sg13g2_nor2_1 _23349_ (.A(_04893_),
    .B(_05334_),
    .Y(_05388_));
 sg13g2_a21oi_1 _23350_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[2] ),
    .A2(_05334_),
    .Y(_05389_),
    .B1(_05388_));
 sg13g2_nor2_1 _23351_ (.A(net10982),
    .B(_05389_),
    .Y(_00305_));
 sg13g2_nor2_1 _23352_ (.A(_04896_),
    .B(net9760),
    .Y(_05390_));
 sg13g2_a21oi_1 _23353_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[30] ),
    .A2(net9760),
    .Y(_05391_),
    .B1(_05390_));
 sg13g2_nor2_1 _23354_ (.A(net11000),
    .B(_05391_),
    .Y(_00306_));
 sg13g2_nor2_1 _23355_ (.A(_04901_),
    .B(net9760),
    .Y(_05392_));
 sg13g2_a21oi_1 _23356_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[31] ),
    .A2(net9760),
    .Y(_05393_),
    .B1(_05392_));
 sg13g2_nor2_1 _23357_ (.A(net11000),
    .B(_05393_),
    .Y(_00307_));
 sg13g2_nor2_1 _23358_ (.A(_04904_),
    .B(net9752),
    .Y(_05394_));
 sg13g2_a21oi_1 _23359_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[3] ),
    .A2(net9752),
    .Y(_05395_),
    .B1(_05394_));
 sg13g2_nor2_1 _23360_ (.A(net10982),
    .B(_05395_),
    .Y(_00308_));
 sg13g2_nor2_1 _23361_ (.A(_04907_),
    .B(net9752),
    .Y(_05396_));
 sg13g2_a21oi_1 _23362_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[4] ),
    .A2(net9752),
    .Y(_05397_),
    .B1(_05396_));
 sg13g2_nor2_1 _23363_ (.A(net10982),
    .B(_05397_),
    .Y(_00309_));
 sg13g2_nor2_1 _23364_ (.A(_04910_),
    .B(net9752),
    .Y(_05398_));
 sg13g2_a21oi_1 _23365_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[5] ),
    .A2(net9753),
    .Y(_05399_),
    .B1(_05398_));
 sg13g2_nor2_1 _23366_ (.A(net10982),
    .B(_05399_),
    .Y(_00310_));
 sg13g2_buf_2 place9882 (.A(net9881),
    .X(net9882));
 sg13g2_nor2_1 _23368_ (.A(_04913_),
    .B(net9753),
    .Y(_05401_));
 sg13g2_a21oi_1 _23369_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[6] ),
    .A2(net9753),
    .Y(_05402_),
    .B1(_05401_));
 sg13g2_nor2_1 _23370_ (.A(net10983),
    .B(_05402_),
    .Y(_00311_));
 sg13g2_nor2_1 _23371_ (.A(_04916_),
    .B(net9753),
    .Y(_05403_));
 sg13g2_a21oi_1 _23372_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[7] ),
    .A2(net9753),
    .Y(_05404_),
    .B1(_05403_));
 sg13g2_nor2_1 _23373_ (.A(net10983),
    .B(_05404_),
    .Y(_00312_));
 sg13g2_nor2_1 _23374_ (.A(_04919_),
    .B(net9753),
    .Y(_05405_));
 sg13g2_a21oi_1 _23375_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[8] ),
    .A2(net9753),
    .Y(_05406_),
    .B1(_05405_));
 sg13g2_nor2_1 _23376_ (.A(net10983),
    .B(_05406_),
    .Y(_00313_));
 sg13g2_nor2_1 _23377_ (.A(_04922_),
    .B(net9754),
    .Y(_05407_));
 sg13g2_a21oi_1 _23378_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[9] ),
    .A2(net9754),
    .Y(_05408_),
    .B1(_05407_));
 sg13g2_nor2_1 _23379_ (.A(net10985),
    .B(_05408_),
    .Y(_00314_));
 sg13g2_xnor2_1 _23380_ (.Y(_05409_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[0] ),
    .B(spi_sensor_clk));
 sg13g2_nor2_1 _23381_ (.A(net11004),
    .B(_05409_),
    .Y(_00315_));
 sg13g2_nand2_1 _23382_ (.Y(_05410_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[0] ),
    .B(spi_sensor_clk));
 sg13g2_xor2_1 _23383_ (.B(_05410_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[1] ),
    .X(_05411_));
 sg13g2_nor2_1 _23384_ (.A(net11004),
    .B(_05411_),
    .Y(_00316_));
 sg13g2_nand3_1 _23385_ (.B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[0] ),
    .C(spi_sensor_clk),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[1] ),
    .Y(_05412_));
 sg13g2_xnor2_1 _23386_ (.Y(_05413_),
    .A(_04319_),
    .B(_05412_));
 sg13g2_nor2_1 _23387_ (.A(net11005),
    .B(_05413_),
    .Y(_00317_));
 sg13g2_nor2_2 _23388_ (.A(_04319_),
    .B(_05412_),
    .Y(_05414_));
 sg13g2_or2_1 _23389_ (.X(_05415_),
    .B(_04331_),
    .A(spi_sensor_clk));
 sg13g2_buf_2 place9880 (.A(net9878),
    .X(net9880));
 sg13g2_nand3b_1 _23391_ (.B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3] ),
    .C(_05415_),
    .Y(_05417_),
    .A_N(_05414_));
 sg13g2_nand2b_1 _23392_ (.Y(_05418_),
    .B(_05414_),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3] ));
 sg13g2_a21oi_1 _23393_ (.A1(_05417_),
    .A2(_05418_),
    .Y(_00318_),
    .B1(net11005));
 sg13g2_nand2_1 _23394_ (.Y(_05419_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3] ),
    .B(_05414_));
 sg13g2_xnor2_1 _23395_ (.Y(_05420_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[4] ),
    .B(_05419_));
 sg13g2_and3_1 _23396_ (.X(_00319_),
    .A(net11037),
    .B(_05415_),
    .C(_05420_));
 sg13g2_nand3_1 _23397_ (.B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[4] ),
    .C(_05414_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3] ),
    .Y(_05421_));
 sg13g2_and2_1 _23398_ (.A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[5] ),
    .B(_05421_),
    .X(_05422_));
 sg13g2_nor2_1 _23399_ (.A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[5] ),
    .B(_05421_),
    .Y(_05423_));
 sg13g2_a21oi_1 _23400_ (.A1(_05415_),
    .A2(_05422_),
    .Y(_05424_),
    .B1(_05423_));
 sg13g2_nor2_1 _23401_ (.A(net11005),
    .B(_05424_),
    .Y(_00320_));
 sg13g2_nor3_2 _23402_ (.A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[5] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[4] ),
    .Y(_05425_));
 sg13g2_nor4_2 _23403_ (.A(spi_sensor_clk),
    .B(_04295_),
    .C(_04554_),
    .Y(_05426_),
    .D(_05425_));
 sg13g2_buf_2 place10001 (.A(net10000),
    .X(net10001));
 sg13g2_buf_2 place9875 (.A(net9874),
    .X(net9875));
 sg13g2_nand2_1 _23406_ (.Y(_05429_),
    .A(spi_sensor_miso),
    .B(net9989));
 sg13g2_buf_2 place9872 (.A(_10932_),
    .X(net9872));
 sg13g2_nand4_1 _23408_ (.B(_00104_),
    .C(_07881_),
    .A(\u_ac_controller_soc_inst.cbus_addr[8] ),
    .Y(_05431_),
    .D(_07882_));
 sg13g2_nor4_2 _23409_ (.A(_00105_),
    .B(_07872_),
    .C(_07880_),
    .Y(_05432_),
    .D(_05431_));
 sg13g2_nand3_1 _23410_ (.B(_04559_),
    .C(_05432_),
    .A(_07887_),
    .Y(_05433_));
 sg13g2_buf_2 place9879 (.A(net9878),
    .X(net9879));
 sg13g2_mux2_1 _23412_ (.A0(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[0] ),
    .A1(_08413_),
    .S(_05433_),
    .X(_05435_));
 sg13g2_nand2b_1 _23413_ (.Y(_05436_),
    .B(_05435_),
    .A_N(net9989));
 sg13g2_a21oi_1 _23414_ (.A1(_05429_),
    .A2(_05436_),
    .Y(_00321_),
    .B1(net10988));
 sg13g2_inv_1 _23415_ (.Y(_05437_),
    .A(_05433_));
 sg13g2_nor3_2 _23416_ (.A(_04295_),
    .B(_05426_),
    .C(_05437_),
    .Y(_05438_));
 sg13g2_buf_2 place9877 (.A(net9876),
    .X(net9877));
 sg13g2_buf_2 place9876 (.A(net9874),
    .X(net9876));
 sg13g2_a22oi_1 _23419_ (.Y(_05441_),
    .B1(net9749),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[10] ),
    .A2(net9990),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[9] ));
 sg13g2_nor2_1 _23420_ (.A(net11005),
    .B(_05441_),
    .Y(_00322_));
 sg13g2_a22oi_1 _23421_ (.Y(_05442_),
    .B1(net9749),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[11] ),
    .A2(net9990),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[10] ));
 sg13g2_nor2_1 _23422_ (.A(net11005),
    .B(_05442_),
    .Y(_00323_));
 sg13g2_buf_2 place9874 (.A(_10932_),
    .X(net9874));
 sg13g2_a22oi_1 _23424_ (.Y(_05444_),
    .B1(net9749),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[12] ),
    .A2(net9990),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[11] ));
 sg13g2_nor2_1 _23425_ (.A(net11006),
    .B(_05444_),
    .Y(_00324_));
 sg13g2_a22oi_1 _23426_ (.Y(_05445_),
    .B1(net9749),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[13] ),
    .A2(net9990),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[12] ));
 sg13g2_nor2_1 _23427_ (.A(net11006),
    .B(_05445_),
    .Y(_00325_));
 sg13g2_a22oi_1 _23428_ (.Y(_05446_),
    .B1(net9749),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[14] ),
    .A2(net9990),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[13] ));
 sg13g2_nor2_1 _23429_ (.A(net11006),
    .B(_05446_),
    .Y(_00326_));
 sg13g2_a22oi_1 _23430_ (.Y(_05447_),
    .B1(net9751),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[15] ),
    .A2(net9992),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[14] ));
 sg13g2_nor2_1 _23431_ (.A(net11008),
    .B(_05447_),
    .Y(_00327_));
 sg13g2_a22oi_1 _23432_ (.Y(_05448_),
    .B1(net9751),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[16] ),
    .A2(net9992),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[15] ));
 sg13g2_nor2_1 _23433_ (.A(net11008),
    .B(_05448_),
    .Y(_00328_));
 sg13g2_a22oi_1 _23434_ (.Y(_05449_),
    .B1(net9751),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[17] ),
    .A2(net9992),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[16] ));
 sg13g2_nor2_1 _23435_ (.A(net11008),
    .B(_05449_),
    .Y(_00329_));
 sg13g2_buf_2 place9878 (.A(_10932_),
    .X(net9878));
 sg13g2_a22oi_1 _23437_ (.Y(_05451_),
    .B1(net9751),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[18] ),
    .A2(net9992),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[17] ));
 sg13g2_nor2_1 _23438_ (.A(net11008),
    .B(_05451_),
    .Y(_00330_));
 sg13g2_a22oi_1 _23439_ (.Y(_05452_),
    .B1(net9751),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[19] ),
    .A2(net9992),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[18] ));
 sg13g2_nor2_1 _23440_ (.A(net11008),
    .B(_05452_),
    .Y(_00331_));
 sg13g2_nand2_1 _23441_ (.Y(_05453_),
    .A(\u_ac_controller_soc_inst.spi_sensor_rdata[0] ),
    .B(net9989));
 sg13g2_inv_1 _23442_ (.Y(_05454_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[1] ));
 sg13g2_nand3_1 _23443_ (.B(_07887_),
    .C(_05433_),
    .A(\u_ac_controller_soc_inst.spi_sensor_rdata[1] ),
    .Y(_05455_));
 sg13g2_o21ai_1 _23444_ (.B1(_05455_),
    .Y(_05456_),
    .A1(_05454_),
    .A2(_05433_));
 sg13g2_nand2b_1 _23445_ (.Y(_05457_),
    .B(_05456_),
    .A_N(_05426_));
 sg13g2_a21oi_1 _23446_ (.A1(_05453_),
    .A2(_05457_),
    .Y(_00332_),
    .B1(net10988));
 sg13g2_buf_2 place9873 (.A(net9872),
    .X(net9873));
 sg13g2_a22oi_1 _23448_ (.Y(_05459_),
    .B1(net9751),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[20] ),
    .A2(net9992),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[19] ));
 sg13g2_nor2_1 _23449_ (.A(net11008),
    .B(_05459_),
    .Y(_00333_));
 sg13g2_a22oi_1 _23450_ (.Y(_05460_),
    .B1(net9750),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[21] ),
    .A2(net9991),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[20] ));
 sg13g2_nor2_1 _23451_ (.A(net11007),
    .B(_05460_),
    .Y(_00334_));
 sg13g2_buf_2 place9936 (.A(_10375_),
    .X(net9936));
 sg13g2_a22oi_1 _23453_ (.Y(_05462_),
    .B1(net9751),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[22] ),
    .A2(net9992),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[21] ));
 sg13g2_nor2_1 _23454_ (.A(net11007),
    .B(_05462_),
    .Y(_00335_));
 sg13g2_a22oi_1 _23455_ (.Y(_05463_),
    .B1(net9751),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[23] ),
    .A2(net9992),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[22] ));
 sg13g2_nor2_1 _23456_ (.A(net11008),
    .B(_05463_),
    .Y(_00336_));
 sg13g2_a22oi_1 _23457_ (.Y(_05464_),
    .B1(net9749),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[24] ),
    .A2(net9990),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[23] ));
 sg13g2_nor2_1 _23458_ (.A(net11006),
    .B(_05464_),
    .Y(_00337_));
 sg13g2_a22oi_1 _23459_ (.Y(_05465_),
    .B1(net9749),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[25] ),
    .A2(net9990),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[24] ));
 sg13g2_nor2_1 _23460_ (.A(net11006),
    .B(_05465_),
    .Y(_00338_));
 sg13g2_a22oi_1 _23461_ (.Y(_05466_),
    .B1(net9750),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[26] ),
    .A2(net9991),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[25] ));
 sg13g2_nor2_1 _23462_ (.A(net11006),
    .B(_05466_),
    .Y(_00339_));
 sg13g2_a22oi_1 _23463_ (.Y(_05467_),
    .B1(net9750),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[27] ),
    .A2(net9991),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[26] ));
 sg13g2_nor2_1 _23464_ (.A(net11007),
    .B(_05467_),
    .Y(_00340_));
 sg13g2_buf_2 place9869 (.A(net9868),
    .X(net9869));
 sg13g2_a22oi_1 _23466_ (.Y(_05469_),
    .B1(net9750),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[28] ),
    .A2(net9991),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[27] ));
 sg13g2_nor2_1 _23467_ (.A(net11007),
    .B(_05469_),
    .Y(_00341_));
 sg13g2_a22oi_1 _23468_ (.Y(_05470_),
    .B1(net9750),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[29] ),
    .A2(net9991),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[28] ));
 sg13g2_nor2_1 _23469_ (.A(net11007),
    .B(_05470_),
    .Y(_00342_));
 sg13g2_buf_2 place10025 (.A(_11043_),
    .X(net10025));
 sg13g2_a22oi_1 _23471_ (.Y(_05472_),
    .B1(_05438_),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[2] ),
    .A2(_05426_),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[1] ));
 sg13g2_nor2_1 _23472_ (.A(net10987),
    .B(_05472_),
    .Y(_00343_));
 sg13g2_a22oi_1 _23473_ (.Y(_05473_),
    .B1(net9750),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[30] ),
    .A2(net9991),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[29] ));
 sg13g2_nor2_1 _23474_ (.A(net11007),
    .B(_05473_),
    .Y(_00344_));
 sg13g2_buf_2 place9868 (.A(_11083_),
    .X(net9868));
 sg13g2_a22oi_1 _23476_ (.Y(_05475_),
    .B1(net9750),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[31] ),
    .A2(net9991),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[30] ));
 sg13g2_nor2_1 _23477_ (.A(net11007),
    .B(_05475_),
    .Y(_00345_));
 sg13g2_a22oi_1 _23478_ (.Y(_05476_),
    .B1(_05438_),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[3] ),
    .A2(_05426_),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[2] ));
 sg13g2_nor2_1 _23479_ (.A(net10987),
    .B(_05476_),
    .Y(_00346_));
 sg13g2_a22oi_1 _23480_ (.Y(_05477_),
    .B1(_05438_),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[4] ),
    .A2(_05426_),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[3] ));
 sg13g2_nor2_1 _23481_ (.A(net10988),
    .B(_05477_),
    .Y(_00347_));
 sg13g2_a22oi_1 _23482_ (.Y(_05478_),
    .B1(net9748),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[5] ),
    .A2(net9989),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[4] ));
 sg13g2_nor2_1 _23483_ (.A(net10988),
    .B(_05478_),
    .Y(_00348_));
 sg13g2_a22oi_1 _23484_ (.Y(_05479_),
    .B1(net9748),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[6] ),
    .A2(net9989),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[5] ));
 sg13g2_nor2_1 _23485_ (.A(net10988),
    .B(_05479_),
    .Y(_00349_));
 sg13g2_a22oi_1 _23486_ (.Y(_05480_),
    .B1(net9748),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[7] ),
    .A2(net9989),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[6] ));
 sg13g2_nor2_1 _23487_ (.A(net10988),
    .B(_05480_),
    .Y(_00350_));
 sg13g2_a22oi_1 _23488_ (.Y(_05481_),
    .B1(net9748),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[8] ),
    .A2(net9989),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[7] ));
 sg13g2_nor2_1 _23489_ (.A(net10988),
    .B(_05481_),
    .Y(_00351_));
 sg13g2_a22oi_1 _23490_ (.Y(_05482_),
    .B1(net9748),
    .B2(\u_ac_controller_soc_inst.spi_sensor_rdata[9] ),
    .A2(net9989),
    .A1(\u_ac_controller_soc_inst.spi_sensor_rdata[8] ));
 sg13g2_nor2_1 _23491_ (.A(net11005),
    .B(_05482_),
    .Y(_00352_));
 sg13g2_buf_2 place9867 (.A(net9864),
    .X(net9867));
 sg13g2_buf_2 place9864 (.A(_11083_),
    .X(net9864));
 sg13g2_nand2b_1 _23494_ (.Y(_05485_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[0] ),
    .A_N(net10748));
 sg13g2_buf_2 place9866 (.A(net9865),
    .X(net9866));
 sg13g2_buf_2 place9853 (.A(_11123_),
    .X(net9853));
 sg13g2_o21ai_1 _23497_ (.B1(net10747),
    .Y(_05488_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[39] ),
    .A2(_04295_));
 sg13g2_and3_1 _23498_ (.X(_05489_),
    .A(net10736),
    .B(_05485_),
    .C(_05488_));
 sg13g2_nor3_1 _23499_ (.A(net10736),
    .B(\u_ac_controller_soc_inst.cbus_wdata[24] ),
    .C(net10149),
    .Y(_05490_));
 sg13g2_buf_2 place10376 (.A(net10372),
    .X(net10376));
 sg13g2_buf_2 place9861 (.A(net9858),
    .X(net9861));
 sg13g2_o21ai_1 _23502_ (.B1(net11039),
    .Y(_05493_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[0] ),
    .A2(net10237));
 sg13g2_nor3_1 _23503_ (.A(_05489_),
    .B(_05490_),
    .C(_05493_),
    .Y(_00353_));
 sg13g2_nand2b_1 _23504_ (.Y(_05494_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[10] ),
    .A_N(net10759));
 sg13g2_o21ai_1 _23505_ (.B1(net10759),
    .Y(_05495_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[9] ),
    .A2(net10158));
 sg13g2_and3_1 _23506_ (.X(_05496_),
    .A(net10743),
    .B(_05494_),
    .C(_05495_));
 sg13g2_nor3_1 _23507_ (.A(net10743),
    .B(\u_ac_controller_soc_inst.cbus_wdata[18] ),
    .C(net10158),
    .Y(_05497_));
 sg13g2_o21ai_1 _23508_ (.B1(net11043),
    .Y(_05498_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[10] ),
    .A2(net10241));
 sg13g2_nor3_1 _23509_ (.A(_05496_),
    .B(_05497_),
    .C(_05498_),
    .Y(_00354_));
 sg13g2_buf_2 place9858 (.A(_11123_),
    .X(net9858));
 sg13g2_nand2b_1 _23511_ (.Y(_05500_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[11] ),
    .A_N(net10760));
 sg13g2_o21ai_1 _23512_ (.B1(net10759),
    .Y(_05501_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[10] ),
    .A2(net10158));
 sg13g2_and3_1 _23513_ (.X(_05502_),
    .A(net10746),
    .B(_05500_),
    .C(_05501_));
 sg13g2_buf_2 place9844 (.A(_11204_),
    .X(net9844));
 sg13g2_nor3_1 _23515_ (.A(net10745),
    .B(\u_ac_controller_soc_inst.cbus_wdata[19] ),
    .C(net10154),
    .Y(_05504_));
 sg13g2_o21ai_1 _23516_ (.B1(net11042),
    .Y(_05505_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[11] ),
    .A2(net10239));
 sg13g2_nor3_1 _23517_ (.A(_05502_),
    .B(_05504_),
    .C(_05505_),
    .Y(_00355_));
 sg13g2_nand2b_1 _23518_ (.Y(_05506_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[12] ),
    .A_N(net10760));
 sg13g2_buf_2 place9850 (.A(net9849),
    .X(net9850));
 sg13g2_buf_2 place9849 (.A(_11204_),
    .X(net9849));
 sg13g2_o21ai_1 _23521_ (.B1(net10760),
    .Y(_05509_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[11] ),
    .A2(net10155));
 sg13g2_and3_1 _23522_ (.X(_05510_),
    .A(net10746),
    .B(_05506_),
    .C(_05509_));
 sg13g2_nor3_1 _23523_ (.A(net10746),
    .B(\u_ac_controller_soc_inst.cbus_wdata[20] ),
    .C(net10155),
    .Y(_05511_));
 sg13g2_o21ai_1 _23524_ (.B1(net11042),
    .Y(_05512_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[12] ),
    .A2(net10239));
 sg13g2_nor3_1 _23525_ (.A(_05510_),
    .B(_05511_),
    .C(_05512_),
    .Y(_00356_));
 sg13g2_nand2b_1 _23526_ (.Y(_05513_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[13] ),
    .A_N(net10760));
 sg13g2_buf_2 place9855 (.A(net9854),
    .X(net9855));
 sg13g2_o21ai_1 _23528_ (.B1(net10760),
    .Y(_05515_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[12] ),
    .A2(net10155));
 sg13g2_and3_1 _23529_ (.X(_05516_),
    .A(net10745),
    .B(_05513_),
    .C(_05515_));
 sg13g2_nor3_1 _23530_ (.A(net10745),
    .B(\u_ac_controller_soc_inst.cbus_wdata[21] ),
    .C(net10154),
    .Y(_05517_));
 sg13g2_o21ai_1 _23531_ (.B1(net11042),
    .Y(_05518_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[13] ),
    .A2(net10240));
 sg13g2_nor3_1 _23532_ (.A(_05516_),
    .B(_05517_),
    .C(_05518_),
    .Y(_00357_));
 sg13g2_nand2b_1 _23533_ (.Y(_05519_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[14] ),
    .A_N(net10758));
 sg13g2_o21ai_1 _23534_ (.B1(net10758),
    .Y(_05520_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[13] ),
    .A2(net10154));
 sg13g2_and3_1 _23535_ (.X(_05521_),
    .A(net10745),
    .B(_05519_),
    .C(_05520_));
 sg13g2_nor3_1 _23536_ (.A(net10744),
    .B(\u_ac_controller_soc_inst.cbus_wdata[22] ),
    .C(net10153),
    .Y(_05522_));
 sg13g2_o21ai_1 _23537_ (.B1(net11042),
    .Y(_05523_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[14] ),
    .A2(net10240));
 sg13g2_nor3_1 _23538_ (.A(_05521_),
    .B(_05522_),
    .C(_05523_),
    .Y(_00358_));
 sg13g2_nand2b_1 _23539_ (.Y(_05524_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[15] ),
    .A_N(net10758));
 sg13g2_o21ai_1 _23540_ (.B1(net10758),
    .Y(_05525_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[14] ),
    .A2(net10153));
 sg13g2_and3_1 _23541_ (.X(_05526_),
    .A(net10744),
    .B(_05524_),
    .C(_05525_));
 sg13g2_nor3_1 _23542_ (.A(net10744),
    .B(\u_ac_controller_soc_inst.cbus_wdata[23] ),
    .C(net10153),
    .Y(_05527_));
 sg13g2_o21ai_1 _23543_ (.B1(net11042),
    .Y(_05528_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[15] ),
    .A2(net10240));
 sg13g2_nor3_1 _23544_ (.A(_05526_),
    .B(_05527_),
    .C(_05528_),
    .Y(_00359_));
 sg13g2_nand2b_1 _23545_ (.Y(_05529_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[16] ),
    .A_N(net10757));
 sg13g2_o21ai_1 _23546_ (.B1(net10756),
    .Y(_05530_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[15] ),
    .A2(net10156));
 sg13g2_and3_1 _23547_ (.X(_05531_),
    .A(net10742),
    .B(_05529_),
    .C(_05530_));
 sg13g2_nor3_1 _23548_ (.A(net10742),
    .B(\u_ac_controller_soc_inst.cbus_wdata[8] ),
    .C(net10156),
    .Y(_05532_));
 sg13g2_o21ai_1 _23549_ (.B1(net11043),
    .Y(_05533_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[16] ),
    .A2(net10241));
 sg13g2_nor3_1 _23550_ (.A(_05531_),
    .B(_05532_),
    .C(_05533_),
    .Y(_00360_));
 sg13g2_nand2b_1 _23551_ (.Y(_05534_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[17] ),
    .A_N(net10757));
 sg13g2_o21ai_1 _23552_ (.B1(net10757),
    .Y(_05535_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[16] ),
    .A2(net10156));
 sg13g2_and3_1 _23553_ (.X(_05536_),
    .A(net10743),
    .B(_05534_),
    .C(_05535_));
 sg13g2_buf_2 place9848 (.A(net9847),
    .X(net9848));
 sg13g2_nor3_1 _23555_ (.A(net10743),
    .B(\u_ac_controller_soc_inst.cbus_wdata[9] ),
    .C(net10158),
    .Y(_05538_));
 sg13g2_o21ai_1 _23556_ (.B1(net11043),
    .Y(_05539_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[17] ),
    .A2(net10241));
 sg13g2_nor3_1 _23557_ (.A(_05536_),
    .B(_05538_),
    .C(_05539_),
    .Y(_00361_));
 sg13g2_nand2b_1 _23558_ (.Y(_05540_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[18] ),
    .A_N(net10760));
 sg13g2_o21ai_1 _23559_ (.B1(net10759),
    .Y(_05541_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[17] ),
    .A2(net10158));
 sg13g2_and3_1 _23560_ (.X(_05542_),
    .A(net10746),
    .B(_05540_),
    .C(_05541_));
 sg13g2_nor3_1 _23561_ (.A(net10746),
    .B(\u_ac_controller_soc_inst.cbus_wdata[10] ),
    .C(net10155),
    .Y(_05543_));
 sg13g2_o21ai_1 _23562_ (.B1(net11042),
    .Y(_05544_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[18] ),
    .A2(net10239));
 sg13g2_nor3_1 _23563_ (.A(_05542_),
    .B(_05543_),
    .C(_05544_),
    .Y(_00362_));
 sg13g2_buf_2 place9862 (.A(_11083_),
    .X(net9862));
 sg13g2_nand2b_1 _23565_ (.Y(_05546_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[19] ),
    .A_N(net10760));
 sg13g2_o21ai_1 _23566_ (.B1(net10759),
    .Y(_05547_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[18] ),
    .A2(net10155));
 sg13g2_and3_1 _23567_ (.X(_05548_),
    .A(net10746),
    .B(_05546_),
    .C(_05547_));
 sg13g2_nor3_1 _23568_ (.A(net10746),
    .B(\u_ac_controller_soc_inst.cbus_wdata[11] ),
    .C(net10155),
    .Y(_05549_));
 sg13g2_buf_2 place9865 (.A(net9864),
    .X(net9865));
 sg13g2_buf_2 place9835 (.A(_11284_),
    .X(net9835));
 sg13g2_o21ai_1 _23571_ (.B1(net11042),
    .Y(_05552_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[19] ),
    .A2(net10239));
 sg13g2_nor3_1 _23572_ (.A(_05548_),
    .B(_05549_),
    .C(_05552_),
    .Y(_00363_));
 sg13g2_nand2b_1 _23573_ (.Y(_05553_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[1] ),
    .A_N(net10748));
 sg13g2_o21ai_1 _23574_ (.B1(net10748),
    .Y(_05554_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[0] ),
    .A2(net10149));
 sg13g2_and3_1 _23575_ (.X(_05555_),
    .A(net10735),
    .B(_05553_),
    .C(_05554_));
 sg13g2_nor3_1 _23576_ (.A(net10737),
    .B(\u_ac_controller_soc_inst.cbus_wdata[25] ),
    .C(net10149),
    .Y(_05556_));
 sg13g2_o21ai_1 _23577_ (.B1(net11040),
    .Y(_05557_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[1] ),
    .A2(net10237));
 sg13g2_nor3_1 _23578_ (.A(_05555_),
    .B(_05556_),
    .C(_05557_),
    .Y(_00364_));
 sg13g2_buf_2 place9860 (.A(net9859),
    .X(net9860));
 sg13g2_nand2b_1 _23580_ (.Y(_05559_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[20] ),
    .A_N(net10757));
 sg13g2_o21ai_1 _23581_ (.B1(net10758),
    .Y(_05560_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[19] ),
    .A2(net10154));
 sg13g2_and3_1 _23582_ (.X(_05561_),
    .A(net10743),
    .B(_05559_),
    .C(_05560_));
 sg13g2_buf_2 place9837 (.A(net9836),
    .X(net9837));
 sg13g2_nor3_1 _23584_ (.A(net10743),
    .B(\u_ac_controller_soc_inst.cbus_wdata[12] ),
    .C(net10157),
    .Y(_05563_));
 sg13g2_o21ai_1 _23585_ (.B1(net11043),
    .Y(_05564_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[20] ),
    .A2(net10241));
 sg13g2_nor3_1 _23586_ (.A(_05561_),
    .B(_05563_),
    .C(_05564_),
    .Y(_00365_));
 sg13g2_nand2b_1 _23587_ (.Y(_05565_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[21] ),
    .A_N(net10756));
 sg13g2_buf_2 place9870 (.A(net9868),
    .X(net9870));
 sg13g2_o21ai_1 _23589_ (.B1(net10757),
    .Y(_05567_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[20] ),
    .A2(net10156));
 sg13g2_and3_1 _23590_ (.X(_05568_),
    .A(net10742),
    .B(_05565_),
    .C(_05567_));
 sg13g2_nor3_1 _23591_ (.A(net10742),
    .B(\u_ac_controller_soc_inst.cbus_wdata[13] ),
    .C(net10157),
    .Y(_05569_));
 sg13g2_o21ai_1 _23592_ (.B1(net11044),
    .Y(_05570_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[21] ),
    .A2(net10241));
 sg13g2_nor3_1 _23593_ (.A(_05568_),
    .B(_05569_),
    .C(_05570_),
    .Y(_00366_));
 sg13g2_nand2b_1 _23594_ (.Y(_05571_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[22] ),
    .A_N(net10756));
 sg13g2_buf_2 place9843 (.A(net9840),
    .X(net9843));
 sg13g2_o21ai_1 _23596_ (.B1(net10756),
    .Y(_05573_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[21] ),
    .A2(net10157));
 sg13g2_and3_1 _23597_ (.X(_05574_),
    .A(net10741),
    .B(_05571_),
    .C(_05573_));
 sg13g2_nor3_1 _23598_ (.A(net10741),
    .B(\u_ac_controller_soc_inst.cbus_wdata[14] ),
    .C(net10157),
    .Y(_05575_));
 sg13g2_o21ai_1 _23599_ (.B1(net11043),
    .Y(_05576_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[22] ),
    .A2(net10241));
 sg13g2_nor3_1 _23600_ (.A(_05574_),
    .B(_05575_),
    .C(_05576_),
    .Y(_00367_));
 sg13g2_nand2b_1 _23601_ (.Y(_05577_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[23] ),
    .A_N(net10756));
 sg13g2_o21ai_1 _23602_ (.B1(net10756),
    .Y(_05578_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[22] ),
    .A2(net10157));
 sg13g2_and3_1 _23603_ (.X(_05579_),
    .A(net10741),
    .B(_05577_),
    .C(_05578_));
 sg13g2_nor3_1 _23604_ (.A(net10741),
    .B(\u_ac_controller_soc_inst.cbus_wdata[15] ),
    .C(net10157),
    .Y(_05580_));
 sg13g2_o21ai_1 _23605_ (.B1(net11043),
    .Y(_05581_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[23] ),
    .A2(net10241));
 sg13g2_nor3_1 _23606_ (.A(_05579_),
    .B(_05580_),
    .C(_05581_),
    .Y(_00368_));
 sg13g2_nand2b_1 _23607_ (.Y(_05582_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[24] ),
    .A_N(net10752));
 sg13g2_o21ai_1 _23608_ (.B1(net10752),
    .Y(_05583_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[23] ),
    .A2(net10151));
 sg13g2_and3_1 _23609_ (.X(_05584_),
    .A(net10740),
    .B(_05582_),
    .C(_05583_));
 sg13g2_nor3_1 _23610_ (.A(net10740),
    .B(net10605),
    .C(net10151),
    .Y(_05585_));
 sg13g2_o21ai_1 _23611_ (.B1(net11046),
    .Y(_05586_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[24] ),
    .A2(net10235));
 sg13g2_nor3_1 _23612_ (.A(_05584_),
    .B(_05585_),
    .C(_05586_),
    .Y(_00369_));
 sg13g2_nand2b_1 _23613_ (.Y(_05587_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[25] ),
    .A_N(net10752));
 sg13g2_o21ai_1 _23614_ (.B1(net10752),
    .Y(_05588_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[24] ),
    .A2(net10151));
 sg13g2_and3_1 _23615_ (.X(_05589_),
    .A(net10740),
    .B(_05587_),
    .C(_05588_));
 sg13g2_nor3_1 _23616_ (.A(net10740),
    .B(\u_ac_controller_soc_inst.cbus_wdata[1] ),
    .C(net10152),
    .Y(_05590_));
 sg13g2_o21ai_1 _23617_ (.B1(net11046),
    .Y(_05591_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[25] ),
    .A2(net10238));
 sg13g2_nor3_1 _23618_ (.A(_05589_),
    .B(_05590_),
    .C(_05591_),
    .Y(_00370_));
 sg13g2_nand2b_1 _23619_ (.Y(_05592_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[26] ),
    .A_N(net10753));
 sg13g2_o21ai_1 _23620_ (.B1(net10753),
    .Y(_05593_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[25] ),
    .A2(net10152));
 sg13g2_and3_1 _23621_ (.X(_05594_),
    .A(net10739),
    .B(_05592_),
    .C(_05593_));
 sg13g2_buf_2 place9857 (.A(_11123_),
    .X(net9857));
 sg13g2_nor3_1 _23623_ (.A(net10739),
    .B(\u_ac_controller_soc_inst.cbus_wdata[2] ),
    .C(net10159),
    .Y(_05596_));
 sg13g2_o21ai_1 _23624_ (.B1(net11046),
    .Y(_05597_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[26] ),
    .A2(net10238));
 sg13g2_nor3_1 _23625_ (.A(_05594_),
    .B(_05596_),
    .C(_05597_),
    .Y(_00371_));
 sg13g2_nand2b_1 _23626_ (.Y(_05598_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[27] ),
    .A_N(net10753));
 sg13g2_o21ai_1 _23627_ (.B1(net10753),
    .Y(_05599_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[26] ),
    .A2(net10159));
 sg13g2_and3_1 _23628_ (.X(_05600_),
    .A(net10739),
    .B(_05598_),
    .C(_05599_));
 sg13g2_nor3_1 _23629_ (.A(net10739),
    .B(\u_ac_controller_soc_inst.cbus_wdata[3] ),
    .C(net10159),
    .Y(_05601_));
 sg13g2_o21ai_1 _23630_ (.B1(net11046),
    .Y(_05602_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[27] ),
    .A2(net10238));
 sg13g2_nor3_1 _23631_ (.A(_05600_),
    .B(_05601_),
    .C(_05602_),
    .Y(_00372_));
 sg13g2_buf_2 place9854 (.A(net9853),
    .X(net9854));
 sg13g2_nand2b_1 _23633_ (.Y(_05604_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[28] ),
    .A_N(net10754));
 sg13g2_o21ai_1 _23634_ (.B1(net10754),
    .Y(_05605_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[27] ),
    .A2(net10159));
 sg13g2_and3_1 _23635_ (.X(_05606_),
    .A(net10739),
    .B(_05604_),
    .C(_05605_));
 sg13g2_nor3_1 _23636_ (.A(net10739),
    .B(\u_ac_controller_soc_inst.cbus_wdata[4] ),
    .C(net10159),
    .Y(_05607_));
 sg13g2_buf_2 place9826 (.A(_11364_),
    .X(net9826));
 sg13g2_buf_2 place9859 (.A(net9858),
    .X(net9859));
 sg13g2_o21ai_1 _23639_ (.B1(net11046),
    .Y(_05610_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[28] ),
    .A2(net10238));
 sg13g2_nor3_1 _23640_ (.A(_05606_),
    .B(_05607_),
    .C(_05610_),
    .Y(_00373_));
 sg13g2_nand2b_1 _23641_ (.Y(_05611_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[29] ),
    .A_N(net10754));
 sg13g2_o21ai_1 _23642_ (.B1(net10754),
    .Y(_05612_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[28] ),
    .A2(net10159));
 sg13g2_and3_1 _23643_ (.X(_05613_),
    .A(net10740),
    .B(_05611_),
    .C(_05612_));
 sg13g2_nor3_1 _23644_ (.A(net10740),
    .B(\u_ac_controller_soc_inst.cbus_wdata[5] ),
    .C(net10159),
    .Y(_05614_));
 sg13g2_o21ai_1 _23645_ (.B1(net11046),
    .Y(_05615_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[29] ),
    .A2(net10238));
 sg13g2_nor3_1 _23646_ (.A(_05613_),
    .B(_05614_),
    .C(_05615_),
    .Y(_00374_));
 sg13g2_buf_2 place9836 (.A(net9835),
    .X(net9836));
 sg13g2_nand2b_1 _23648_ (.Y(_05617_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[2] ),
    .A_N(net10750));
 sg13g2_o21ai_1 _23649_ (.B1(net10750),
    .Y(_05618_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[1] ),
    .A2(net10149));
 sg13g2_and3_1 _23650_ (.X(_05619_),
    .A(net10737),
    .B(_05617_),
    .C(_05618_));
 sg13g2_buf_2 place9829 (.A(net9828),
    .X(net9829));
 sg13g2_nor3_1 _23652_ (.A(net10737),
    .B(\u_ac_controller_soc_inst.cbus_wdata[26] ),
    .C(net10149),
    .Y(_05621_));
 sg13g2_o21ai_1 _23653_ (.B1(net11040),
    .Y(_05622_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[2] ),
    .A2(net10237));
 sg13g2_nor3_1 _23654_ (.A(_05619_),
    .B(_05621_),
    .C(_05622_),
    .Y(_00375_));
 sg13g2_nand2b_1 _23655_ (.Y(_05623_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[30] ),
    .A_N(net10754));
 sg13g2_o21ai_1 _23656_ (.B1(net10754),
    .Y(_05624_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[29] ),
    .A2(net10152));
 sg13g2_and3_1 _23657_ (.X(_05625_),
    .A(net10740),
    .B(_05623_),
    .C(_05624_));
 sg13g2_nor3_1 _23658_ (.A(net10740),
    .B(\u_ac_controller_soc_inst.cbus_wdata[6] ),
    .C(net10152),
    .Y(_05626_));
 sg13g2_o21ai_1 _23659_ (.B1(net11046),
    .Y(_05627_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[30] ),
    .A2(net10238));
 sg13g2_nor3_1 _23660_ (.A(_05625_),
    .B(_05626_),
    .C(_05627_),
    .Y(_00376_));
 sg13g2_nand2b_1 _23661_ (.Y(_05628_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[31] ),
    .A_N(net10751));
 sg13g2_o21ai_1 _23662_ (.B1(net10751),
    .Y(_05629_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[30] ),
    .A2(net10151));
 sg13g2_and3_1 _23663_ (.X(_05630_),
    .A(net10738),
    .B(_05628_),
    .C(_05629_));
 sg13g2_nor3_1 _23664_ (.A(net10738),
    .B(\u_ac_controller_soc_inst.cbus_wdata[7] ),
    .C(net10151),
    .Y(_05631_));
 sg13g2_o21ai_1 _23665_ (.B1(net11040),
    .Y(_05632_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[31] ),
    .A2(net10235));
 sg13g2_nor3_1 _23666_ (.A(_05630_),
    .B(_05631_),
    .C(_05632_),
    .Y(_00377_));
 sg13g2_nor2b_2 _23667_ (.A(net10735),
    .B_N(net10234),
    .Y(_05633_));
 sg13g2_buf_2 place9828 (.A(net9826),
    .X(net9828));
 sg13g2_buf_2 place9827 (.A(net9826),
    .X(net9827));
 sg13g2_nand3b_1 _23670_ (.B(net10237),
    .C(net10750),
    .Y(_05636_),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[31] ));
 sg13g2_o21ai_1 _23671_ (.B1(_05636_),
    .Y(_05637_),
    .A1(net10748),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[32] ));
 sg13g2_o21ai_1 _23672_ (.B1(net11039),
    .Y(_05638_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[32] ),
    .A2(net10237));
 sg13g2_a221oi_1 _23673_ (.B2(net10735),
    .C1(_05638_),
    .B1(_05637_),
    .A1(net10459),
    .Y(_00378_),
    .A2(_05633_));
 sg13g2_nand3b_1 _23674_ (.B(net10237),
    .C(net10748),
    .Y(_05639_),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[32] ));
 sg13g2_o21ai_1 _23675_ (.B1(_05639_),
    .Y(_05640_),
    .A1(net10749),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[33] ));
 sg13g2_o21ai_1 _23676_ (.B1(net11039),
    .Y(_05641_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[33] ),
    .A2(net10236));
 sg13g2_a221oi_1 _23677_ (.B2(net10736),
    .C1(_05641_),
    .B1(_05640_),
    .A1(_08126_),
    .Y(_00379_),
    .A2(_05633_));
 sg13g2_nand3_1 _23678_ (.B(_04310_),
    .C(net10236),
    .A(net10749),
    .Y(_05642_));
 sg13g2_o21ai_1 _23679_ (.B1(_05642_),
    .Y(_05643_),
    .A1(net10749),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[36] ));
 sg13g2_o21ai_1 _23680_ (.B1(net11039),
    .Y(_05644_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[36] ),
    .A2(net10237));
 sg13g2_a221oi_1 _23681_ (.B2(net10736),
    .C1(_05644_),
    .B1(_05643_),
    .A1(_07707_),
    .Y(_00382_),
    .A2(_05633_));
 sg13g2_nand3b_1 _23682_ (.B(net10237),
    .C(net10748),
    .Y(_05645_),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[36] ));
 sg13g2_o21ai_1 _23683_ (.B1(_05645_),
    .Y(_05646_),
    .A1(net10749),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[37] ));
 sg13g2_o21ai_1 _23684_ (.B1(net11039),
    .Y(_05647_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[37] ),
    .A2(net10236));
 sg13g2_a221oi_1 _23685_ (.B2(net10735),
    .C1(_05647_),
    .B1(_05646_),
    .A1(_08078_),
    .Y(_00383_),
    .A2(_05633_));
 sg13g2_inv_1 _23686_ (.Y(_05648_),
    .A(net10614));
 sg13g2_nand3b_1 _23687_ (.B(net10236),
    .C(net10747),
    .Y(_05649_),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[37] ));
 sg13g2_o21ai_1 _23688_ (.B1(_05649_),
    .Y(_05650_),
    .A1(net10747),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[38] ));
 sg13g2_o21ai_1 _23689_ (.B1(net11039),
    .Y(_05651_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[38] ),
    .A2(net10236));
 sg13g2_a221oi_1 _23690_ (.B2(net10735),
    .C1(_05651_),
    .B1(_05650_),
    .A1(_05648_),
    .Y(_00384_),
    .A2(_05633_));
 sg13g2_inv_1 _23691_ (.Y(_05652_),
    .A(net10613));
 sg13g2_nand3b_1 _23692_ (.B(net10234),
    .C(net10747),
    .Y(_05653_),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[38] ));
 sg13g2_o21ai_1 _23693_ (.B1(_05653_),
    .Y(_05654_),
    .A1(net10747),
    .A2(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[39] ));
 sg13g2_o21ai_1 _23694_ (.B1(net11038),
    .Y(_05655_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[39] ),
    .A2(net10234));
 sg13g2_a221oi_1 _23695_ (.B2(net10735),
    .C1(_05655_),
    .B1(_05654_),
    .A1(_05652_),
    .Y(_00385_),
    .A2(_05633_));
 sg13g2_nand2b_1 _23696_ (.Y(_05656_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[3] ),
    .A_N(net10750));
 sg13g2_o21ai_1 _23697_ (.B1(net10750),
    .Y(_05657_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[2] ),
    .A2(net10150));
 sg13g2_and3_1 _23698_ (.X(_05658_),
    .A(net10737),
    .B(_05656_),
    .C(_05657_));
 sg13g2_nor3_1 _23699_ (.A(net10737),
    .B(\u_ac_controller_soc_inst.cbus_wdata[27] ),
    .C(net10150),
    .Y(_05659_));
 sg13g2_o21ai_1 _23700_ (.B1(net11040),
    .Y(_05660_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[3] ),
    .A2(net10235));
 sg13g2_nor3_1 _23701_ (.A(_05658_),
    .B(_05659_),
    .C(_05660_),
    .Y(_00386_));
 sg13g2_nand2b_1 _23702_ (.Y(_05661_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[4] ),
    .A_N(net10751));
 sg13g2_o21ai_1 _23703_ (.B1(net10750),
    .Y(_05662_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[3] ),
    .A2(net10150));
 sg13g2_and3_1 _23704_ (.X(_05663_),
    .A(_00103_),
    .B(_05661_),
    .C(_05662_));
 sg13g2_nor3_1 _23705_ (.A(net10737),
    .B(\u_ac_controller_soc_inst.cbus_wdata[28] ),
    .C(net10150),
    .Y(_05664_));
 sg13g2_o21ai_1 _23706_ (.B1(net11040),
    .Y(_05665_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[4] ),
    .A2(net10238));
 sg13g2_nor3_1 _23707_ (.A(_05663_),
    .B(_05664_),
    .C(_05665_),
    .Y(_00387_));
 sg13g2_nand2b_1 _23708_ (.Y(_05666_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[5] ),
    .A_N(net10751));
 sg13g2_o21ai_1 _23709_ (.B1(net10751),
    .Y(_05667_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[4] ),
    .A2(net10150));
 sg13g2_and3_1 _23710_ (.X(_05668_),
    .A(net10738),
    .B(_05666_),
    .C(_05667_));
 sg13g2_nor3_1 _23711_ (.A(net10738),
    .B(\u_ac_controller_soc_inst.cbus_wdata[29] ),
    .C(net10151),
    .Y(_05669_));
 sg13g2_o21ai_1 _23712_ (.B1(net11040),
    .Y(_05670_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[5] ),
    .A2(net10238));
 sg13g2_nor3_1 _23713_ (.A(_05668_),
    .B(_05669_),
    .C(_05670_),
    .Y(_00388_));
 sg13g2_nand2b_1 _23714_ (.Y(_05671_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[6] ),
    .A_N(net10752));
 sg13g2_o21ai_1 _23715_ (.B1(net10751),
    .Y(_05672_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[5] ),
    .A2(net10151));
 sg13g2_and3_1 _23716_ (.X(_05673_),
    .A(net10738),
    .B(_05671_),
    .C(_05672_));
 sg13g2_nor3_1 _23717_ (.A(net10738),
    .B(\u_ac_controller_soc_inst.cbus_wdata[30] ),
    .C(net10151),
    .Y(_05674_));
 sg13g2_o21ai_1 _23718_ (.B1(net11041),
    .Y(_05675_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[6] ),
    .A2(net10235));
 sg13g2_nor3_1 _23719_ (.A(_05673_),
    .B(_05674_),
    .C(_05675_),
    .Y(_00389_));
 sg13g2_nand2b_1 _23720_ (.Y(_05676_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[7] ),
    .A_N(net10755));
 sg13g2_o21ai_1 _23721_ (.B1(net10756),
    .Y(_05677_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[6] ),
    .A2(net10153));
 sg13g2_and3_1 _23722_ (.X(_05678_),
    .A(net10741),
    .B(_05676_),
    .C(_05677_));
 sg13g2_nor3_1 _23723_ (.A(net10738),
    .B(\u_ac_controller_soc_inst.cbus_wdata[31] ),
    .C(net10153),
    .Y(_05679_));
 sg13g2_o21ai_1 _23724_ (.B1(net11041),
    .Y(_05680_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[7] ),
    .A2(net10235));
 sg13g2_nor3_1 _23725_ (.A(_05678_),
    .B(_05679_),
    .C(_05680_),
    .Y(_00390_));
 sg13g2_nand2b_1 _23726_ (.Y(_05681_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[8] ),
    .A_N(net10755));
 sg13g2_o21ai_1 _23727_ (.B1(net10755),
    .Y(_05682_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[7] ),
    .A2(net10153));
 sg13g2_and3_1 _23728_ (.X(_05683_),
    .A(net10744),
    .B(_05681_),
    .C(_05682_));
 sg13g2_nor3_1 _23729_ (.A(net10744),
    .B(\u_ac_controller_soc_inst.cbus_wdata[16] ),
    .C(net10153),
    .Y(_05684_));
 sg13g2_o21ai_1 _23730_ (.B1(net11042),
    .Y(_05685_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[8] ),
    .A2(net10240));
 sg13g2_nor3_1 _23731_ (.A(_05683_),
    .B(_05684_),
    .C(_05685_),
    .Y(_00391_));
 sg13g2_nand2b_1 _23732_ (.Y(_05686_),
    .B(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[9] ),
    .A_N(net10757));
 sg13g2_o21ai_1 _23733_ (.B1(net10758),
    .Y(_05687_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[8] ),
    .A2(net10154));
 sg13g2_and3_1 _23734_ (.X(_05688_),
    .A(net10743),
    .B(_05686_),
    .C(_05687_));
 sg13g2_nor3_1 _23735_ (.A(net10743),
    .B(\u_ac_controller_soc_inst.cbus_wdata[17] ),
    .C(net10158),
    .Y(_05689_));
 sg13g2_o21ai_1 _23736_ (.B1(net11043),
    .Y(_05690_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[9] ),
    .A2(net10241));
 sg13g2_nor3_1 _23737_ (.A(_05688_),
    .B(_05689_),
    .C(_05690_),
    .Y(_00392_));
 sg13g2_nand2_1 _23738_ (.Y(_05691_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[5] ),
    .B(_04325_));
 sg13g2_nor2_1 _23739_ (.A(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[5] ),
    .B(_04325_),
    .Y(_05692_));
 sg13g2_a21oi_1 _23740_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[5] ),
    .A2(_05691_),
    .Y(_05693_),
    .B1(_05692_));
 sg13g2_nand2b_1 _23741_ (.Y(_05694_),
    .B(_00043_),
    .A_N(spi_sensor_cs_n));
 sg13g2_nor4_1 _23742_ (.A(net11004),
    .B(_04327_),
    .C(_05693_),
    .D(_05694_),
    .Y(_00393_));
 sg13g2_nor2b_1 _23743_ (.A(_04316_),
    .B_N(_04331_),
    .Y(_05695_));
 sg13g2_nor3_1 _23744_ (.A(net11004),
    .B(_04317_),
    .C(_05695_),
    .Y(_00395_));
 sg13g2_and3_1 _23745_ (.X(_00396_),
    .A(net11038),
    .B(_05454_),
    .C(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[0] ));
 sg13g2_nor2_1 _23746_ (.A(net10988),
    .B(_05454_),
    .Y(_00398_));
 sg13g2_nand2b_1 _23747_ (.Y(_00397_),
    .B(_00398_),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[0] ));
 sg13g2_nand3_1 _23748_ (.B(_04554_),
    .C(_05432_),
    .A(net10234),
    .Y(_05696_));
 sg13g2_mux2_1 _23749_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[0] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[0] ),
    .S(_05696_),
    .X(_05697_));
 sg13g2_and2_1 _23750_ (.A(net11038),
    .B(_05697_),
    .X(_00399_));
 sg13g2_mux2_1 _23751_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[1] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[1] ),
    .S(_05696_),
    .X(_05698_));
 sg13g2_and2_1 _23752_ (.A(net11038),
    .B(_05698_),
    .X(_00400_));
 sg13g2_xor2_1 _23753_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[1] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[2] ),
    .X(_05699_));
 sg13g2_xnor2_1 _23754_ (.Y(_05700_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[28] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[27] ));
 sg13g2_xnor2_1 _23755_ (.Y(_05701_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[3] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2] ));
 sg13g2_xnor2_1 _23756_ (.Y(_05702_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[6] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[5] ));
 sg13g2_xnor2_1 _23757_ (.Y(_05703_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[27] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[26] ));
 sg13g2_nand4_1 _23758_ (.B(_05701_),
    .C(_05702_),
    .A(_05700_),
    .Y(_05704_),
    .D(_05703_));
 sg13g2_xnor2_1 _23759_ (.Y(_05705_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[11] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[10] ));
 sg13g2_xnor2_1 _23760_ (.Y(_05706_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[17] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[16] ));
 sg13g2_xnor2_1 _23761_ (.Y(_05707_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[21] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[20] ));
 sg13g2_xnor2_1 _23762_ (.Y(_05708_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[24] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[23] ));
 sg13g2_nand4_1 _23763_ (.B(_05706_),
    .C(_05707_),
    .A(_05705_),
    .Y(_05709_),
    .D(_05708_));
 sg13g2_xor2_1 _23764_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[25] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[26] ),
    .X(_05710_));
 sg13g2_xor2_1 _23765_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[24] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[25] ),
    .X(_05711_));
 sg13g2_xor2_1 _23766_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[29] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[30] ),
    .X(_05712_));
 sg13g2_xor2_1 _23767_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[7] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[8] ),
    .X(_05713_));
 sg13g2_nor4_1 _23768_ (.A(_05710_),
    .B(_05711_),
    .C(_05712_),
    .D(_05713_),
    .Y(_05714_));
 sg13g2_xnor2_1 _23769_ (.Y(_05715_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[4] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[3] ));
 sg13g2_xnor2_1 _23770_ (.Y(_05716_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[29] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[28] ));
 sg13g2_nand4_1 _23771_ (.B(_05714_),
    .C(_05715_),
    .A(_04572_),
    .Y(_05717_),
    .D(_05716_));
 sg13g2_nor4_1 _23772_ (.A(_05699_),
    .B(_05704_),
    .C(_05709_),
    .D(_05717_),
    .Y(_05718_));
 sg13g2_xor2_1 _23773_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[8] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[9] ),
    .X(_05719_));
 sg13g2_xor2_1 _23774_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[11] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[12] ),
    .X(_05720_));
 sg13g2_xor2_1 _23775_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[19] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[20] ),
    .X(_05721_));
 sg13g2_xor2_1 _23776_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[15] ),
    .X(_05722_));
 sg13g2_nor4_2 _23777_ (.A(_05719_),
    .B(_05720_),
    .C(_05721_),
    .Y(_05723_),
    .D(_05722_));
 sg13g2_xnor2_1 _23778_ (.Y(_05724_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[5] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[4] ));
 sg13g2_nand4_1 _23779_ (.B(_05718_),
    .C(_05723_),
    .A(_04498_),
    .Y(_05725_),
    .D(_05724_));
 sg13g2_xnor2_1 _23780_ (.Y(_05726_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[23] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22] ));
 sg13g2_xnor2_1 _23781_ (.Y(_05727_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[1] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[0] ));
 sg13g2_xnor2_1 _23782_ (.Y(_05728_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[13] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[12] ));
 sg13g2_nand3_1 _23783_ (.B(_05727_),
    .C(_05728_),
    .A(_05726_),
    .Y(_05729_));
 sg13g2_xnor2_1 _23784_ (.Y(_05730_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[22] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[21] ));
 sg13g2_xnor2_1 _23785_ (.Y(_05731_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[18] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[17] ));
 sg13g2_xnor2_1 _23786_ (.Y(_05732_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[14] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13] ));
 sg13g2_xnor2_1 _23787_ (.Y(_05733_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[16] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[15] ));
 sg13g2_nand4_1 _23788_ (.B(_05731_),
    .C(_05732_),
    .A(_05730_),
    .Y(_05734_),
    .D(_05733_));
 sg13g2_xnor2_1 _23789_ (.Y(_05735_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[7] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[6] ));
 sg13g2_xnor2_1 _23790_ (.Y(_05736_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[19] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[18] ));
 sg13g2_xnor2_1 _23791_ (.Y(_05737_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[31] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[30] ));
 sg13g2_xnor2_1 _23792_ (.Y(_05738_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[10] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9] ));
 sg13g2_nand4_1 _23793_ (.B(_05736_),
    .C(_05737_),
    .A(_05735_),
    .Y(_05739_),
    .D(_05738_));
 sg13g2_nor4_2 _23794_ (.A(_05725_),
    .B(_05729_),
    .C(_05734_),
    .Y(_05740_),
    .D(_05739_));
 sg13g2_nor3_2 _23795_ (.A(net10734),
    .B(net10733),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2] ),
    .Y(_05741_));
 sg13g2_nand3_1 _23796_ (.B(_05740_),
    .C(_05741_),
    .A(_00137_),
    .Y(_05742_));
 sg13g2_and4_2 _23797_ (.A(_07899_),
    .B(_07895_),
    .C(_07902_),
    .D(_04554_),
    .X(_05743_));
 sg13g2_buf_2 place9825 (.A(net9824),
    .X(net9825));
 sg13g2_nor2b_2 _23799_ (.A(_05743_),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync ),
    .Y(_05745_));
 sg13g2_buf_2 place9824 (.A(net9823),
    .X(net9824));
 sg13g2_and2_1 _23801_ (.A(_05740_),
    .B(_05745_),
    .X(_05747_));
 sg13g2_a22oi_1 _23802_ (.Y(_05748_),
    .B1(_05747_),
    .B2(_05741_),
    .A2(_05742_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[0] ));
 sg13g2_nor2_1 _23803_ (.A(net10980),
    .B(_05748_),
    .Y(_00436_));
 sg13g2_and2_1 _23804_ (.A(_04573_),
    .B(_05740_),
    .X(_05749_));
 sg13g2_buf_2 place9823 (.A(_04811_),
    .X(net9823));
 sg13g2_nand2_1 _23806_ (.Y(_05751_),
    .A(_04592_),
    .B(_05749_));
 sg13g2_nor2_2 _23807_ (.A(_00137_),
    .B(_05741_),
    .Y(_05752_));
 sg13g2_nand2_1 _23808_ (.Y(_05753_),
    .A(_05745_),
    .B(_05752_));
 sg13g2_nor2b_2 _23809_ (.A(net10734),
    .B_N(net10733),
    .Y(_05754_));
 sg13g2_buf_2 place9839 (.A(net9838),
    .X(net9839));
 sg13g2_nor2_1 _23811_ (.A(_04592_),
    .B(_05754_),
    .Y(_05756_));
 sg13g2_nor2_1 _23812_ (.A(_05753_),
    .B(_05756_),
    .Y(_05757_));
 sg13g2_a22oi_1 _23813_ (.Y(_05758_),
    .B1(_05757_),
    .B2(_05749_),
    .A2(_05751_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[1] ));
 sg13g2_nor2_1 _23814_ (.A(net10980),
    .B(_05758_),
    .Y(_00437_));
 sg13g2_nand3_1 _23815_ (.B(_05749_),
    .C(_05754_),
    .A(_05745_),
    .Y(_05759_));
 sg13g2_inv_1 _23816_ (.Y(_05760_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[2] ));
 sg13g2_a21o_1 _23817_ (.A2(_05754_),
    .A1(_05749_),
    .B1(_05760_),
    .X(_05761_));
 sg13g2_a21oi_1 _23818_ (.A1(_05759_),
    .A2(_05761_),
    .Y(_00438_),
    .B1(net10980));
 sg13g2_and2_1 _23819_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2] ),
    .B(_05740_),
    .X(_05762_));
 sg13g2_buf_16 clkbuf_leaf_380_clk (.X(clknet_leaf_380_clk),
    .A(clknet_8_120_0_clk));
 sg13g2_inv_1 _23821_ (.Y(_05764_),
    .A(_05762_));
 sg13g2_nor3_1 _23822_ (.A(net10733),
    .B(_05753_),
    .C(_05764_),
    .Y(_05765_));
 sg13g2_o21ai_1 _23823_ (.B1(_04574_),
    .Y(_05766_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[3] ),
    .A2(_05765_));
 sg13g2_inv_2 _23824_ (.Y(_05767_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[3] ));
 sg13g2_a21oi_1 _23825_ (.A1(net10733),
    .A2(_05749_),
    .Y(_05768_),
    .B1(_05767_));
 sg13g2_nand4_1 _23826_ (.B(_05745_),
    .C(_05749_),
    .A(_04595_),
    .Y(_05769_),
    .D(_05752_));
 sg13g2_nor2b_1 _23827_ (.A(_05768_),
    .B_N(_05769_),
    .Y(_05770_));
 sg13g2_a21oi_1 _23828_ (.A1(_05766_),
    .A2(_05770_),
    .Y(_00439_),
    .B1(net10979));
 sg13g2_nor2_2 _23829_ (.A(net10734),
    .B(net10733),
    .Y(_05771_));
 sg13g2_nand3_1 _23830_ (.B(_05745_),
    .C(_05762_),
    .A(_05771_),
    .Y(_05772_));
 sg13g2_inv_1 _23831_ (.Y(_05773_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[4] ));
 sg13g2_a21o_1 _23832_ (.A2(_05762_),
    .A1(_05771_),
    .B1(_05773_),
    .X(_05774_));
 sg13g2_a21oi_1 _23833_ (.A1(_05772_),
    .A2(_05774_),
    .Y(_00440_),
    .B1(net10980));
 sg13g2_buf_2 place9831 (.A(net9830),
    .X(net9831));
 sg13g2_buf_2 place9814 (.A(net9813),
    .X(net9814));
 sg13g2_nand2_1 _23836_ (.Y(_05777_),
    .A(_04592_),
    .B(_05762_));
 sg13g2_a22oi_1 _23837_ (.Y(_05778_),
    .B1(_05777_),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[5] ),
    .A2(_05762_),
    .A1(_05757_));
 sg13g2_nor2_1 _23838_ (.A(net10980),
    .B(_05778_),
    .Y(_00441_));
 sg13g2_nand2_1 _23839_ (.Y(_05779_),
    .A(_05754_),
    .B(_05762_));
 sg13g2_xnor2_1 _23840_ (.Y(_05780_),
    .A(_04573_),
    .B(_05771_));
 sg13g2_and3_2 _23841_ (.X(_05781_),
    .A(_05740_),
    .B(_05745_),
    .C(_05780_));
 sg13g2_a22oi_1 _23842_ (.Y(_05782_),
    .B1(_05781_),
    .B2(_05754_),
    .A2(_05779_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[6] ));
 sg13g2_nor2_1 _23843_ (.A(net10980),
    .B(_05782_),
    .Y(_00442_));
 sg13g2_nand2_1 _23844_ (.Y(_05783_),
    .A(_04595_),
    .B(_05762_));
 sg13g2_a22oi_1 _23845_ (.Y(_05784_),
    .B1(_05783_),
    .B2(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[7] ),
    .A2(_05781_),
    .A1(_05752_));
 sg13g2_buf_2 place9820 (.A(net9819),
    .X(net9820));
 sg13g2_o21ai_1 _23847_ (.B1(net11039),
    .Y(_05786_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[7] ),
    .A2(_05756_));
 sg13g2_nor2_1 _23848_ (.A(_05784_),
    .B(_05786_),
    .Y(_00443_));
 sg13g2_inv_1 _23849_ (.Y(_05787_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[8] ));
 sg13g2_nor2_1 _23850_ (.A(net10987),
    .B(_05787_),
    .Y(_00444_));
 sg13g2_nand2b_1 _23851_ (.Y(_00445_),
    .B(net11055),
    .A_N(ser_rx));
 sg13g2_nand2b_1 _23852_ (.Y(_00446_),
    .B(net11055),
    .A_N(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync1 ));
 sg13g2_inv_1 _23853_ (.Y(_05788_),
    .A(_04563_));
 sg13g2_and3_2 _23854_ (.X(_05789_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_done ),
    .B(_07927_),
    .C(_05788_));
 sg13g2_buf_2 place9817 (.A(net9816),
    .X(net9817));
 sg13g2_buf_16 clkbuf_leaf_391_clk (.X(clknet_leaf_391_clk),
    .A(clknet_8_109_0_clk));
 sg13g2_buf_16 clkbuf_leaf_389_clk (.X(clknet_leaf_389_clk),
    .A(clknet_8_105_0_clk));
 sg13g2_inv_1 _23858_ (.Y(_05793_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[0] ));
 sg13g2_nand3_1 _23859_ (.B(_05793_),
    .C(net9987),
    .A(net10310),
    .Y(_05794_));
 sg13g2_o21ai_1 _23860_ (.B1(_05794_),
    .Y(_05795_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[0] ),
    .A2(_05789_));
 sg13g2_nor2_1 _23861_ (.A(net10986),
    .B(_05795_),
    .Y(_00450_));
 sg13g2_inv_1 _23862_ (.Y(_05796_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[1] ));
 sg13g2_nand3_1 _23863_ (.B(_05796_),
    .C(net9988),
    .A(net10310),
    .Y(_05797_));
 sg13g2_o21ai_1 _23864_ (.B1(_05797_),
    .Y(_05798_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[1] ),
    .A2(net9988));
 sg13g2_nor2_1 _23865_ (.A(net10986),
    .B(_05798_),
    .Y(_00451_));
 sg13g2_nand3_1 _23866_ (.B(_05760_),
    .C(net9987),
    .A(net10310),
    .Y(_05799_));
 sg13g2_o21ai_1 _23867_ (.B1(_05799_),
    .Y(_05800_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[2] ),
    .A2(_05789_));
 sg13g2_nor2_1 _23868_ (.A(net10986),
    .B(_05800_),
    .Y(_00452_));
 sg13g2_nand3_1 _23869_ (.B(_05767_),
    .C(net9987),
    .A(net10310),
    .Y(_05801_));
 sg13g2_o21ai_1 _23870_ (.B1(_05801_),
    .Y(_05802_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[3] ),
    .A2(net9987));
 sg13g2_nor2_1 _23871_ (.A(net10986),
    .B(_05802_),
    .Y(_00453_));
 sg13g2_nand3_1 _23872_ (.B(_05773_),
    .C(net9988),
    .A(net10310),
    .Y(_05803_));
 sg13g2_o21ai_1 _23873_ (.B1(_05803_),
    .Y(_05804_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[4] ),
    .A2(net9988));
 sg13g2_nor2_1 _23874_ (.A(net10979),
    .B(_05804_),
    .Y(_00454_));
 sg13g2_inv_1 _23875_ (.Y(_05805_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[5] ));
 sg13g2_nand3_1 _23876_ (.B(_05805_),
    .C(net9988),
    .A(net10310),
    .Y(_05806_));
 sg13g2_o21ai_1 _23877_ (.B1(_05806_),
    .Y(_05807_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[5] ),
    .A2(net9988));
 sg13g2_nor2_1 _23878_ (.A(net10986),
    .B(_05807_),
    .Y(_00455_));
 sg13g2_inv_1 _23879_ (.Y(_05808_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[6] ));
 sg13g2_nand3_1 _23880_ (.B(_05808_),
    .C(net9988),
    .A(net10310),
    .Y(_05809_));
 sg13g2_o21ai_1 _23881_ (.B1(_05809_),
    .Y(_05810_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[6] ),
    .A2(net9988));
 sg13g2_nor2_1 _23882_ (.A(net10989),
    .B(_05810_),
    .Y(_00456_));
 sg13g2_buf_16 clkbuf_leaf_386_clk (.X(clknet_leaf_386_clk),
    .A(clknet_8_110_0_clk));
 sg13g2_inv_1 _23884_ (.Y(_05812_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[7] ));
 sg13g2_nand3_1 _23885_ (.B(_05812_),
    .C(net9987),
    .A(net10310),
    .Y(_05813_));
 sg13g2_o21ai_1 _23886_ (.B1(_05813_),
    .Y(_05814_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[7] ),
    .A2(net9987));
 sg13g2_nor2_1 _23887_ (.A(net10986),
    .B(_05814_),
    .Y(_00457_));
 sg13g2_nand3_1 _23888_ (.B(_05787_),
    .C(_05789_),
    .A(_04546_),
    .Y(_05815_));
 sg13g2_o21ai_1 _23889_ (.B1(_05815_),
    .Y(_05816_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[8] ),
    .A2(_05789_));
 sg13g2_nor2_1 _23890_ (.A(net10987),
    .B(_05816_),
    .Y(_00458_));
 sg13g2_and2_1 _23891_ (.A(\u_ac_controller_soc_inst.cbus_addr[3] ),
    .B(_04560_),
    .X(_05817_));
 sg13g2_nand2_1 _23892_ (.Y(_05818_),
    .A(_04550_),
    .B(_05817_));
 sg13g2_nor2_1 _23893_ (.A(_08410_),
    .B(_04563_),
    .Y(_05819_));
 sg13g2_o21ai_1 _23894_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_done ),
    .Y(_05820_),
    .A1(_04558_),
    .A2(_05819_));
 sg13g2_o21ai_1 _23895_ (.B1(_05820_),
    .Y(_05821_),
    .A1(_04556_),
    .A2(_05818_));
 sg13g2_and2_1 _23896_ (.A(net11038),
    .B(_05821_),
    .X(_00459_));
 sg13g2_nor2_1 _23897_ (.A(net10615),
    .B(net10617),
    .Y(_05822_));
 sg13g2_nand2_1 _23898_ (.Y(_05823_),
    .A(_07927_),
    .B(_04554_));
 sg13g2_nor3_1 _23899_ (.A(net10606),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_ready ),
    .C(_05823_),
    .Y(_05824_));
 sg13g2_nand4_1 _23900_ (.B(_05822_),
    .C(_04550_),
    .A(\u_ac_controller_soc_inst.cbus_addr[3] ),
    .Y(_05825_),
    .D(_05824_));
 sg13g2_buf_2 place9830 (.A(_11364_),
    .X(net9830));
 sg13g2_o21ai_1 _23902_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[0] ),
    .Y(_05827_),
    .A1(net10621),
    .A2(_05825_));
 sg13g2_nor2_1 _23903_ (.A(net10621),
    .B(_05825_),
    .Y(_05828_));
 sg13g2_nand3_1 _23904_ (.B(_07927_),
    .C(_05828_),
    .A(net10605),
    .Y(_05829_));
 sg13g2_a21oi_1 _23905_ (.A1(_05827_),
    .A2(_05829_),
    .Y(_00460_),
    .B1(net10976));
 sg13g2_o21ai_1 _23906_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[1] ),
    .Y(_05830_),
    .A1(net10621),
    .A2(_05825_));
 sg13g2_nand3_1 _23907_ (.B(_07927_),
    .C(_05828_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[1] ),
    .Y(_05831_));
 sg13g2_a21oi_1 _23908_ (.A1(_05830_),
    .A2(_05831_),
    .Y(_00461_),
    .B1(net10976));
 sg13g2_o21ai_1 _23909_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[2] ),
    .Y(_05832_),
    .A1(net10621),
    .A2(_05825_));
 sg13g2_nand3_1 _23910_ (.B(_07927_),
    .C(_05828_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[2] ),
    .Y(_05833_));
 sg13g2_buf_2 place9806 (.A(_07936_),
    .X(net9806));
 sg13g2_buf_16 clkbuf_leaf_385_clk (.X(clknet_leaf_385_clk),
    .A(clknet_8_111_0_clk));
 sg13g2_a21oi_1 _23913_ (.A1(_05832_),
    .A2(_05833_),
    .Y(_00462_),
    .B1(net10976));
 sg13g2_nand4_1 _23914_ (.B(_04550_),
    .C(_05743_),
    .A(net10621),
    .Y(_05836_),
    .D(_05817_));
 sg13g2_buf_2 place9813 (.A(net9812),
    .X(net9813));
 sg13g2_buf_16 clkbuf_leaf_384_clk (.X(clknet_leaf_384_clk),
    .A(clknet_8_122_0_clk));
 sg13g2_mux2_1 _23917_ (.A0(net10605),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[0] ),
    .S(net10147),
    .X(_05839_));
 sg13g2_and2_1 _23918_ (.A(net11047),
    .B(_05839_),
    .X(_00463_));
 sg13g2_inv_2 _23919_ (.Y(_05840_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[10] ));
 sg13g2_nand2_1 _23920_ (.Y(_05841_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[10] ),
    .B(net10148));
 sg13g2_o21ai_1 _23921_ (.B1(_05841_),
    .Y(_05842_),
    .A1(_05840_),
    .A2(net10148));
 sg13g2_and2_1 _23922_ (.A(net11044),
    .B(_05842_),
    .X(_00464_));
 sg13g2_inv_2 _23923_ (.Y(_05843_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[11] ));
 sg13g2_nand2_1 _23924_ (.Y(_05844_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[11] ),
    .B(net10148));
 sg13g2_o21ai_1 _23925_ (.B1(_05844_),
    .Y(_05845_),
    .A1(_05843_),
    .A2(net10148));
 sg13g2_and2_1 _23926_ (.A(net11044),
    .B(_05845_),
    .X(_00465_));
 sg13g2_mux2_1 _23927_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[12] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[12] ),
    .S(net10145),
    .X(_05846_));
 sg13g2_and2_1 _23928_ (.A(net11045),
    .B(_05846_),
    .X(_00466_));
 sg13g2_buf_16 clkbuf_leaf_382_clk (.X(clknet_leaf_382_clk),
    .A(clknet_8_123_0_clk));
 sg13g2_mux2_1 _23930_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[13] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[13] ),
    .S(net10145),
    .X(_05848_));
 sg13g2_and2_1 _23931_ (.A(net11045),
    .B(_05848_),
    .X(_00467_));
 sg13g2_mux2_1 _23932_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[14] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[14] ),
    .S(net10145),
    .X(_05849_));
 sg13g2_and2_1 _23933_ (.A(net11045),
    .B(_05849_),
    .X(_00468_));
 sg13g2_mux2_1 _23934_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[15] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[15] ),
    .S(net10145),
    .X(_05850_));
 sg13g2_and2_1 _23935_ (.A(net11045),
    .B(_05850_),
    .X(_00469_));
 sg13g2_mux2_1 _23936_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[16] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[16] ),
    .S(net10146),
    .X(_05851_));
 sg13g2_and2_1 _23937_ (.A(net11045),
    .B(_05851_),
    .X(_00470_));
 sg13g2_buf_2 place9812 (.A(_04974_),
    .X(net9812));
 sg13g2_mux2_1 _23939_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[17] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[17] ),
    .S(net10146),
    .X(_05853_));
 sg13g2_and2_1 _23940_ (.A(net11057),
    .B(_05853_),
    .X(_00471_));
 sg13g2_mux2_1 _23941_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[18] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[18] ),
    .S(net10146),
    .X(_05854_));
 sg13g2_and2_1 _23942_ (.A(net11057),
    .B(_05854_),
    .X(_00472_));
 sg13g2_mux2_1 _23943_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[19] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[19] ),
    .S(net10146),
    .X(_05855_));
 sg13g2_and2_1 _23944_ (.A(net11057),
    .B(_05855_),
    .X(_00473_));
 sg13g2_mux2_1 _23945_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[1] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[1] ),
    .S(net10147),
    .X(_05856_));
 sg13g2_and2_1 _23946_ (.A(net11047),
    .B(_05856_),
    .X(_00474_));
 sg13g2_mux2_1 _23947_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[20] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[20] ),
    .S(net10146),
    .X(_05857_));
 sg13g2_and2_1 _23948_ (.A(net11057),
    .B(_05857_),
    .X(_00475_));
 sg13g2_mux2_1 _23949_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[21] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[21] ),
    .S(net10146),
    .X(_05858_));
 sg13g2_and2_1 _23950_ (.A(net11057),
    .B(_05858_),
    .X(_00476_));
 sg13g2_buf_16 clkbuf_leaf_388_clk (.X(clknet_leaf_388_clk),
    .A(clknet_8_110_0_clk));
 sg13g2_mux2_1 _23952_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[22] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[22] ),
    .S(net10146),
    .X(_05860_));
 sg13g2_and2_1 _23953_ (.A(net11045),
    .B(_05860_),
    .X(_00477_));
 sg13g2_mux2_1 _23954_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[23] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[23] ),
    .S(net10145),
    .X(_05861_));
 sg13g2_and2_1 _23955_ (.A(net11045),
    .B(_05861_),
    .X(_00478_));
 sg13g2_mux2_1 _23956_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[24] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[24] ),
    .S(net10144),
    .X(_05862_));
 sg13g2_and2_1 _23957_ (.A(net11056),
    .B(_05862_),
    .X(_00479_));
 sg13g2_mux2_1 _23958_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[25] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[25] ),
    .S(net10144),
    .X(_05863_));
 sg13g2_and2_1 _23959_ (.A(net11056),
    .B(_05863_),
    .X(_00480_));
 sg13g2_buf_16 clkbuf_leaf_387_clk (.X(clknet_leaf_387_clk),
    .A(clknet_8_111_0_clk));
 sg13g2_mux2_1 _23961_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[26] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[26] ),
    .S(net10144),
    .X(_05865_));
 sg13g2_and2_1 _23962_ (.A(net11056),
    .B(_05865_),
    .X(_00481_));
 sg13g2_mux2_1 _23963_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[27] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[27] ),
    .S(net10144),
    .X(_05866_));
 sg13g2_and2_1 _23964_ (.A(net11056),
    .B(_05866_),
    .X(_00482_));
 sg13g2_mux2_1 _23965_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[28] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[28] ),
    .S(net10144),
    .X(_05867_));
 sg13g2_and2_1 _23966_ (.A(net11057),
    .B(_05867_),
    .X(_00483_));
 sg13g2_mux2_1 _23967_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[29] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[29] ),
    .S(net10144),
    .X(_05868_));
 sg13g2_and2_1 _23968_ (.A(net11057),
    .B(_05868_),
    .X(_00484_));
 sg13g2_mux2_1 _23969_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[2] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[2] ),
    .S(net10147),
    .X(_05869_));
 sg13g2_and2_1 _23970_ (.A(net11047),
    .B(_05869_),
    .X(_00485_));
 sg13g2_mux2_1 _23971_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[30] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[30] ),
    .S(net10144),
    .X(_05870_));
 sg13g2_and2_1 _23972_ (.A(net11057),
    .B(_05870_),
    .X(_00486_));
 sg13g2_buf_16 clkbuf_leaf_394_clk (.X(clknet_leaf_394_clk),
    .A(clknet_8_108_0_clk));
 sg13g2_mux2_1 _23974_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[31] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[31] ),
    .S(net10145),
    .X(_05872_));
 sg13g2_and2_1 _23975_ (.A(net11047),
    .B(_05872_),
    .X(_00487_));
 sg13g2_mux2_1 _23976_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[3] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[3] ),
    .S(net10147),
    .X(_05873_));
 sg13g2_and2_1 _23977_ (.A(net11047),
    .B(_05873_),
    .X(_00488_));
 sg13g2_mux2_1 _23978_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[4] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[4] ),
    .S(net10144),
    .X(_05874_));
 sg13g2_and2_1 _23979_ (.A(net11047),
    .B(_05874_),
    .X(_00489_));
 sg13g2_mux2_1 _23980_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[5] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[5] ),
    .S(net10147),
    .X(_05875_));
 sg13g2_and2_1 _23981_ (.A(net11047),
    .B(_05875_),
    .X(_00490_));
 sg13g2_mux2_1 _23982_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[6] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[6] ),
    .S(net10147),
    .X(_05876_));
 sg13g2_and2_1 _23983_ (.A(net11045),
    .B(_05876_),
    .X(_00491_));
 sg13g2_mux2_1 _23984_ (.A0(\u_ac_controller_soc_inst.cbus_wdata[7] ),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[7] ),
    .S(net10147),
    .X(_05877_));
 sg13g2_and2_1 _23985_ (.A(net11047),
    .B(_05877_),
    .X(_00492_));
 sg13g2_inv_2 _23986_ (.Y(_05878_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[8] ));
 sg13g2_nand2_1 _23987_ (.Y(_05879_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[8] ),
    .B(net10148));
 sg13g2_o21ai_1 _23988_ (.B1(_05879_),
    .Y(_05880_),
    .A1(_05878_),
    .A2(net10148));
 sg13g2_and2_1 _23989_ (.A(net11044),
    .B(_05880_),
    .X(_00493_));
 sg13g2_inv_2 _23990_ (.Y(_05881_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[9] ));
 sg13g2_nand2_1 _23991_ (.Y(_05882_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[9] ),
    .B(net10148));
 sg13g2_o21ai_1 _23992_ (.B1(_05882_),
    .Y(_05883_),
    .A1(_05881_),
    .A2(net10148));
 sg13g2_and2_1 _23993_ (.A(net11044),
    .B(_05883_),
    .X(_00494_));
 sg13g2_nor2_1 _23994_ (.A(_04460_),
    .B(_04703_),
    .Y(_05884_));
 sg13g2_nand2_1 _23995_ (.Y(_05885_),
    .A(_04566_),
    .B(_05884_));
 sg13g2_a21oi_1 _23996_ (.A1(_04548_),
    .A2(_05885_),
    .Y(_00495_),
    .B1(_08213_));
 sg13g2_a21oi_2 _23997_ (.B1(_05743_),
    .Y(_05886_),
    .A2(_00111_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout ));
 sg13g2_buf_16 clkbuf_leaf_393_clk (.X(clknet_leaf_393_clk),
    .A(clknet_8_109_0_clk));
 sg13g2_inv_4 _23999_ (.A(_05886_),
    .Y(_05888_));
 sg13g2_inv_1 _24000_ (.Y(_05889_),
    .A(_00111_));
 sg13g2_nor4_1 _24001_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[0] ),
    .C(_05889_),
    .D(_05743_),
    .Y(_05890_));
 sg13g2_a21oi_1 _24002_ (.A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[0] ),
    .A2(_05888_),
    .Y(_05891_),
    .B1(_05890_));
 sg13g2_nor2_1 _24003_ (.A(net11012),
    .B(_05891_),
    .Y(_00497_));
 sg13g2_a21oi_1 _24004_ (.A1(_04546_),
    .A2(_04737_),
    .Y(_05892_),
    .B1(_05889_));
 sg13g2_o21ai_1 _24005_ (.B1(net11049),
    .Y(_05893_),
    .A1(_05743_),
    .A2(_05892_));
 sg13g2_buf_2 place9822 (.A(net9821),
    .X(net9822));
 sg13g2_buf_2 place9808 (.A(net9807),
    .X(net9808));
 sg13g2_nor2_2 _24008_ (.A(_04729_),
    .B(_05888_),
    .Y(_05896_));
 sg13g2_and4_1 _24009_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[9] ),
    .B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[8] ),
    .C(_04720_),
    .D(_05896_),
    .X(_05897_));
 sg13g2_xnor2_1 _24010_ (.Y(_05898_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[10] ),
    .B(_05897_));
 sg13g2_nor2_1 _24011_ (.A(net9730),
    .B(_05898_),
    .Y(_00498_));
 sg13g2_nand2b_2 _24012_ (.Y(_05899_),
    .B(_05886_),
    .A_N(_04729_));
 sg13g2_nor2_2 _24013_ (.A(_04722_),
    .B(_05899_),
    .Y(_05900_));
 sg13g2_xnor2_1 _24014_ (.Y(_05901_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[11] ),
    .B(_05900_));
 sg13g2_nor2_1 _24015_ (.A(net9732),
    .B(_05901_),
    .Y(_00499_));
 sg13g2_nand2_1 _24016_ (.Y(_05902_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[11] ),
    .B(_05900_));
 sg13g2_xor2_1 _24017_ (.B(_05902_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[12] ),
    .X(_05903_));
 sg13g2_nor2_1 _24018_ (.A(net9732),
    .B(_05903_),
    .Y(_00500_));
 sg13g2_nand3_1 _24019_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[11] ),
    .C(_05900_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[12] ),
    .Y(_05904_));
 sg13g2_xor2_1 _24020_ (.B(_05904_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[13] ),
    .X(_05905_));
 sg13g2_nor2_1 _24021_ (.A(_05893_),
    .B(_05905_),
    .Y(_00501_));
 sg13g2_nand2_2 _24022_ (.Y(_05906_),
    .A(_04732_),
    .B(_05886_));
 sg13g2_xor2_1 _24023_ (.B(_05906_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[14] ),
    .X(_05907_));
 sg13g2_nor2_1 _24024_ (.A(net9732),
    .B(_05907_),
    .Y(_00502_));
 sg13g2_nor2_2 _24025_ (.A(_04733_),
    .B(_05888_),
    .Y(_05908_));
 sg13g2_buf_2 place9809 (.A(net9806),
    .X(net9809));
 sg13g2_nand2_1 _24027_ (.Y(_05910_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[14] ),
    .B(_05908_));
 sg13g2_xor2_1 _24028_ (.B(_05910_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[15] ),
    .X(_05911_));
 sg13g2_nor2_1 _24029_ (.A(net9732),
    .B(_05911_),
    .Y(_00503_));
 sg13g2_nand3_1 _24030_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[14] ),
    .C(_05908_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[15] ),
    .Y(_05912_));
 sg13g2_xor2_1 _24031_ (.B(_05912_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[16] ),
    .X(_05913_));
 sg13g2_nor2_1 _24032_ (.A(net9732),
    .B(_05913_),
    .Y(_00504_));
 sg13g2_nand4_1 _24033_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[15] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[14] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[16] ),
    .Y(_05914_),
    .D(_05908_));
 sg13g2_xor2_1 _24034_ (.B(_05914_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[17] ),
    .X(_05915_));
 sg13g2_nor2_1 _24035_ (.A(net9732),
    .B(_05915_),
    .Y(_00505_));
 sg13g2_nor2_1 _24036_ (.A(_04709_),
    .B(_05906_),
    .Y(_05916_));
 sg13g2_xnor2_1 _24037_ (.Y(_05917_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[18] ),
    .B(_05916_));
 sg13g2_nor2_1 _24038_ (.A(net9732),
    .B(_05917_),
    .Y(_00506_));
 sg13g2_nand2_1 _24039_ (.Y(_05918_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[18] ),
    .B(_05916_));
 sg13g2_xor2_1 _24040_ (.B(_05918_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[19] ),
    .X(_05919_));
 sg13g2_nor2_1 _24041_ (.A(net9732),
    .B(_05919_),
    .Y(_00507_));
 sg13g2_buf_2 place10940 (.A(net10939),
    .X(net10940));
 sg13g2_nand2_2 _24043_ (.Y(_05921_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[0] ),
    .B(_05886_));
 sg13g2_xor2_1 _24044_ (.B(_05921_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[1] ),
    .X(_05922_));
 sg13g2_nor2_1 _24045_ (.A(net9730),
    .B(_05922_),
    .Y(_00508_));
 sg13g2_nand2_1 _24046_ (.Y(_05923_),
    .A(_04711_),
    .B(_05908_));
 sg13g2_xor2_1 _24047_ (.B(_05923_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[20] ),
    .X(_05924_));
 sg13g2_nor2_1 _24048_ (.A(net9733),
    .B(_05924_),
    .Y(_00509_));
 sg13g2_nand3_1 _24049_ (.B(_04711_),
    .C(_05908_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[20] ),
    .Y(_05925_));
 sg13g2_xor2_1 _24050_ (.B(_05925_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[21] ),
    .X(_05926_));
 sg13g2_nor2_1 _24051_ (.A(net9733),
    .B(_05926_),
    .Y(_00510_));
 sg13g2_nand2_1 _24052_ (.Y(_05927_),
    .A(_04712_),
    .B(_05908_));
 sg13g2_xor2_1 _24053_ (.B(_05927_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[22] ),
    .X(_05928_));
 sg13g2_nor2_1 _24054_ (.A(net9733),
    .B(_05928_),
    .Y(_00511_));
 sg13g2_and3_2 _24055_ (.X(_05929_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[22] ),
    .B(_04712_),
    .C(_05908_));
 sg13g2_buf_2 place9821 (.A(_04811_),
    .X(net9821));
 sg13g2_xnor2_1 _24057_ (.Y(_05931_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[23] ),
    .B(_05929_));
 sg13g2_nor2_1 _24058_ (.A(net9733),
    .B(_05931_),
    .Y(_00512_));
 sg13g2_nand2_1 _24059_ (.Y(_05932_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[23] ),
    .B(_05929_));
 sg13g2_xor2_1 _24060_ (.B(_05932_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[24] ),
    .X(_05933_));
 sg13g2_nor2_1 _24061_ (.A(net9733),
    .B(_05933_),
    .Y(_00513_));
 sg13g2_nand3_1 _24062_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[23] ),
    .C(_05929_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[24] ),
    .Y(_05934_));
 sg13g2_xor2_1 _24063_ (.B(_05934_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[25] ),
    .X(_05935_));
 sg13g2_nor2_1 _24064_ (.A(net9733),
    .B(_05935_),
    .Y(_00514_));
 sg13g2_nand4_1 _24065_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[24] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[23] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[25] ),
    .Y(_05936_),
    .D(_05929_));
 sg13g2_xor2_1 _24066_ (.B(_05936_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[26] ),
    .X(_05937_));
 sg13g2_nor2_1 _24067_ (.A(net9733),
    .B(_05937_),
    .Y(_00515_));
 sg13g2_and2_1 _24068_ (.A(_04717_),
    .B(_05929_),
    .X(_05938_));
 sg13g2_xnor2_1 _24069_ (.Y(_05939_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[27] ),
    .B(_05938_));
 sg13g2_nor2_1 _24070_ (.A(net9733),
    .B(_05939_),
    .Y(_00516_));
 sg13g2_nor2_2 _24071_ (.A(_04718_),
    .B(_05906_),
    .Y(_05940_));
 sg13g2_xnor2_1 _24072_ (.Y(_05941_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[28] ),
    .B(_05940_));
 sg13g2_nor2_1 _24073_ (.A(net9731),
    .B(_05941_),
    .Y(_00517_));
 sg13g2_buf_2 place9863 (.A(net9862),
    .X(net9863));
 sg13g2_nand2_1 _24075_ (.Y(_05943_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[28] ),
    .B(_05940_));
 sg13g2_xor2_1 _24076_ (.B(_05943_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[29] ),
    .X(_05944_));
 sg13g2_nor2_1 _24077_ (.A(_05893_),
    .B(_05944_),
    .Y(_00518_));
 sg13g2_nand3_1 _24078_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[0] ),
    .C(_05886_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[1] ),
    .Y(_05945_));
 sg13g2_xor2_1 _24079_ (.B(_05945_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[2] ),
    .X(_05946_));
 sg13g2_nor2_1 _24080_ (.A(net9731),
    .B(_05946_),
    .Y(_00519_));
 sg13g2_nand3_1 _24081_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[28] ),
    .C(_05940_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[29] ),
    .Y(_05947_));
 sg13g2_xor2_1 _24082_ (.B(_05947_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[30] ),
    .X(_05948_));
 sg13g2_nor2_1 _24083_ (.A(net9731),
    .B(_05948_),
    .Y(_00520_));
 sg13g2_inv_1 _24084_ (.Y(_05949_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[31] ));
 sg13g2_nand4_1 _24085_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[29] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[28] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[30] ),
    .Y(_05950_),
    .D(_05940_));
 sg13g2_a21oi_1 _24086_ (.A1(_05949_),
    .A2(_05950_),
    .Y(_00521_),
    .B1(net9731));
 sg13g2_nand4_1 _24087_ (.B(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[1] ),
    .C(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[0] ),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[2] ),
    .Y(_05951_),
    .D(_05886_));
 sg13g2_xor2_1 _24088_ (.B(_05951_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[3] ),
    .X(_05952_));
 sg13g2_nor2_1 _24089_ (.A(net9731),
    .B(_05952_),
    .Y(_00522_));
 sg13g2_o21ai_1 _24090_ (.B1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[4] ),
    .Y(_05953_),
    .A1(_04724_),
    .A2(_05921_));
 sg13g2_or3_1 _24091_ (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[4] ),
    .B(_04724_),
    .C(_05921_),
    .X(_05954_));
 sg13g2_a21oi_1 _24092_ (.A1(_05953_),
    .A2(_05954_),
    .Y(_00523_),
    .B1(net9730));
 sg13g2_nand2_1 _24093_ (.Y(_05955_),
    .A(_04728_),
    .B(_05886_));
 sg13g2_xor2_1 _24094_ (.B(_05955_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[5] ),
    .X(_05956_));
 sg13g2_nor2_1 _24095_ (.A(net9730),
    .B(_05956_),
    .Y(_00524_));
 sg13g2_xor2_1 _24096_ (.B(_05899_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[6] ),
    .X(_05957_));
 sg13g2_nor2_1 _24097_ (.A(net9730),
    .B(_05957_),
    .Y(_00525_));
 sg13g2_nand2_1 _24098_ (.Y(_05958_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[6] ),
    .B(_05896_));
 sg13g2_xor2_1 _24099_ (.B(_05958_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[7] ),
    .X(_05959_));
 sg13g2_nor2_1 _24100_ (.A(net9730),
    .B(_05959_),
    .Y(_00526_));
 sg13g2_nand2_1 _24101_ (.Y(_05960_),
    .A(_04720_),
    .B(_05896_));
 sg13g2_xor2_1 _24102_ (.B(_05960_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[8] ),
    .X(_05961_));
 sg13g2_nor2_1 _24103_ (.A(net9730),
    .B(_05961_),
    .Y(_00527_));
 sg13g2_nand3_1 _24104_ (.B(_04720_),
    .C(_05896_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[8] ),
    .Y(_05962_));
 sg13g2_xor2_1 _24105_ (.B(_05962_),
    .A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[9] ),
    .X(_05963_));
 sg13g2_nor2_1 _24106_ (.A(net9730),
    .B(_05963_),
    .Y(_00528_));
 sg13g2_o21ai_1 _24107_ (.B1(_05885_),
    .Y(_05964_),
    .A1(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfering ),
    .A2(_04689_));
 sg13g2_a21oi_1 _24108_ (.A1(_04548_),
    .A2(_05964_),
    .Y(_00529_),
    .B1(_08213_));
 sg13g2_and2_1 _24109_ (.A(net11048),
    .B(_00140_),
    .X(_00530_));
 sg13g2_inv_2 _24110_ (.Y(_05965_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[10] ));
 sg13g2_and4_2 _24111_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[0] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[1] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[2] ),
    .D(\u_ac_controller_soc_inst.u_picorv32.count_cycle[3] ),
    .X(_05966_));
 sg13g2_buf_2 place9818 (.A(net9816),
    .X(net9818));
 sg13g2_and3_2 _24113_ (.X(_05968_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[4] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[5] ),
    .C(_05966_));
 sg13g2_buf_2 place9805 (.A(_08417_),
    .X(net9805));
 sg13g2_and3_1 _24115_ (.X(_05970_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[6] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[7] ),
    .C(_05968_));
 sg13g2_nand3_1 _24116_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[9] ),
    .C(_05970_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[8] ),
    .Y(_05971_));
 sg13g2_xnor2_1 _24117_ (.Y(_05972_),
    .A(_05965_),
    .B(_05971_));
 sg13g2_nor2_1 _24118_ (.A(net11015),
    .B(_05972_),
    .Y(_00531_));
 sg13g2_nor2_2 _24119_ (.A(_05965_),
    .B(_05971_),
    .Y(_05973_));
 sg13g2_xnor2_1 _24120_ (.Y(_05974_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[11] ),
    .B(_05973_));
 sg13g2_nor2_1 _24121_ (.A(net11015),
    .B(_05974_),
    .Y(_00532_));
 sg13g2_nand2_1 _24122_ (.Y(_05975_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[11] ),
    .B(_05973_));
 sg13g2_xor2_1 _24123_ (.B(_05975_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[12] ),
    .X(_05976_));
 sg13g2_nor2_1 _24124_ (.A(net11015),
    .B(_05976_),
    .Y(_00533_));
 sg13g2_inv_2 _24125_ (.Y(_05977_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[8] ));
 sg13g2_and2_1 _24126_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[6] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[7] ),
    .X(_05978_));
 sg13g2_nand4_1 _24127_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[5] ),
    .C(_05966_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[4] ),
    .Y(_05979_),
    .D(_05978_));
 sg13g2_buf_2 place9807 (.A(net9806),
    .X(net9807));
 sg13g2_nand2_1 _24129_ (.Y(_05981_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[9] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[10] ));
 sg13g2_nand2_1 _24130_ (.Y(_05982_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[11] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[12] ));
 sg13g2_nor4_2 _24131_ (.A(_05977_),
    .B(_05979_),
    .C(_05981_),
    .Y(_05983_),
    .D(_05982_));
 sg13g2_xnor2_1 _24132_ (.Y(_05984_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[13] ),
    .B(_05983_));
 sg13g2_nor2_1 _24133_ (.A(net11015),
    .B(_05984_),
    .Y(_00534_));
 sg13g2_and4_2 _24134_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[11] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[12] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[13] ),
    .D(_05973_),
    .X(_05985_));
 sg13g2_buf_16 clkbuf_leaf_395_clk (.X(clknet_leaf_395_clk),
    .A(clknet_8_100_0_clk));
 sg13g2_xnor2_1 _24136_ (.Y(_05987_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[14] ),
    .B(_05985_));
 sg13g2_nor2_1 _24137_ (.A(net11027),
    .B(_05987_),
    .Y(_00535_));
 sg13g2_nand2_1 _24138_ (.Y(_05988_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[14] ),
    .B(_05985_));
 sg13g2_xor2_1 _24139_ (.B(_05988_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[15] ),
    .X(_05989_));
 sg13g2_nor2_1 _24140_ (.A(net11026),
    .B(_05989_),
    .Y(_00536_));
 sg13g2_and2_1 _24141_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[14] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[15] ),
    .X(_05990_));
 sg13g2_nand3_1 _24142_ (.B(_05983_),
    .C(_05990_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[13] ),
    .Y(_05991_));
 sg13g2_xor2_1 _24143_ (.B(_05991_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[16] ),
    .X(_05992_));
 sg13g2_nor2_1 _24144_ (.A(net11026),
    .B(_05992_),
    .Y(_00537_));
 sg13g2_buf_2 place9816 (.A(_04971_),
    .X(net9816));
 sg13g2_and4_2 _24146_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[13] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[16] ),
    .C(_05983_),
    .D(_05990_),
    .X(_05994_));
 sg13g2_xnor2_1 _24147_ (.Y(_05995_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[17] ),
    .B(_05994_));
 sg13g2_nor2_1 _24148_ (.A(net11020),
    .B(_05995_),
    .Y(_00538_));
 sg13g2_inv_1 _24149_ (.Y(_05996_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[17] ));
 sg13g2_nand4_1 _24150_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[15] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[16] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[14] ),
    .Y(_05997_),
    .D(_05985_));
 sg13g2_nor2_1 _24151_ (.A(_05996_),
    .B(_05997_),
    .Y(_05998_));
 sg13g2_xnor2_1 _24152_ (.Y(_05999_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[18] ),
    .B(_05998_));
 sg13g2_nor2_1 _24153_ (.A(net11022),
    .B(_05999_),
    .Y(_00539_));
 sg13g2_nand2_1 _24154_ (.Y(_06000_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[18] ),
    .B(_05998_));
 sg13g2_xor2_1 _24155_ (.B(_06000_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[19] ),
    .X(_06001_));
 sg13g2_nor2_1 _24156_ (.A(net11022),
    .B(_06001_),
    .Y(_00540_));
 sg13g2_xnor2_1 _24157_ (.Y(_06002_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[0] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[1] ));
 sg13g2_nor2_1 _24158_ (.A(net11009),
    .B(_06002_),
    .Y(_00541_));
 sg13g2_inv_2 _24159_ (.Y(_06003_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[20] ));
 sg13g2_nand4_1 _24160_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[18] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[19] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[17] ),
    .Y(_06004_),
    .D(_05994_));
 sg13g2_buf_2 place9802 (.A(net9801),
    .X(net9802));
 sg13g2_xnor2_1 _24162_ (.Y(_06006_),
    .A(_06003_),
    .B(_06004_));
 sg13g2_nor2_1 _24163_ (.A(net11023),
    .B(_06006_),
    .Y(_00542_));
 sg13g2_nor2_1 _24164_ (.A(_06003_),
    .B(_06004_),
    .Y(_06007_));
 sg13g2_xnor2_1 _24165_ (.Y(_06008_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[21] ),
    .B(_06007_));
 sg13g2_nor2_1 _24166_ (.A(net11022),
    .B(_06008_),
    .Y(_00543_));
 sg13g2_nand2_1 _24167_ (.Y(_06009_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[21] ),
    .B(_06007_));
 sg13g2_xor2_1 _24168_ (.B(_06009_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[22] ),
    .X(_06010_));
 sg13g2_nor2_1 _24169_ (.A(net11022),
    .B(_06010_),
    .Y(_00544_));
 sg13g2_nand2_2 _24170_ (.Y(_06011_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[21] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[22] ));
 sg13g2_nor3_2 _24171_ (.A(_06003_),
    .B(_06004_),
    .C(_06011_),
    .Y(_06012_));
 sg13g2_xnor2_1 _24172_ (.Y(_06013_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[23] ),
    .B(_06012_));
 sg13g2_nor2_1 _24173_ (.A(net11023),
    .B(_06013_),
    .Y(_00545_));
 sg13g2_nand2_1 _24174_ (.Y(_06014_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[23] ),
    .B(_06012_));
 sg13g2_xor2_1 _24175_ (.B(_06014_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[24] ),
    .X(_06015_));
 sg13g2_nor2_1 _24176_ (.A(net11023),
    .B(_06015_),
    .Y(_00546_));
 sg13g2_nand3_1 _24177_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[24] ),
    .C(_06012_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[23] ),
    .Y(_06016_));
 sg13g2_xnor2_1 _24178_ (.Y(_06017_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[25] ),
    .B(_06016_));
 sg13g2_and2_1 _24179_ (.A(net11055),
    .B(_06017_),
    .X(_00547_));
 sg13g2_inv_1 _24180_ (.Y(_06018_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[25] ));
 sg13g2_nor2_1 _24181_ (.A(_06018_),
    .B(_06016_),
    .Y(_06019_));
 sg13g2_xnor2_1 _24182_ (.Y(_06020_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[26] ),
    .B(_06019_));
 sg13g2_nor2_1 _24183_ (.A(net11023),
    .B(_06020_),
    .Y(_00548_));
 sg13g2_buf_2 place9819 (.A(net9818),
    .X(net9819));
 sg13g2_nand2_1 _24185_ (.Y(_06022_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[26] ),
    .B(_06019_));
 sg13g2_xor2_1 _24186_ (.B(_06022_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[27] ),
    .X(_06023_));
 sg13g2_nor2_1 _24187_ (.A(net11023),
    .B(_06023_),
    .Y(_00549_));
 sg13g2_and2_1 _24188_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[25] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[26] ),
    .X(_06024_));
 sg13g2_nand4_1 _24189_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[24] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[27] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[23] ),
    .Y(_06025_),
    .D(_06024_));
 sg13g2_nor4_2 _24190_ (.A(_06003_),
    .B(_06004_),
    .C(_06011_),
    .Y(_06026_),
    .D(_06025_));
 sg13g2_xnor2_1 _24191_ (.Y(_06027_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[28] ),
    .B(_06026_));
 sg13g2_nor2_1 _24192_ (.A(net11023),
    .B(_06027_),
    .Y(_00550_));
 sg13g2_nand2_1 _24193_ (.Y(_06028_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[28] ),
    .B(_06026_));
 sg13g2_xor2_1 _24194_ (.B(_06028_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[29] ),
    .X(_06029_));
 sg13g2_nor2_1 _24195_ (.A(net11022),
    .B(_06029_),
    .Y(_00551_));
 sg13g2_nand2_1 _24196_ (.Y(_06030_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[0] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[1] ));
 sg13g2_xor2_1 _24197_ (.B(_06030_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[2] ),
    .X(_06031_));
 sg13g2_nor2_1 _24198_ (.A(net11009),
    .B(_06031_),
    .Y(_00552_));
 sg13g2_and3_1 _24199_ (.X(_06032_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[28] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[29] ),
    .C(_06026_));
 sg13g2_xnor2_1 _24200_ (.Y(_06033_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[30] ),
    .B(_06032_));
 sg13g2_nor2_1 _24201_ (.A(net11020),
    .B(_06033_),
    .Y(_00553_));
 sg13g2_nand4_1 _24202_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[29] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[30] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[28] ),
    .Y(_06034_),
    .D(_06026_));
 sg13g2_buf_2 place9846 (.A(net9845),
    .X(net9846));
 sg13g2_xor2_1 _24204_ (.B(_06034_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[31] ),
    .X(_06036_));
 sg13g2_nor2_1 _24205_ (.A(net11026),
    .B(_06036_),
    .Y(_00554_));
 sg13g2_and2_1 _24206_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[30] ),
    .B(_06032_),
    .X(_06037_));
 sg13g2_nand2_2 _24207_ (.Y(_06038_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[31] ),
    .B(_06037_));
 sg13g2_buf_2 place9800 (.A(net9799),
    .X(net9800));
 sg13g2_xor2_1 _24209_ (.B(_06038_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[32] ),
    .X(_06040_));
 sg13g2_nor2_1 _24210_ (.A(net11015),
    .B(_06040_),
    .Y(_00555_));
 sg13g2_and3_1 _24211_ (.X(_06041_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[32] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[31] ),
    .C(_06037_));
 sg13g2_xnor2_1 _24212_ (.Y(_06042_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[33] ),
    .B(_06041_));
 sg13g2_nor2_1 _24213_ (.A(net11015),
    .B(_06042_),
    .Y(_00556_));
 sg13g2_nand2_2 _24214_ (.Y(_06043_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[32] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[33] ));
 sg13g2_nor2_2 _24215_ (.A(_06038_),
    .B(_06043_),
    .Y(_06044_));
 sg13g2_xnor2_1 _24216_ (.Y(_06045_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[34] ),
    .B(_06044_));
 sg13g2_nor2_1 _24217_ (.A(net11012),
    .B(_06045_),
    .Y(_00557_));
 sg13g2_buf_2 place9845 (.A(net9844),
    .X(net9845));
 sg13g2_nand2_1 _24219_ (.Y(_06047_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[34] ),
    .B(_06044_));
 sg13g2_xnor2_1 _24220_ (.Y(_06048_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[35] ),
    .B(_06047_));
 sg13g2_and2_1 _24221_ (.A(net11048),
    .B(_06048_),
    .X(_00558_));
 sg13g2_and3_2 _24222_ (.X(_06049_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[34] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[35] ),
    .C(_06044_));
 sg13g2_buf_2 place9840 (.A(_11284_),
    .X(net9840));
 sg13g2_xnor2_1 _24224_ (.Y(_06051_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[36] ),
    .B(_06049_));
 sg13g2_nor2_1 _24225_ (.A(net11012),
    .B(_06051_),
    .Y(_00559_));
 sg13g2_nand2_1 _24226_ (.Y(_06052_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[36] ),
    .B(_06049_));
 sg13g2_xnor2_1 _24227_ (.Y(_06053_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[37] ),
    .B(_06052_));
 sg13g2_and2_1 _24228_ (.A(net11049),
    .B(_06053_),
    .X(_00560_));
 sg13g2_and2_1 _24229_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[36] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[37] ),
    .X(_06054_));
 sg13g2_nand2_1 _24230_ (.Y(_06055_),
    .A(_06049_),
    .B(_06054_));
 sg13g2_xnor2_1 _24231_ (.Y(_06056_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[38] ),
    .B(_06055_));
 sg13g2_and2_1 _24232_ (.A(net11049),
    .B(_06056_),
    .X(_00561_));
 sg13g2_buf_2 place9801 (.A(net9800),
    .X(net9801));
 sg13g2_nand4_1 _24234_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[35] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[38] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[34] ),
    .Y(_06058_),
    .D(_06054_));
 sg13g2_nor3_2 _24235_ (.A(_06038_),
    .B(_06043_),
    .C(_06058_),
    .Y(_06059_));
 sg13g2_xnor2_1 _24236_ (.Y(_06060_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[39] ),
    .B(_06059_));
 sg13g2_nor2_1 _24237_ (.A(net11010),
    .B(_06060_),
    .Y(_00562_));
 sg13g2_nand3_1 _24238_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[1] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[2] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[0] ),
    .Y(_06061_));
 sg13g2_xor2_1 _24239_ (.B(_06061_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[3] ),
    .X(_06062_));
 sg13g2_nor2_1 _24240_ (.A(net11012),
    .B(_06062_),
    .Y(_00563_));
 sg13g2_nand2_1 _24241_ (.Y(_06063_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[39] ),
    .B(_06059_));
 sg13g2_xor2_1 _24242_ (.B(_06063_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[40] ),
    .X(_06064_));
 sg13g2_nor2_1 _24243_ (.A(net11010),
    .B(_06064_),
    .Y(_00564_));
 sg13g2_nand3_1 _24244_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[40] ),
    .C(_06059_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[39] ),
    .Y(_06065_));
 sg13g2_xor2_1 _24245_ (.B(_06065_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[41] ),
    .X(_06066_));
 sg13g2_nor2_1 _24246_ (.A(net11010),
    .B(_06066_),
    .Y(_00565_));
 sg13g2_nand3_1 _24247_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[40] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[41] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[39] ),
    .Y(_06067_));
 sg13g2_or3_1 _24248_ (.A(_06043_),
    .B(_06058_),
    .C(_06067_),
    .X(_06068_));
 sg13g2_buf_2 place9803 (.A(net9802),
    .X(net9803));
 sg13g2_nor2_2 _24250_ (.A(_06038_),
    .B(_06068_),
    .Y(_06070_));
 sg13g2_xnor2_1 _24251_ (.Y(_06071_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[42] ),
    .B(_06070_));
 sg13g2_nor2_1 _24252_ (.A(net11016),
    .B(_06071_),
    .Y(_00566_));
 sg13g2_nand2_1 _24253_ (.Y(_06072_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[42] ),
    .B(_06070_));
 sg13g2_xnor2_1 _24254_ (.Y(_06073_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[43] ),
    .B(_06072_));
 sg13g2_and2_1 _24255_ (.A(net11049),
    .B(_06073_),
    .X(_00567_));
 sg13g2_nand3_1 _24256_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[43] ),
    .C(_06070_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[42] ),
    .Y(_06074_));
 sg13g2_xnor2_1 _24257_ (.Y(_06075_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[44] ),
    .B(_06074_));
 sg13g2_and2_1 _24258_ (.A(net11049),
    .B(_06075_),
    .X(_00568_));
 sg13g2_nand3_1 _24259_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[43] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[44] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[42] ),
    .Y(_06076_));
 sg13g2_nor3_1 _24260_ (.A(_06038_),
    .B(_06068_),
    .C(_06076_),
    .Y(_06077_));
 sg13g2_xnor2_1 _24261_ (.Y(_06078_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[45] ),
    .B(_06077_));
 sg13g2_nor2_1 _24262_ (.A(net11016),
    .B(_06078_),
    .Y(_00569_));
 sg13g2_nand2_1 _24263_ (.Y(_06079_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[45] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[31] ));
 sg13g2_or3_1 _24264_ (.A(_06068_),
    .B(_06076_),
    .C(_06079_),
    .X(_06080_));
 sg13g2_nor2_1 _24265_ (.A(_06034_),
    .B(_06080_),
    .Y(_06081_));
 sg13g2_xnor2_1 _24266_ (.Y(_06082_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[46] ),
    .B(_06081_));
 sg13g2_nor2_1 _24267_ (.A(net11026),
    .B(_06082_),
    .Y(_00570_));
 sg13g2_nand2_1 _24268_ (.Y(_06083_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[46] ),
    .B(_06081_));
 sg13g2_xor2_1 _24269_ (.B(_06083_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[47] ),
    .X(_06084_));
 sg13g2_nor2_1 _24270_ (.A(net11027),
    .B(_06084_),
    .Y(_00571_));
 sg13g2_inv_2 _24271_ (.Y(_06085_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[48] ));
 sg13g2_nand2_1 _24272_ (.Y(_06086_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[46] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[47] ));
 sg13g2_or2_1 _24273_ (.X(_06087_),
    .B(_06086_),
    .A(_06080_));
 sg13g2_or2_1 _24274_ (.X(_06088_),
    .B(_06087_),
    .A(_06034_));
 sg13g2_xnor2_1 _24275_ (.Y(_06089_),
    .A(_06085_),
    .B(_06088_));
 sg13g2_nor2_1 _24276_ (.A(net11026),
    .B(_06089_),
    .Y(_00572_));
 sg13g2_nor2_1 _24277_ (.A(_06085_),
    .B(_06088_),
    .Y(_06090_));
 sg13g2_xnor2_1 _24278_ (.Y(_06091_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[49] ),
    .B(_06090_));
 sg13g2_nor2_1 _24279_ (.A(net11020),
    .B(_06091_),
    .Y(_00573_));
 sg13g2_buf_16 clkbuf_leaf_396_clk (.X(clknet_leaf_396_clk),
    .A(clknet_8_100_0_clk));
 sg13g2_xnor2_1 _24281_ (.Y(_06093_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[4] ),
    .B(_05966_));
 sg13g2_nor2_1 _24282_ (.A(net11009),
    .B(_06093_),
    .Y(_00574_));
 sg13g2_and2_1 _24283_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[49] ),
    .B(_06090_),
    .X(_06094_));
 sg13g2_buf_2 place9815 (.A(_04974_),
    .X(net9815));
 sg13g2_xnor2_1 _24285_ (.Y(_06096_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[50] ),
    .B(_06094_));
 sg13g2_nor2_1 _24286_ (.A(net11021),
    .B(_06096_),
    .Y(_00575_));
 sg13g2_nand2_1 _24287_ (.Y(_06097_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[50] ),
    .B(_06094_));
 sg13g2_xor2_1 _24288_ (.B(_06097_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[51] ),
    .X(_06098_));
 sg13g2_nor2_1 _24289_ (.A(net11021),
    .B(_06098_),
    .Y(_00576_));
 sg13g2_and2_1 _24290_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[50] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[51] ),
    .X(_06099_));
 sg13g2_buf_2 place10329 (.A(net10326),
    .X(net10329));
 sg13g2_nand2_1 _24292_ (.Y(_06101_),
    .A(_06094_),
    .B(_06099_));
 sg13g2_xor2_1 _24293_ (.B(_06101_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[52] ),
    .X(_06102_));
 sg13g2_nor2_1 _24294_ (.A(net11020),
    .B(_06102_),
    .Y(_00577_));
 sg13g2_nand3_1 _24295_ (.B(_06094_),
    .C(_06099_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[52] ),
    .Y(_06103_));
 sg13g2_xor2_1 _24296_ (.B(_06103_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[53] ),
    .X(_06104_));
 sg13g2_nor2_1 _24297_ (.A(net11020),
    .B(_06104_),
    .Y(_00578_));
 sg13g2_inv_1 _24298_ (.Y(_06105_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[54] ));
 sg13g2_nand4_1 _24299_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[52] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[53] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[49] ),
    .Y(_06106_),
    .D(_06099_));
 sg13g2_or4_1 _24300_ (.A(_06085_),
    .B(_06034_),
    .C(_06087_),
    .D(_06106_),
    .X(_06107_));
 sg13g2_buf_2 place9799 (.A(_09885_),
    .X(net9799));
 sg13g2_xnor2_1 _24302_ (.Y(_06109_),
    .A(_06105_),
    .B(_06107_));
 sg13g2_nor2_1 _24303_ (.A(net11024),
    .B(_06109_),
    .Y(_00579_));
 sg13g2_nor2_1 _24304_ (.A(_06105_),
    .B(_06107_),
    .Y(_06110_));
 sg13g2_xnor2_1 _24305_ (.Y(_06111_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[55] ),
    .B(_06110_));
 sg13g2_nor2_1 _24306_ (.A(net11024),
    .B(_06111_),
    .Y(_00580_));
 sg13g2_nand2_1 _24307_ (.Y(_06112_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[54] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[55] ));
 sg13g2_nor2_1 _24308_ (.A(_06107_),
    .B(_06112_),
    .Y(_06113_));
 sg13g2_xnor2_1 _24309_ (.Y(_06114_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[56] ),
    .B(_06113_));
 sg13g2_nor2_1 _24310_ (.A(net11024),
    .B(_06114_),
    .Y(_00581_));
 sg13g2_inv_1 _24311_ (.Y(_06115_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[56] ));
 sg13g2_nor3_1 _24312_ (.A(_06115_),
    .B(_06107_),
    .C(_06112_),
    .Y(_06116_));
 sg13g2_xnor2_1 _24313_ (.Y(_06117_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[57] ),
    .B(_06116_));
 sg13g2_nor2_1 _24314_ (.A(net11024),
    .B(_06117_),
    .Y(_00582_));
 sg13g2_nand4_1 _24315_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[55] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_cycle[56] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[54] ),
    .Y(_06118_),
    .D(\u_ac_controller_soc_inst.u_picorv32.count_cycle[57] ));
 sg13g2_nor2_1 _24316_ (.A(_06107_),
    .B(_06118_),
    .Y(_06119_));
 sg13g2_xnor2_1 _24317_ (.Y(_06120_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[58] ),
    .B(_06119_));
 sg13g2_nor2_1 _24318_ (.A(net11024),
    .B(_06120_),
    .Y(_00583_));
 sg13g2_buf_2 place9841 (.A(net9840),
    .X(net9841));
 sg13g2_inv_1 _24320_ (.Y(_06122_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[58] ));
 sg13g2_nor3_2 _24321_ (.A(_06122_),
    .B(_06107_),
    .C(_06118_),
    .Y(_06123_));
 sg13g2_xnor2_1 _24322_ (.Y(_06124_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[59] ),
    .B(_06123_));
 sg13g2_nor2_1 _24323_ (.A(net11021),
    .B(_06124_),
    .Y(_00584_));
 sg13g2_nand2_1 _24324_ (.Y(_06125_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[4] ),
    .B(_05966_));
 sg13g2_xor2_1 _24325_ (.B(_06125_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[5] ),
    .X(_06126_));
 sg13g2_nor2_1 _24326_ (.A(net11010),
    .B(_06126_),
    .Y(_00585_));
 sg13g2_nand2_1 _24327_ (.Y(_06127_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[59] ),
    .B(_06123_));
 sg13g2_xor2_1 _24328_ (.B(_06127_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[60] ),
    .X(_06128_));
 sg13g2_nor2_1 _24329_ (.A(net11021),
    .B(_06128_),
    .Y(_00586_));
 sg13g2_and3_2 _24330_ (.X(_06129_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[59] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[60] ),
    .C(_06123_));
 sg13g2_xnor2_1 _24331_ (.Y(_06130_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[61] ),
    .B(_06129_));
 sg13g2_nor2_1 _24332_ (.A(net11029),
    .B(_06130_),
    .Y(_00587_));
 sg13g2_and2_1 _24333_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[61] ),
    .B(_06129_),
    .X(_06131_));
 sg13g2_xnor2_1 _24334_ (.Y(_06132_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[62] ),
    .B(_06131_));
 sg13g2_nor2_1 _24335_ (.A(net11029),
    .B(_06132_),
    .Y(_00588_));
 sg13g2_nand2_1 _24336_ (.Y(_06133_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[62] ),
    .B(_06131_));
 sg13g2_xnor2_1 _24337_ (.Y(_06134_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[63] ),
    .B(_06133_));
 sg13g2_and2_1 _24338_ (.A(net11053),
    .B(_06134_),
    .X(_00589_));
 sg13g2_xnor2_1 _24339_ (.Y(_06135_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[6] ),
    .B(_05968_));
 sg13g2_nor2_1 _24340_ (.A(net11009),
    .B(_06135_),
    .Y(_00590_));
 sg13g2_nand2_1 _24341_ (.Y(_06136_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[6] ),
    .B(_05968_));
 sg13g2_xor2_1 _24342_ (.B(_06136_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_cycle[7] ),
    .X(_06137_));
 sg13g2_nor2_1 _24343_ (.A(net11009),
    .B(_06137_),
    .Y(_00591_));
 sg13g2_xnor2_1 _24344_ (.Y(_06138_),
    .A(_05977_),
    .B(_05979_));
 sg13g2_nor2_1 _24345_ (.A(net11010),
    .B(_06138_),
    .Y(_00592_));
 sg13g2_o21ai_1 _24346_ (.B1(\u_ac_controller_soc_inst.u_picorv32.count_cycle[9] ),
    .Y(_06139_),
    .A1(_05977_),
    .A2(_05979_));
 sg13g2_or3_1 _24347_ (.A(_05977_),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_cycle[9] ),
    .C(_05979_),
    .X(_06140_));
 sg13g2_a21oi_1 _24348_ (.A1(_06139_),
    .A2(_06140_),
    .Y(_00593_),
    .B1(net11010));
 sg13g2_buf_2 place9842 (.A(net9840),
    .X(net9842));
 sg13g2_buf_2 place10330 (.A(net10326),
    .X(net10330));
 sg13g2_buf_2 place9838 (.A(net9835),
    .X(net9838));
 sg13g2_nand3_1 _24352_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoder_trigger ),
    .C(_00141_),
    .A(net10715),
    .Y(_06144_));
 sg13g2_nand2_2 _24353_ (.Y(_06145_),
    .A(net10715),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoder_trigger ));
 sg13g2_nand2_1 _24354_ (.Y(_06146_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[0] ),
    .B(_06145_));
 sg13g2_a21oi_1 _24355_ (.A1(_06144_),
    .A2(_06146_),
    .Y(_00594_),
    .B1(net11022));
 sg13g2_and4_2 _24356_ (.A(\u_ac_controller_soc_inst.u_picorv32.cpu_state[1] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoder_trigger ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[0] ),
    .D(\u_ac_controller_soc_inst.u_picorv32.count_instr[1] ),
    .X(_06147_));
 sg13g2_buf_2 place9796 (.A(net9795),
    .X(net9796));
 sg13g2_nand4_1 _24358_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[3] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[4] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[2] ),
    .Y(_06149_),
    .D(_06147_));
 sg13g2_buf_2 place9795 (.A(_09902_),
    .X(net9795));
 sg13g2_and2_1 _24360_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_instr[7] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_instr[8] ),
    .X(_06151_));
 sg13g2_nand4_1 _24361_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[6] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[9] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[5] ),
    .Y(_06152_),
    .D(_06151_));
 sg13g2_buf_2 place9804 (.A(_08417_),
    .X(net9804));
 sg13g2_nor2_2 _24363_ (.A(_06149_),
    .B(_06152_),
    .Y(_06154_));
 sg13g2_xnor2_1 _24364_ (.Y(_06155_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[10] ),
    .B(_06154_));
 sg13g2_nor2_1 _24365_ (.A(net11017),
    .B(_06155_),
    .Y(_00595_));
 sg13g2_nand2_1 _24366_ (.Y(_06156_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[10] ),
    .B(_06154_));
 sg13g2_xnor2_1 _24367_ (.Y(_06157_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[11] ),
    .B(_06156_));
 sg13g2_and2_1 _24368_ (.A(net11049),
    .B(_06157_),
    .X(_00596_));
 sg13g2_nand3_1 _24369_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[11] ),
    .C(_06154_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[10] ),
    .Y(_06158_));
 sg13g2_xor2_1 _24370_ (.B(_06158_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[12] ),
    .X(_06159_));
 sg13g2_nor2_1 _24371_ (.A(net11017),
    .B(_06159_),
    .Y(_00597_));
 sg13g2_buf_2 place9791 (.A(_09911_),
    .X(net9791));
 sg13g2_buf_2 place9832 (.A(_11364_),
    .X(net9832));
 sg13g2_nand4_1 _24374_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[11] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[12] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[10] ),
    .Y(_06162_),
    .D(_06154_));
 sg13g2_xor2_1 _24375_ (.B(_06162_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[13] ),
    .X(_06163_));
 sg13g2_nor2_1 _24376_ (.A(net11017),
    .B(_06163_),
    .Y(_00598_));
 sg13g2_inv_2 _24377_ (.Y(_06164_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[14] ));
 sg13g2_nand4_1 _24378_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[11] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[12] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[10] ),
    .Y(_06165_),
    .D(\u_ac_controller_soc_inst.u_picorv32.count_instr[13] ));
 sg13g2_or3_1 _24379_ (.A(_06149_),
    .B(_06152_),
    .C(_06165_),
    .X(_06166_));
 sg13g2_xnor2_1 _24380_ (.Y(_06167_),
    .A(_06164_),
    .B(_06166_));
 sg13g2_nor2_1 _24381_ (.A(net11028),
    .B(_06167_),
    .Y(_00599_));
 sg13g2_nor2_2 _24382_ (.A(_06164_),
    .B(_06166_),
    .Y(_06168_));
 sg13g2_xnor2_1 _24383_ (.Y(_06169_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[15] ),
    .B(_06168_));
 sg13g2_nor2_1 _24384_ (.A(net11028),
    .B(_06169_),
    .Y(_00600_));
 sg13g2_nand2_1 _24385_ (.Y(_06170_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[15] ),
    .B(_06168_));
 sg13g2_xor2_1 _24386_ (.B(_06170_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[16] ),
    .X(_06171_));
 sg13g2_nor2_1 _24387_ (.A(net11028),
    .B(_06171_),
    .Y(_00601_));
 sg13g2_inv_2 _24388_ (.Y(_06172_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[17] ));
 sg13g2_nand3_1 _24389_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[16] ),
    .C(_06168_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[15] ),
    .Y(_06173_));
 sg13g2_xnor2_1 _24390_ (.Y(_06174_),
    .A(_06172_),
    .B(_06173_));
 sg13g2_nor2_1 _24391_ (.A(net11028),
    .B(_06174_),
    .Y(_00602_));
 sg13g2_nor2_2 _24392_ (.A(_06172_),
    .B(_06173_),
    .Y(_06175_));
 sg13g2_xnor2_1 _24393_ (.Y(_06176_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[18] ),
    .B(_06175_));
 sg13g2_nor2_1 _24394_ (.A(net11028),
    .B(_06176_),
    .Y(_00603_));
 sg13g2_nand2_1 _24395_ (.Y(_06177_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[18] ),
    .B(_06175_));
 sg13g2_xor2_1 _24396_ (.B(_06177_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[19] ),
    .X(_06178_));
 sg13g2_nor2_1 _24397_ (.A(net11028),
    .B(_06178_),
    .Y(_00604_));
 sg13g2_nand3_1 _24398_ (.B(\u_ac_controller_soc_inst.u_picorv32.decoder_trigger ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[0] ),
    .A(net10715),
    .Y(_06179_));
 sg13g2_xor2_1 _24399_ (.B(_06179_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[1] ),
    .X(_06180_));
 sg13g2_nor2_1 _24400_ (.A(net11022),
    .B(_06180_),
    .Y(_00605_));
 sg13g2_nand3_1 _24401_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[19] ),
    .C(_06175_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[18] ),
    .Y(_06181_));
 sg13g2_xor2_1 _24402_ (.B(_06181_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[20] ),
    .X(_06182_));
 sg13g2_nor2_1 _24403_ (.A(net11028),
    .B(_06182_),
    .Y(_00606_));
 sg13g2_or2_1 _24404_ (.X(_06183_),
    .B(_06165_),
    .A(_06164_));
 sg13g2_and4_1 _24405_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_instr[15] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_instr[16] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[17] ),
    .D(\u_ac_controller_soc_inst.u_picorv32.count_instr[18] ),
    .X(_06184_));
 sg13g2_nand3_1 _24406_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[20] ),
    .C(_06184_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[19] ),
    .Y(_06185_));
 sg13g2_nor4_2 _24407_ (.A(_06149_),
    .B(_06152_),
    .C(_06183_),
    .Y(_06186_),
    .D(_06185_));
 sg13g2_xnor2_1 _24408_ (.Y(_06187_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[21] ),
    .B(_06186_));
 sg13g2_nor2_1 _24409_ (.A(net11031),
    .B(_06187_),
    .Y(_00607_));
 sg13g2_buf_2 place9792 (.A(_09911_),
    .X(net9792));
 sg13g2_nand2_1 _24411_ (.Y(_06189_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[21] ),
    .B(_06186_));
 sg13g2_xor2_1 _24412_ (.B(_06189_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[22] ),
    .X(_06190_));
 sg13g2_nor2_1 _24413_ (.A(net11031),
    .B(_06190_),
    .Y(_00608_));
 sg13g2_and3_2 _24414_ (.X(_06191_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[21] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_instr[22] ),
    .C(_06186_));
 sg13g2_buf_2 place9810 (.A(_07936_),
    .X(net9810));
 sg13g2_xnor2_1 _24416_ (.Y(_06193_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[23] ),
    .B(_06191_));
 sg13g2_nor2_1 _24417_ (.A(net11031),
    .B(_06193_),
    .Y(_00609_));
 sg13g2_nand2_1 _24418_ (.Y(_06194_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[23] ),
    .B(_06191_));
 sg13g2_xor2_1 _24419_ (.B(_06194_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[24] ),
    .X(_06195_));
 sg13g2_nor2_1 _24420_ (.A(net11031),
    .B(_06195_),
    .Y(_00610_));
 sg13g2_inv_2 _24421_ (.Y(_06196_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[25] ));
 sg13g2_nand3_1 _24422_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[24] ),
    .C(_06191_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[23] ),
    .Y(_06197_));
 sg13g2_xnor2_1 _24423_ (.Y(_06198_),
    .A(_06196_),
    .B(_06197_));
 sg13g2_nor2_1 _24424_ (.A(net11029),
    .B(_06198_),
    .Y(_00611_));
 sg13g2_nor2_1 _24425_ (.A(_06196_),
    .B(_06197_),
    .Y(_06199_));
 sg13g2_xor2_1 _24426_ (.B(_06199_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[26] ),
    .X(_06200_));
 sg13g2_and2_1 _24427_ (.A(net11053),
    .B(_06200_),
    .X(_00612_));
 sg13g2_nand2_1 _24428_ (.Y(_06201_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[26] ),
    .B(_06199_));
 sg13g2_xor2_1 _24429_ (.B(_06201_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[27] ),
    .X(_06202_));
 sg13g2_nor2_1 _24430_ (.A(net11029),
    .B(_06202_),
    .Y(_00613_));
 sg13g2_inv_2 _24431_ (.Y(_06203_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[28] ));
 sg13g2_nand4_1 _24432_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[22] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[23] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[21] ),
    .Y(_06204_),
    .D(\u_ac_controller_soc_inst.u_picorv32.count_instr[24] ));
 sg13g2_nor2_1 _24433_ (.A(_06196_),
    .B(_06204_),
    .Y(_06205_));
 sg13g2_nand4_1 _24434_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[27] ),
    .C(_06186_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[26] ),
    .Y(_06206_),
    .D(_06205_));
 sg13g2_xnor2_1 _24435_ (.Y(_06207_),
    .A(_06203_),
    .B(_06206_));
 sg13g2_nor2_1 _24436_ (.A(net11029),
    .B(_06207_),
    .Y(_00614_));
 sg13g2_nor2_2 _24437_ (.A(_06203_),
    .B(_06206_),
    .Y(_06208_));
 sg13g2_xnor2_1 _24438_ (.Y(_06209_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[29] ),
    .B(_06208_));
 sg13g2_nor2_1 _24439_ (.A(net11030),
    .B(_06209_),
    .Y(_00615_));
 sg13g2_xnor2_1 _24440_ (.Y(_06210_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[2] ),
    .B(_06147_));
 sg13g2_nor2_1 _24441_ (.A(net11016),
    .B(_06210_),
    .Y(_00616_));
 sg13g2_nand2_1 _24442_ (.Y(_06211_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[29] ),
    .B(_06208_));
 sg13g2_xor2_1 _24443_ (.B(_06211_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[30] ),
    .X(_06212_));
 sg13g2_nor2_1 _24444_ (.A(net11030),
    .B(_06212_),
    .Y(_00617_));
 sg13g2_inv_2 _24445_ (.Y(_06213_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[31] ));
 sg13g2_nand3_1 _24446_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[30] ),
    .C(_06208_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[29] ),
    .Y(_06214_));
 sg13g2_xnor2_1 _24447_ (.Y(_06215_),
    .A(_06213_),
    .B(_06214_));
 sg13g2_nor2_1 _24448_ (.A(net11029),
    .B(_06215_),
    .Y(_00618_));
 sg13g2_buf_2 place9794 (.A(net9793),
    .X(net9794));
 sg13g2_nor2_2 _24450_ (.A(_06213_),
    .B(_06214_),
    .Y(_06217_));
 sg13g2_xnor2_1 _24451_ (.Y(_06218_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[32] ),
    .B(_06217_));
 sg13g2_nor2_1 _24452_ (.A(net11029),
    .B(_06218_),
    .Y(_00619_));
 sg13g2_nand2_1 _24453_ (.Y(_06219_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[32] ),
    .B(_06217_));
 sg13g2_xor2_1 _24454_ (.B(_06219_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[33] ),
    .X(_06220_));
 sg13g2_nor2_1 _24455_ (.A(net11027),
    .B(_06220_),
    .Y(_00620_));
 sg13g2_nand3_1 _24456_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[33] ),
    .C(_06217_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[32] ),
    .Y(_06221_));
 sg13g2_xor2_1 _24457_ (.B(_06221_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[34] ),
    .X(_06222_));
 sg13g2_nor2_1 _24458_ (.A(net11027),
    .B(_06222_),
    .Y(_00621_));
 sg13g2_nand4_1 _24459_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[33] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[34] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[32] ),
    .Y(_06223_),
    .D(_06217_));
 sg13g2_xor2_1 _24460_ (.B(_06223_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[35] ),
    .X(_06224_));
 sg13g2_nor2_1 _24461_ (.A(net11027),
    .B(_06224_),
    .Y(_00622_));
 sg13g2_nand4_1 _24462_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[33] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[34] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[32] ),
    .Y(_06225_),
    .D(\u_ac_controller_soc_inst.u_picorv32.count_instr[35] ));
 sg13g2_nor2_1 _24463_ (.A(_06213_),
    .B(_06225_),
    .Y(_06226_));
 sg13g2_and4_2 _24464_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_instr[29] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_instr[30] ),
    .C(_06208_),
    .D(_06226_),
    .X(_06227_));
 sg13g2_buf_2 place9789 (.A(net9788),
    .X(net9789));
 sg13g2_xnor2_1 _24466_ (.Y(_06229_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[36] ),
    .B(_06227_));
 sg13g2_nor2_1 _24467_ (.A(net11016),
    .B(_06229_),
    .Y(_00623_));
 sg13g2_nand2_1 _24468_ (.Y(_06230_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[36] ),
    .B(_06227_));
 sg13g2_xor2_1 _24469_ (.B(_06230_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[37] ),
    .X(_06231_));
 sg13g2_nor2_1 _24470_ (.A(net11016),
    .B(_06231_),
    .Y(_00624_));
 sg13g2_inv_2 _24471_ (.Y(_06232_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[38] ));
 sg13g2_nand3_1 _24472_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[37] ),
    .C(_06227_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[36] ),
    .Y(_06233_));
 sg13g2_buf_2 place9793 (.A(net9792),
    .X(net9793));
 sg13g2_xnor2_1 _24474_ (.Y(_06235_),
    .A(_06232_),
    .B(_06233_));
 sg13g2_nor2_1 _24475_ (.A(net11011),
    .B(_06235_),
    .Y(_00625_));
 sg13g2_nor2_2 _24476_ (.A(_06232_),
    .B(_06233_),
    .Y(_06236_));
 sg13g2_xnor2_1 _24477_ (.Y(_06237_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[39] ),
    .B(_06236_));
 sg13g2_nor2_1 _24478_ (.A(net11011),
    .B(_06237_),
    .Y(_00626_));
 sg13g2_nand2_1 _24479_ (.Y(_06238_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[2] ),
    .B(_06147_));
 sg13g2_xor2_1 _24480_ (.B(_06238_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[3] ),
    .X(_06239_));
 sg13g2_nor2_1 _24481_ (.A(net11016),
    .B(_06239_),
    .Y(_00627_));
 sg13g2_nand2_1 _24482_ (.Y(_06240_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[39] ),
    .B(_06236_));
 sg13g2_xor2_1 _24483_ (.B(_06240_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[40] ),
    .X(_06241_));
 sg13g2_nor2_1 _24484_ (.A(net11011),
    .B(_06241_),
    .Y(_00628_));
 sg13g2_buf_2 place9779 (.A(net9778),
    .X(net9779));
 sg13g2_and3_1 _24486_ (.X(_06243_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[39] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_instr[40] ),
    .C(_06236_));
 sg13g2_xnor2_1 _24487_ (.Y(_06244_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[41] ),
    .B(_06243_));
 sg13g2_nor2_1 _24488_ (.A(net11011),
    .B(_06244_),
    .Y(_00629_));
 sg13g2_nand2_1 _24489_ (.Y(_06245_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[41] ),
    .B(_06243_));
 sg13g2_xor2_1 _24490_ (.B(_06245_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[42] ),
    .X(_06246_));
 sg13g2_nor2_1 _24491_ (.A(net11011),
    .B(_06246_),
    .Y(_00630_));
 sg13g2_inv_2 _24492_ (.Y(_06247_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[43] ));
 sg13g2_or2_1 _24493_ (.X(_06248_),
    .B(_06233_),
    .A(_06232_));
 sg13g2_nand4_1 _24494_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[40] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[41] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[39] ),
    .Y(_06249_),
    .D(\u_ac_controller_soc_inst.u_picorv32.count_instr[42] ));
 sg13g2_or2_1 _24495_ (.X(_06250_),
    .B(_06249_),
    .A(_06248_));
 sg13g2_xnor2_1 _24496_ (.Y(_06251_),
    .A(_06247_),
    .B(_06250_));
 sg13g2_nor2_1 _24497_ (.A(net11017),
    .B(_06251_),
    .Y(_00631_));
 sg13g2_nor2_2 _24498_ (.A(_06247_),
    .B(_06250_),
    .Y(_06252_));
 sg13g2_xnor2_1 _24499_ (.Y(_06253_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[44] ),
    .B(_06252_));
 sg13g2_nor2_1 _24500_ (.A(net11017),
    .B(_06253_),
    .Y(_00632_));
 sg13g2_inv_2 _24501_ (.Y(_06254_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[45] ));
 sg13g2_nand2_2 _24502_ (.Y(_06255_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[44] ),
    .B(_06252_));
 sg13g2_xnor2_1 _24503_ (.Y(_06256_),
    .A(_06254_),
    .B(_06255_));
 sg13g2_nor2_1 _24504_ (.A(net11017),
    .B(_06256_),
    .Y(_00633_));
 sg13g2_nor2_1 _24505_ (.A(_06254_),
    .B(_06255_),
    .Y(_06257_));
 sg13g2_xnor2_1 _24506_ (.Y(_06258_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[46] ),
    .B(_06257_));
 sg13g2_nor2_1 _24507_ (.A(net11017),
    .B(_06258_),
    .Y(_00634_));
 sg13g2_inv_1 _24508_ (.Y(_06259_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[46] ));
 sg13g2_nor3_1 _24509_ (.A(_06254_),
    .B(_06259_),
    .C(_06255_),
    .Y(_06260_));
 sg13g2_xnor2_1 _24510_ (.Y(_06261_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[47] ),
    .B(_06260_));
 sg13g2_nor2_1 _24511_ (.A(net11017),
    .B(_06261_),
    .Y(_00635_));
 sg13g2_nand4_1 _24512_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[45] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[46] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[44] ),
    .Y(_06262_),
    .D(\u_ac_controller_soc_inst.u_picorv32.count_instr[47] ));
 sg13g2_nor4_2 _24513_ (.A(_06247_),
    .B(_06248_),
    .C(_06249_),
    .Y(_06263_),
    .D(_06262_));
 sg13g2_xnor2_1 _24514_ (.Y(_06264_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[48] ),
    .B(_06263_));
 sg13g2_nor2_1 _24515_ (.A(net11027),
    .B(_06264_),
    .Y(_00636_));
 sg13g2_and2_1 _24516_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_instr[48] ),
    .B(_06263_),
    .X(_06265_));
 sg13g2_buf_2 place9788 (.A(net9787),
    .X(net9788));
 sg13g2_xnor2_1 _24518_ (.Y(_06267_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[49] ),
    .B(net9682));
 sg13g2_nor2_1 _24519_ (.A(net11031),
    .B(_06267_),
    .Y(_00637_));
 sg13g2_nand3_1 _24520_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[3] ),
    .C(_06147_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[2] ),
    .Y(_06268_));
 sg13g2_xor2_1 _24521_ (.B(_06268_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[4] ),
    .X(_06269_));
 sg13g2_nor2_1 _24522_ (.A(net11016),
    .B(_06269_),
    .Y(_00638_));
 sg13g2_buf_2 place9787 (.A(net9786),
    .X(net9787));
 sg13g2_nand2_2 _24524_ (.Y(_06271_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[49] ),
    .B(net9682));
 sg13g2_xor2_1 _24525_ (.B(_06271_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[50] ),
    .X(_06272_));
 sg13g2_nor2_1 _24526_ (.A(net11031),
    .B(_06272_),
    .Y(_00639_));
 sg13g2_nand3_1 _24527_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[50] ),
    .C(net9682),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[49] ),
    .Y(_06273_));
 sg13g2_xor2_1 _24528_ (.B(_06273_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[51] ),
    .X(_06274_));
 sg13g2_nor2_1 _24529_ (.A(net11030),
    .B(_06274_),
    .Y(_00640_));
 sg13g2_nand4_1 _24530_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[50] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[51] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[49] ),
    .Y(_06275_),
    .D(_06265_));
 sg13g2_xor2_1 _24531_ (.B(_06275_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[52] ),
    .X(_06276_));
 sg13g2_nor2_1 _24532_ (.A(net11030),
    .B(_06276_),
    .Y(_00641_));
 sg13g2_nand3_1 _24533_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[51] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[52] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[50] ),
    .Y(_06277_));
 sg13g2_nor2_1 _24534_ (.A(_06271_),
    .B(_06277_),
    .Y(_06278_));
 sg13g2_xnor2_1 _24535_ (.Y(_06279_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[53] ),
    .B(_06278_));
 sg13g2_nor2_1 _24536_ (.A(net11030),
    .B(_06279_),
    .Y(_00642_));
 sg13g2_nand4_1 _24537_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[51] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[52] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[50] ),
    .Y(_06280_),
    .D(\u_ac_controller_soc_inst.u_picorv32.count_instr[53] ));
 sg13g2_nor2_1 _24538_ (.A(_06271_),
    .B(_06280_),
    .Y(_06281_));
 sg13g2_xnor2_1 _24539_ (.Y(_06282_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[54] ),
    .B(_06281_));
 sg13g2_nor2_1 _24540_ (.A(net11031),
    .B(_06282_),
    .Y(_00643_));
 sg13g2_nand2_1 _24541_ (.Y(_06283_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[49] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_instr[54] ));
 sg13g2_nor2_1 _24542_ (.A(_06280_),
    .B(_06283_),
    .Y(_06284_));
 sg13g2_nand2_1 _24543_ (.Y(_06285_),
    .A(net9682),
    .B(_06284_));
 sg13g2_xor2_1 _24544_ (.B(_06285_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[55] ),
    .X(_06286_));
 sg13g2_nor2_1 _24545_ (.A(net11031),
    .B(_06286_),
    .Y(_00644_));
 sg13g2_and2_1 _24546_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_instr[55] ),
    .B(_06284_),
    .X(_06287_));
 sg13g2_buf_2 place9834 (.A(net9833),
    .X(net9834));
 sg13g2_nand2_1 _24548_ (.Y(_06289_),
    .A(net9682),
    .B(_06287_));
 sg13g2_xor2_1 _24549_ (.B(_06289_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[56] ),
    .X(_06290_));
 sg13g2_nor2_1 _24550_ (.A(net11021),
    .B(_06290_),
    .Y(_00645_));
 sg13g2_nand3_1 _24551_ (.B(net9682),
    .C(_06287_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[56] ),
    .Y(_06291_));
 sg13g2_xor2_1 _24552_ (.B(_06291_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[57] ),
    .X(_06292_));
 sg13g2_nor2_1 _24553_ (.A(net11021),
    .B(_06292_),
    .Y(_00646_));
 sg13g2_and3_2 _24554_ (.X(_06293_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[56] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_instr[57] ),
    .C(_06287_));
 sg13g2_buf_2 place9770 (.A(net9766),
    .X(net9770));
 sg13g2_nand2_1 _24556_ (.Y(_06295_),
    .A(net9682),
    .B(_06293_));
 sg13g2_xor2_1 _24557_ (.B(_06295_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[58] ),
    .X(_06296_));
 sg13g2_nor2_1 _24558_ (.A(net11021),
    .B(_06296_),
    .Y(_00647_));
 sg13g2_nand3_1 _24559_ (.B(net9682),
    .C(_06293_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[58] ),
    .Y(_06297_));
 sg13g2_xor2_1 _24560_ (.B(_06297_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[59] ),
    .X(_06298_));
 sg13g2_nor2_1 _24561_ (.A(net11021),
    .B(_06298_),
    .Y(_00648_));
 sg13g2_buf_2 place9775 (.A(net9773),
    .X(net9775));
 sg13g2_xor2_1 _24563_ (.B(_06149_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[5] ),
    .X(_06300_));
 sg13g2_nor2_1 _24564_ (.A(net11011),
    .B(_06300_),
    .Y(_00649_));
 sg13g2_and4_2 _24565_ (.A(\u_ac_controller_soc_inst.u_picorv32.count_instr[58] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_instr[59] ),
    .C(_06265_),
    .D(_06293_),
    .X(_06301_));
 sg13g2_buf_2 place9777 (.A(net9772),
    .X(net9777));
 sg13g2_xnor2_1 _24567_ (.Y(_06303_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[60] ),
    .B(_06301_));
 sg13g2_nor2_1 _24568_ (.A(net11024),
    .B(_06303_),
    .Y(_00650_));
 sg13g2_nand2_1 _24569_ (.Y(_06304_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[60] ),
    .B(_06301_));
 sg13g2_xor2_1 _24570_ (.B(_06304_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[61] ),
    .X(_06305_));
 sg13g2_nor2_1 _24571_ (.A(net11024),
    .B(_06305_),
    .Y(_00651_));
 sg13g2_nand3_1 _24572_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[61] ),
    .C(_06301_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[60] ),
    .Y(_06306_));
 sg13g2_xor2_1 _24573_ (.B(_06306_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[62] ),
    .X(_06307_));
 sg13g2_nor2_1 _24574_ (.A(net11024),
    .B(_06307_),
    .Y(_00652_));
 sg13g2_nand4_1 _24575_ (.B(\u_ac_controller_soc_inst.u_picorv32.count_instr[61] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.count_instr[62] ),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[60] ),
    .Y(_06308_),
    .D(_06301_));
 sg13g2_xor2_1 _24576_ (.B(_06308_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[63] ),
    .X(_06309_));
 sg13g2_nor2_1 _24577_ (.A(net11020),
    .B(_06309_),
    .Y(_00653_));
 sg13g2_inv_1 _24578_ (.Y(_06310_),
    .A(_06149_));
 sg13g2_nand2_1 _24579_ (.Y(_06311_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[5] ),
    .B(_06310_));
 sg13g2_xnor2_1 _24580_ (.Y(_06312_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[6] ),
    .B(_06311_));
 sg13g2_and2_1 _24581_ (.A(net11049),
    .B(_06312_),
    .X(_00654_));
 sg13g2_and3_2 _24582_ (.X(_06313_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[5] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.count_instr[6] ),
    .C(_06310_));
 sg13g2_buf_2 place9778 (.A(net9777),
    .X(net9778));
 sg13g2_xnor2_1 _24584_ (.Y(_06315_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[7] ),
    .B(_06313_));
 sg13g2_nor2_1 _24585_ (.A(net11010),
    .B(_06315_),
    .Y(_00655_));
 sg13g2_nand2_1 _24586_ (.Y(_06316_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[7] ),
    .B(_06313_));
 sg13g2_xor2_1 _24587_ (.B(_06316_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[8] ),
    .X(_06317_));
 sg13g2_nor2_1 _24588_ (.A(net11011),
    .B(_06317_),
    .Y(_00656_));
 sg13g2_nand2_1 _24589_ (.Y(_06318_),
    .A(_06151_),
    .B(_06313_));
 sg13g2_xor2_1 _24590_ (.B(_06318_),
    .A(\u_ac_controller_soc_inst.u_picorv32.count_instr[9] ),
    .X(_06319_));
 sg13g2_nor2_1 _24591_ (.A(net11011),
    .B(_06319_),
    .Y(_00657_));
 sg13g2_inv_1 _24592_ (.Y(_01729_),
    .A(_08387_));
 sg13g2_buf_2 place10736 (.A(net10735),
    .X(net10736));
 sg13g2_and2_1 _24594_ (.A(\u_ac_controller_soc_inst.u_picorv32.is_alu_reg_reg ),
    .B(_11570_),
    .X(_06321_));
 sg13g2_buf_2 place9762 (.A(net9761),
    .X(net9762));
 sg13g2_nor2_1 _24596_ (.A(net10376),
    .B(_11526_),
    .Y(_06323_));
 sg13g2_a22oi_1 _24597_ (.Y(_06324_),
    .B1(_06321_),
    .B2(_06323_),
    .A2(net10378),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_add ));
 sg13g2_nor2_1 _24598_ (.A(net11014),
    .B(_06324_),
    .Y(_01730_));
 sg13g2_and2_1 _24599_ (.A(_00121_),
    .B(_11525_),
    .X(_06325_));
 sg13g2_buf_2 place9755 (.A(_05334_),
    .X(net9755));
 sg13g2_a22oi_1 _24601_ (.Y(_06327_),
    .B1(_06325_),
    .B2(_11575_),
    .A2(net10378),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_addi ));
 sg13g2_nor2_1 _24602_ (.A(net11015),
    .B(_06327_),
    .Y(_01731_));
 sg13g2_nand3_1 _24603_ (.B(\u_ac_controller_soc_inst.u_picorv32.instr_and ),
    .C(net10373),
    .A(net11053),
    .Y(_06328_));
 sg13g2_nor2b_2 _24604_ (.A(_00123_),
    .B_N(_11570_),
    .Y(_06329_));
 sg13g2_nand3_1 _24605_ (.B(net10607),
    .C(net10608),
    .A(net11053),
    .Y(_06330_));
 sg13g2_nor2_2 _24606_ (.A(_00121_),
    .B(_06330_),
    .Y(_06331_));
 sg13g2_nand3_1 _24607_ (.B(_06329_),
    .C(_06331_),
    .A(net10273),
    .Y(_06332_));
 sg13g2_nand2_1 _24608_ (.Y(_01732_),
    .A(_06328_),
    .B(_06332_));
 sg13g2_and3_1 _24609_ (.X(_06333_),
    .A(net11053),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_andi ),
    .C(net10373));
 sg13g2_a21o_1 _24610_ (.A2(_06331_),
    .A1(_11571_),
    .B1(_06333_),
    .X(_01733_));
 sg13g2_buf_2 place9833 (.A(net9832),
    .X(net9833));
 sg13g2_nor2_2 _24612_ (.A(_00102_),
    .B(net10376),
    .Y(_06335_));
 sg13g2_a22oi_1 _24613_ (.Y(_06336_),
    .B1(_06325_),
    .B2(_06335_),
    .A2(net10378),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_beq ));
 sg13g2_nor2_1 _24614_ (.A(net11014),
    .B(_06336_),
    .Y(_01735_));
 sg13g2_nand2_1 _24615_ (.Y(_06337_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_bge ),
    .B(net10365));
 sg13g2_nand2b_1 _24616_ (.Y(_06338_),
    .B(_06335_),
    .A_N(_11539_));
 sg13g2_a21oi_1 _24617_ (.A1(_06337_),
    .A2(_06338_),
    .Y(_01736_),
    .B1(net11019));
 sg13g2_nor2_2 _24618_ (.A(_08861_),
    .B(_11418_),
    .Y(_06339_));
 sg13g2_nor3_1 _24619_ (.A(net11019),
    .B(_08850_),
    .C(net10273),
    .Y(_06340_));
 sg13g2_a21o_1 _24620_ (.A2(_06339_),
    .A1(_06331_),
    .B1(_06340_),
    .X(_01737_));
 sg13g2_a22oi_1 _24621_ (.Y(_06341_),
    .B1(_11532_),
    .B2(_06339_),
    .A2(net10375),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_blt ));
 sg13g2_nor2_1 _24622_ (.A(net11025),
    .B(_06341_),
    .Y(_01738_));
 sg13g2_nor2_2 _24623_ (.A(_00121_),
    .B(_11544_),
    .Y(_06342_));
 sg13g2_a22oi_1 _24624_ (.Y(_06343_),
    .B1(_06339_),
    .B2(_06342_),
    .A2(net10375),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_bltu ));
 sg13g2_nor2_1 _24625_ (.A(net11025),
    .B(_06343_),
    .Y(_01739_));
 sg13g2_a22oi_1 _24626_ (.Y(_06344_),
    .B1(_11537_),
    .B2(_06339_),
    .A2(net10373),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_bne ));
 sg13g2_nor2_1 _24627_ (.A(net11019),
    .B(_06344_),
    .Y(_01740_));
 sg13g2_nand2_1 _24628_ (.Y(_06345_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_fence ),
    .B(net10378));
 sg13g2_nor4_2 _24629_ (.A(_11551_),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[4] ),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[5] ),
    .Y(_06346_),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[6] ));
 sg13g2_nand4_1 _24630_ (.B(_06325_),
    .C(_04017_),
    .A(net10274),
    .Y(_06347_),
    .D(_06346_));
 sg13g2_a21oi_1 _24631_ (.A1(_06345_),
    .A2(_06347_),
    .Y(_01741_),
    .B1(net11014));
 sg13g2_nand2_1 _24632_ (.Y(_06348_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_or ),
    .B(net10375));
 sg13g2_nand3_1 _24633_ (.B(_06329_),
    .C(_06342_),
    .A(net10273),
    .Y(_06349_));
 sg13g2_a21oi_1 _24634_ (.A1(_06348_),
    .A2(_06349_),
    .Y(_01750_),
    .B1(net11026));
 sg13g2_a22oi_1 _24635_ (.Y(_06350_),
    .B1(_11571_),
    .B2(_06342_),
    .A2(net10375),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_ori ));
 sg13g2_nor2_1 _24636_ (.A(net11025),
    .B(_06350_),
    .Y(_01751_));
 sg13g2_nor2_1 _24637_ (.A(net10372),
    .B(_11567_),
    .Y(_06351_));
 sg13g2_a22oi_1 _24638_ (.Y(_06352_),
    .B1(_06329_),
    .B2(_06351_),
    .A2(net10372),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_sll ));
 sg13g2_nor2_1 _24639_ (.A(net11018),
    .B(_06352_),
    .Y(_01758_));
 sg13g2_nor2_1 _24640_ (.A(net10374),
    .B(_11541_),
    .Y(_06353_));
 sg13g2_a22oi_1 _24641_ (.Y(_06354_),
    .B1(_06321_),
    .B2(_06353_),
    .A2(net10374),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_slt ));
 sg13g2_nor2_1 _24642_ (.A(net11025),
    .B(_06354_),
    .Y(_01760_));
 sg13g2_nor2_1 _24643_ (.A(_11541_),
    .B(_11577_),
    .Y(_06355_));
 sg13g2_a21oi_1 _24644_ (.A1(\u_ac_controller_soc_inst.u_picorv32.instr_slti ),
    .A2(net10374),
    .Y(_06356_),
    .B1(_06355_));
 sg13g2_nor2_1 _24645_ (.A(net11025),
    .B(_06356_),
    .Y(_01761_));
 sg13g2_nand4_1 _24646_ (.B(net10607),
    .C(net10608),
    .A(net11053),
    .Y(_06357_),
    .D(_00121_));
 sg13g2_nand3_1 _24647_ (.B(\u_ac_controller_soc_inst.u_picorv32.instr_sltiu ),
    .C(net10374),
    .A(net11053),
    .Y(_06358_));
 sg13g2_o21ai_1 _24648_ (.B1(_06358_),
    .Y(_01762_),
    .A1(_11577_),
    .A2(_06357_));
 sg13g2_nand3_1 _24649_ (.B(\u_ac_controller_soc_inst.u_picorv32.instr_sltu ),
    .C(net10374),
    .A(net11053),
    .Y(_06359_));
 sg13g2_inv_1 _24650_ (.Y(_06360_),
    .A(_06357_));
 sg13g2_nand3_1 _24651_ (.B(_06321_),
    .C(_06360_),
    .A(net10273),
    .Y(_06361_));
 sg13g2_nand2_1 _24652_ (.Y(_01763_),
    .A(_06359_),
    .B(_06361_));
 sg13g2_inv_1 _24653_ (.Y(_06362_),
    .A(_11585_));
 sg13g2_a22oi_1 _24654_ (.Y(_06363_),
    .B1(_11574_),
    .B2(_06362_),
    .A2(net10372),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_sra ));
 sg13g2_nor2_1 _24655_ (.A(net11018),
    .B(_06363_),
    .Y(_01764_));
 sg13g2_nor2_1 _24656_ (.A(net10374),
    .B(_11539_),
    .Y(_06364_));
 sg13g2_a22oi_1 _24657_ (.Y(_06365_),
    .B1(_06321_),
    .B2(_06364_),
    .A2(net10374),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_srl ));
 sg13g2_nor2_1 _24658_ (.A(net11018),
    .B(_06365_),
    .Y(_01766_));
 sg13g2_buf_2 place9763 (.A(net9762),
    .X(net9763));
 sg13g2_buf_2 place9761 (.A(_05143_),
    .X(net9761));
 sg13g2_buf_2 place9754 (.A(net9753),
    .X(net9754));
 sg13g2_nor3_1 _24662_ (.A(_11526_),
    .B(_11573_),
    .C(_11585_),
    .Y(_06369_));
 sg13g2_a21oi_1 _24663_ (.A1(net10633),
    .A2(net10376),
    .Y(_06370_),
    .B1(_06369_));
 sg13g2_nor2_1 _24664_ (.A(net11014),
    .B(_06370_),
    .Y(_01768_));
 sg13g2_nand2_1 _24665_ (.Y(_06371_),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_xor ),
    .B(net10373));
 sg13g2_nand3_1 _24666_ (.B(_11532_),
    .C(_06329_),
    .A(net10273),
    .Y(_06372_));
 sg13g2_a21oi_1 _24667_ (.A1(_06371_),
    .A2(_06372_),
    .Y(_01770_),
    .B1(net11018));
 sg13g2_a22oi_1 _24668_ (.Y(_06373_),
    .B1(_11532_),
    .B2(_11571_),
    .A2(net10375),
    .A1(\u_ac_controller_soc_inst.u_picorv32.instr_xori ));
 sg13g2_nor2_1 _24669_ (.A(net11025),
    .B(_06373_),
    .Y(_01771_));
 sg13g2_a22oi_1 _24670_ (.Y(_06374_),
    .B1(_04027_),
    .B2(_04033_),
    .A2(_08581_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.is_beq_bne_blt_bge_bltu_bgeu ));
 sg13g2_nor2_1 _24671_ (.A(net11013),
    .B(_06374_),
    .Y(_01774_));
 sg13g2_a21oi_1 _24672_ (.A1(_08859_),
    .A2(_08864_),
    .Y(_06375_),
    .B1(_08861_));
 sg13g2_nor2_1 _24673_ (.A(\u_ac_controller_soc_inst.u_picorv32.is_beq_bne_blt_bge_bltu_bgeu ),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_jalr ),
    .Y(_06376_));
 sg13g2_or2_1 _24674_ (.X(_06377_),
    .B(_06376_),
    .A(_08378_));
 sg13g2_nand2_2 _24675_ (.Y(_06378_),
    .A(net10658),
    .B(net10661));
 sg13g2_nand2_1 _24676_ (.Y(_06379_),
    .A(\u_ac_controller_soc_inst.u_picorv32.latched_branch ),
    .B(_09847_));
 sg13g2_o21ai_1 _24677_ (.B1(_06379_),
    .Y(_06380_),
    .A1(_09847_),
    .A2(_06378_));
 sg13g2_nand3_1 _24678_ (.B(_08395_),
    .C(_06380_),
    .A(net11052),
    .Y(_06381_));
 sg13g2_o21ai_1 _24679_ (.B1(_06381_),
    .Y(_01781_),
    .A1(_06375_),
    .A2(_06377_));
 sg13g2_mux2_1 _24680_ (.A0(_11933_),
    .A1(_00088_),
    .S(_07942_),
    .X(_06382_));
 sg13g2_o21ai_1 _24681_ (.B1(_06382_),
    .Y(_06383_),
    .A1(net10695),
    .A2(net10722));
 sg13g2_a21oi_1 _24682_ (.A1(_07697_),
    .A2(_07940_),
    .Y(_06384_),
    .B1(net10610));
 sg13g2_a21oi_1 _24683_ (.A1(_00088_),
    .A2(_07942_),
    .Y(_06385_),
    .B1(_06384_));
 sg13g2_nor2_1 _24684_ (.A(_07949_),
    .B(_06385_),
    .Y(_06386_));
 sg13g2_a22oi_1 _24685_ (.Y(_06387_),
    .B1(_06386_),
    .B2(\u_ac_controller_soc_inst.u_picorv32.instr_lb ),
    .A2(_06383_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.latched_is_lb ));
 sg13g2_nor2_1 _24686_ (.A(net11013),
    .B(_06387_),
    .Y(_01782_));
 sg13g2_a22oi_1 _24687_ (.Y(_06388_),
    .B1(_06386_),
    .B2(\u_ac_controller_soc_inst.u_picorv32.instr_lh ),
    .A2(_06383_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.latched_is_lh ));
 sg13g2_nor2_1 _24688_ (.A(net11013),
    .B(_06388_),
    .Y(_01783_));
 sg13g2_o21ai_1 _24689_ (.B1(\u_ac_controller_soc_inst.u_picorv32.latched_stalu ),
    .Y(_06389_),
    .A1(_09847_),
    .A2(net10710));
 sg13g2_nand2_1 _24690_ (.Y(_06390_),
    .A(net10709),
    .B(_00102_));
 sg13g2_a21oi_1 _24691_ (.A1(_06389_),
    .A2(_06390_),
    .Y(_01789_),
    .B1(net11034));
 sg13g2_a22oi_1 _24692_ (.Y(_06391_),
    .B1(_08945_),
    .B2(_04749_),
    .A2(_08322_),
    .A1(net10714));
 sg13g2_nor2_1 _24693_ (.A(\u_ac_controller_soc_inst.u_picorv32.latched_store ),
    .B(_06391_),
    .Y(_06392_));
 sg13g2_nor2_1 _24694_ (.A(net11034),
    .B(_06392_),
    .Y(_06393_));
 sg13g2_nand3b_1 _24695_ (.B(_06393_),
    .C(\u_ac_controller_soc_inst.u_picorv32.cpu_state[3] ),
    .Y(_06394_),
    .A_N(_00110_));
 sg13g2_nand3_1 _24696_ (.B(_08390_),
    .C(_09819_),
    .A(_07949_),
    .Y(_06395_));
 sg13g2_buf_2 place9753 (.A(net9752),
    .X(net9753));
 sg13g2_nor2b_1 _24698_ (.A(net10722),
    .B_N(_00110_),
    .Y(_06397_));
 sg13g2_o21ai_1 _24699_ (.B1(_06393_),
    .Y(_06398_),
    .A1(_06395_),
    .A2(_06397_));
 sg13g2_o21ai_1 _24700_ (.B1(_06398_),
    .Y(_01790_),
    .A1(_06375_),
    .A2(_06394_));
 sg13g2_buf_2 place9752 (.A(_05334_),
    .X(net9752));
 sg13g2_nor2_1 _24702_ (.A(net10725),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[10] ),
    .Y(_06400_));
 sg13g2_buf_2 place9750 (.A(net9749),
    .X(net9750));
 sg13g2_mux2_1 _24704_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[8] ),
    .A1(_10107_),
    .S(net10350),
    .X(_06402_));
 sg13g2_buf_2 place9756 (.A(net9755),
    .X(net9756));
 sg13g2_nor2_2 _24706_ (.A(net10663),
    .B(net10259),
    .Y(_06404_));
 sg13g2_mux2_1 _24707_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[7] ),
    .A1(_10101_),
    .S(net10352),
    .X(_06405_));
 sg13g2_buf_2 place9748 (.A(_05438_),
    .X(net9748));
 sg13g2_inv_2 _24709_ (.Y(_06407_),
    .A(_06405_));
 sg13g2_mux2_1 _24710_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[2] ),
    .A1(_10045_),
    .S(net10353),
    .X(_06408_));
 sg13g2_buf_2 place9751 (.A(net9750),
    .X(net9751));
 sg13g2_nand2_2 _24712_ (.Y(_06410_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2] ),
    .B(_06408_));
 sg13g2_mux2_1 _24713_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[1] ),
    .A1(_09952_),
    .S(net10353),
    .X(_06411_));
 sg13g2_buf_2 place9747 (.A(_08207_),
    .X(net9747));
 sg13g2_or3_1 _24715_ (.A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[2] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2] ),
    .C(net10351),
    .X(_06413_));
 sg13g2_or3_1 _24716_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2] ),
    .B(_10045_),
    .C(_11612_),
    .X(_06414_));
 sg13g2_nand4_1 _24717_ (.B(_06411_),
    .C(_06413_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1] ),
    .Y(_06415_),
    .D(_06414_));
 sg13g2_buf_2 place9785 (.A(net9784),
    .X(net9785));
 sg13g2_nand2_1 _24719_ (.Y(_06417_),
    .A(_06410_),
    .B(_06415_));
 sg13g2_inv_2 _24720_ (.Y(_06418_),
    .A(_00131_));
 sg13g2_mux2_1 _24721_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[3] ),
    .A1(_10069_),
    .S(net10353),
    .X(_06419_));
 sg13g2_buf_2 place9784 (.A(net9783),
    .X(net9784));
 sg13g2_mux2_1 _24723_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[4] ),
    .A1(_10076_),
    .S(net10353),
    .X(_06421_));
 sg13g2_buf_2 place9745 (.A(net9744),
    .X(net9745));
 sg13g2_o21ai_1 _24725_ (.B1(_06421_),
    .Y(_06423_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3] ),
    .A2(_06419_));
 sg13g2_nor2_1 _24726_ (.A(_06418_),
    .B(_06423_),
    .Y(_06424_));
 sg13g2_nor2_1 _24727_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3] ),
    .B(_06419_),
    .Y(_06425_));
 sg13g2_nor3_1 _24728_ (.A(_00131_),
    .B(_06421_),
    .C(_06425_),
    .Y(_06426_));
 sg13g2_nand2_1 _24729_ (.Y(_06427_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3] ),
    .B(_06419_));
 sg13g2_nand3_1 _24730_ (.B(_06410_),
    .C(_06415_),
    .A(_06427_),
    .Y(_06428_));
 sg13g2_nand3_1 _24731_ (.B(_06421_),
    .C(_06419_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3] ),
    .Y(_06429_));
 sg13g2_nand2_1 _24732_ (.Y(_06430_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[4] ),
    .B(_06421_));
 sg13g2_o21ai_1 _24733_ (.B1(_06430_),
    .Y(_06431_),
    .A1(_06418_),
    .A2(_06429_));
 sg13g2_a221oi_1 _24734_ (.B2(_06428_),
    .C1(_06431_),
    .B1(_06426_),
    .A1(_06417_),
    .Y(_06432_),
    .A2(_06424_));
 sg13g2_buf_2 place9764 (.A(net9763),
    .X(net9764));
 sg13g2_mux2_1 _24736_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[6] ),
    .A1(_10092_),
    .S(net10353),
    .X(_06434_));
 sg13g2_buf_2 place9744 (.A(net9743),
    .X(net9744));
 sg13g2_and2_1 _24738_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[6] ),
    .B(_06434_),
    .X(_06436_));
 sg13g2_mux2_1 _24739_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[5] ),
    .A1(_10084_),
    .S(net10353),
    .X(_06437_));
 sg13g2_buf_2 place9746 (.A(_09919_),
    .X(net9746));
 sg13g2_nand2_1 _24741_ (.Y(_06439_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[5] ),
    .B(_06437_));
 sg13g2_nor2b_2 _24742_ (.A(_06436_),
    .B_N(_06439_),
    .Y(_06440_));
 sg13g2_or2_1 _24743_ (.X(_06441_),
    .B(_06437_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[5] ));
 sg13g2_or2_1 _24744_ (.X(_06442_),
    .B(_06434_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[6] ));
 sg13g2_a21oi_1 _24745_ (.A1(_06441_),
    .A2(_06442_),
    .Y(_06443_),
    .B1(_06436_));
 sg13g2_a221oi_1 _24746_ (.B2(_06440_),
    .C1(_06443_),
    .B1(_06432_),
    .A1(_04005_),
    .Y(_06444_),
    .A2(_06407_));
 sg13g2_buf_2 place9743 (.A(_09919_),
    .X(net9743));
 sg13g2_a221oi_1 _24748_ (.B2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[7] ),
    .C1(_06444_),
    .B1(_06405_),
    .A1(net10663),
    .Y(_06446_),
    .A2(net10259));
 sg13g2_buf_2 place9811 (.A(net9810),
    .X(net9811));
 sg13g2_nand2_1 _24750_ (.Y(_06448_),
    .A(_10115_),
    .B(net10351));
 sg13g2_and2_1 _24751_ (.A(_11786_),
    .B(_06448_),
    .X(_06449_));
 sg13g2_buf_2 place9735 (.A(_09938_),
    .X(net9735));
 sg13g2_o21ai_1 _24753_ (.B1(_06449_),
    .Y(_06451_),
    .A1(_06404_),
    .A2(_06446_));
 sg13g2_nor3_1 _24754_ (.A(_06449_),
    .B(_06404_),
    .C(_06446_),
    .Y(_06452_));
 sg13g2_a21oi_2 _24755_ (.B1(_06452_),
    .Y(_06453_),
    .A2(_06451_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[9] ));
 sg13g2_xnor2_1 _24756_ (.Y(_06454_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[10] ),
    .B(_06453_));
 sg13g2_and4_2 _24757_ (.A(_06421_),
    .B(net10258),
    .C(_06408_),
    .D(_06437_),
    .X(_06455_));
 sg13g2_buf_2 place9742 (.A(net9740),
    .X(net9742));
 sg13g2_nand3_1 _24759_ (.B(_06434_),
    .C(_06455_),
    .A(_06405_),
    .Y(_06457_));
 sg13g2_nand2b_2 _24760_ (.Y(_06458_),
    .B(_06402_),
    .A_N(_06457_));
 sg13g2_buf_2 place9741 (.A(net9740),
    .X(net9741));
 sg13g2_nor3_1 _24762_ (.A(net10653),
    .B(_06458_),
    .C(_06449_),
    .Y(_06460_));
 sg13g2_a21o_1 _24763_ (.A2(_06454_),
    .A1(net10653),
    .B1(_06460_),
    .X(_06461_));
 sg13g2_mux2_1 _24764_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[10] ),
    .A1(_09860_),
    .S(net10350),
    .X(_06462_));
 sg13g2_buf_2 place9739 (.A(_09928_),
    .X(net9739));
 sg13g2_inv_2 _24766_ (.Y(_06464_),
    .A(_06462_));
 sg13g2_a21oi_1 _24767_ (.A1(net10660),
    .A2(_06461_),
    .Y(_06465_),
    .B1(_06464_));
 sg13g2_and3_1 _24768_ (.X(_06466_),
    .A(net10660),
    .B(_06464_),
    .C(_06461_));
 sg13g2_nor3_1 _24769_ (.A(_09847_),
    .B(_06465_),
    .C(_06466_),
    .Y(_06467_));
 sg13g2_nor3_1 _24770_ (.A(net11033),
    .B(_06400_),
    .C(_06467_),
    .Y(_01864_));
 sg13g2_nor2_2 _24771_ (.A(_11501_),
    .B(net10380),
    .Y(_06468_));
 sg13g2_a21oi_1 _24772_ (.A1(_06464_),
    .A2(_06453_),
    .Y(_06469_),
    .B1(_03994_));
 sg13g2_nor2_1 _24773_ (.A(_06464_),
    .B(_06453_),
    .Y(_06470_));
 sg13g2_or3_1 _24774_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11] ),
    .B(_06469_),
    .C(_06470_),
    .X(_06471_));
 sg13g2_o21ai_1 _24775_ (.B1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11] ),
    .Y(_06472_),
    .A1(_06469_),
    .A2(_06470_));
 sg13g2_nand3_1 _24776_ (.B(_06471_),
    .C(_06472_),
    .A(_06468_),
    .Y(_06473_));
 sg13g2_mux2_1 _24777_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[9] ),
    .A1(_10115_),
    .S(net10351),
    .X(_06474_));
 sg13g2_buf_16 clkbuf_leaf_397_clk (.X(clknet_leaf_397_clk),
    .A(clknet_8_108_0_clk));
 sg13g2_nand2_2 _24779_ (.Y(_06476_),
    .A(_06462_),
    .B(_06474_));
 sg13g2_or3_1 _24780_ (.A(_04739_),
    .B(_06458_),
    .C(_06476_),
    .X(_06477_));
 sg13g2_nand2_1 _24781_ (.Y(_06478_),
    .A(_09872_),
    .B(_11605_));
 sg13g2_and2_1 _24782_ (.A(_11634_),
    .B(_06478_),
    .X(_06479_));
 sg13g2_buf_2 place9737 (.A(net9736),
    .X(net9737));
 sg13g2_nand2_1 _24784_ (.Y(_06481_),
    .A(net10275),
    .B(_06479_));
 sg13g2_a21oi_1 _24785_ (.A1(_06473_),
    .A2(_06477_),
    .Y(_06482_),
    .B1(_06481_));
 sg13g2_mux2_1 _24786_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[11] ),
    .A1(_09872_),
    .S(_11605_),
    .X(_06483_));
 sg13g2_buf_2 place9736 (.A(net9735),
    .X(net9736));
 sg13g2_nand4_1 _24788_ (.B(_06473_),
    .C(_06477_),
    .A(net10275),
    .Y(_06485_),
    .D(_06483_));
 sg13g2_nor2_2 _24789_ (.A(net11019),
    .B(net10715),
    .Y(_06486_));
 sg13g2_nand2_1 _24790_ (.Y(_06487_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[11] ),
    .B(_06486_));
 sg13g2_nand3b_1 _24791_ (.B(_06485_),
    .C(_06487_),
    .Y(_01865_),
    .A_N(_06482_));
 sg13g2_buf_2 place9734 (.A(_03758_),
    .X(net9734));
 sg13g2_mux2_1 _24793_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[12] ),
    .A1(_09881_),
    .S(net10351),
    .X(_06489_));
 sg13g2_buf_2 place9738 (.A(net9735),
    .X(net9738));
 sg13g2_nor2_2 _24795_ (.A(_04005_),
    .B(_06407_),
    .Y(_06491_));
 sg13g2_nand2_1 _24796_ (.Y(_06492_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[10] ),
    .B(_06462_));
 sg13g2_nand2b_1 _24797_ (.Y(_06493_),
    .B(_03994_),
    .A_N(_06462_));
 sg13g2_xnor2_1 _24798_ (.Y(_06494_),
    .A(_08527_),
    .B(_06483_));
 sg13g2_xnor2_1 _24799_ (.Y(_06495_),
    .A(_04011_),
    .B(_06474_));
 sg13g2_nand4_1 _24800_ (.B(_06493_),
    .C(_06494_),
    .A(_06492_),
    .Y(_06496_),
    .D(_06495_));
 sg13g2_xnor2_1 _24801_ (.Y(_06497_),
    .A(net10663),
    .B(net10259));
 sg13g2_nor2_1 _24802_ (.A(_06496_),
    .B(_06497_),
    .Y(_06498_));
 sg13g2_o21ai_1 _24803_ (.B1(_06498_),
    .Y(_06499_),
    .A1(_06444_),
    .A2(_06491_));
 sg13g2_a21oi_1 _24804_ (.A1(net10663),
    .A2(net10259),
    .Y(_06500_),
    .B1(_06474_));
 sg13g2_nand3_1 _24805_ (.B(net10259),
    .C(_06474_),
    .A(net10663),
    .Y(_06501_));
 sg13g2_o21ai_1 _24806_ (.B1(_06501_),
    .Y(_06502_),
    .A1(_04011_),
    .A2(_06500_));
 sg13g2_nor2_1 _24807_ (.A(_03994_),
    .B(_06464_),
    .Y(_06503_));
 sg13g2_a21oi_1 _24808_ (.A1(_06493_),
    .A2(_06502_),
    .Y(_06504_),
    .B1(_06503_));
 sg13g2_o21ai_1 _24809_ (.B1(_08527_),
    .Y(_06505_),
    .A1(_06479_),
    .A2(_06504_));
 sg13g2_nand2_1 _24810_ (.Y(_06506_),
    .A(_06479_),
    .B(_06504_));
 sg13g2_nand2_1 _24811_ (.Y(_06507_),
    .A(_06505_),
    .B(_06506_));
 sg13g2_nand2_1 _24812_ (.Y(_06508_),
    .A(_06499_),
    .B(_06507_));
 sg13g2_xor2_1 _24813_ (.B(_06508_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12] ),
    .X(_06509_));
 sg13g2_nor4_1 _24814_ (.A(net10653),
    .B(_06458_),
    .C(_06476_),
    .D(_06479_),
    .Y(_06510_));
 sg13g2_a21oi_2 _24815_ (.B1(_06510_),
    .Y(_06511_),
    .A2(_06509_),
    .A1(net10654));
 sg13g2_nor2_1 _24816_ (.A(net10379),
    .B(_06511_),
    .Y(_06512_));
 sg13g2_xnor2_1 _24817_ (.Y(_06513_),
    .A(_06489_),
    .B(_06512_));
 sg13g2_nor2_1 _24818_ (.A(net10726),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[12] ),
    .Y(_06514_));
 sg13g2_a21oi_1 _24819_ (.A1(net10726),
    .A2(_06513_),
    .Y(_06515_),
    .B1(_06514_));
 sg13g2_and2_1 _24820_ (.A(net11037),
    .B(_06515_),
    .X(_01866_));
 sg13g2_buf_2 place9733 (.A(_05893_),
    .X(net9733));
 sg13g2_mux2_1 _24822_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[13] ),
    .A1(_09889_),
    .S(_11605_),
    .X(_06517_));
 sg13g2_buf_2 place9731 (.A(_05893_),
    .X(net9731));
 sg13g2_buf_2 place9730 (.A(_05893_),
    .X(net9730));
 sg13g2_inv_1 _24825_ (.Y(_06520_),
    .A(_06489_));
 sg13g2_nand3_1 _24826_ (.B(_06499_),
    .C(_06507_),
    .A(_06520_),
    .Y(_06521_));
 sg13g2_a21oi_1 _24827_ (.A1(_06499_),
    .A2(_06507_),
    .Y(_06522_),
    .B1(_06520_));
 sg13g2_a21oi_2 _24828_ (.B1(_06522_),
    .Y(_06523_),
    .A2(_06521_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12] ));
 sg13g2_xnor2_1 _24829_ (.Y(_06524_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[13] ),
    .B(_06523_));
 sg13g2_or4_1 _24830_ (.A(_06458_),
    .B(_06476_),
    .C(_06479_),
    .D(_06520_),
    .X(_06525_));
 sg13g2_buf_2 place9732 (.A(_05893_),
    .X(net9732));
 sg13g2_nor2_1 _24832_ (.A(net10654),
    .B(_06525_),
    .Y(_06527_));
 sg13g2_a21oi_1 _24833_ (.A1(net10654),
    .A2(_06524_),
    .Y(_06528_),
    .B1(_06527_));
 sg13g2_nor2_1 _24834_ (.A(net10379),
    .B(_06528_),
    .Y(_06529_));
 sg13g2_xnor2_1 _24835_ (.Y(_06530_),
    .A(_06517_),
    .B(_06529_));
 sg13g2_o21ai_1 _24836_ (.B1(net11054),
    .Y(_06531_),
    .A1(net10725),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[13] ));
 sg13g2_a21oi_1 _24837_ (.A1(net10723),
    .A2(_06530_),
    .Y(_01867_),
    .B1(_06531_));
 sg13g2_nand2_1 _24838_ (.Y(_06532_),
    .A(_09898_),
    .B(net10349));
 sg13g2_nand2_2 _24839_ (.Y(_06533_),
    .A(_11651_),
    .B(_06532_));
 sg13g2_buf_2 place9726 (.A(_08209_),
    .X(net9726));
 sg13g2_nand2_1 _24841_ (.Y(_06535_),
    .A(_09889_),
    .B(net10349));
 sg13g2_and2_1 _24842_ (.A(_11646_),
    .B(_06535_),
    .X(_06536_));
 sg13g2_buf_2 place9727 (.A(net9726),
    .X(net9727));
 sg13g2_nand2_1 _24844_ (.Y(_06538_),
    .A(_06536_),
    .B(_06523_));
 sg13g2_o21ai_1 _24845_ (.B1(_03996_),
    .Y(_06539_),
    .A1(_06536_),
    .A2(_06523_));
 sg13g2_a21o_1 _24846_ (.A2(_06539_),
    .A1(_06538_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[14] ),
    .X(_06540_));
 sg13g2_a21oi_1 _24847_ (.A1(_06536_),
    .A2(_06523_),
    .Y(_06541_),
    .B1(_03998_));
 sg13g2_a21oi_1 _24848_ (.A1(_06539_),
    .A2(_06541_),
    .Y(_06542_),
    .B1(net10362));
 sg13g2_nor2_1 _24849_ (.A(_06536_),
    .B(_06525_),
    .Y(_06543_));
 sg13g2_a22oi_1 _24850_ (.Y(_06544_),
    .B1(_06543_),
    .B2(net10362),
    .A2(_06542_),
    .A1(_06540_));
 sg13g2_nor4_1 _24851_ (.A(_11410_),
    .B(_08332_),
    .C(_06533_),
    .D(_06544_),
    .Y(_06545_));
 sg13g2_nand3_1 _24852_ (.B(_06533_),
    .C(_06544_),
    .A(net10275),
    .Y(_06546_));
 sg13g2_nor2_2 _24853_ (.A(net10661),
    .B(_08332_),
    .Y(_06547_));
 sg13g2_a22oi_1 _24854_ (.Y(_06548_),
    .B1(_06533_),
    .B2(_06547_),
    .A2(_06486_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[14] ));
 sg13g2_nand3b_1 _24855_ (.B(_06546_),
    .C(_06548_),
    .Y(_01868_),
    .A_N(_06545_));
 sg13g2_mux2_1 _24856_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[15] ),
    .A1(_09906_),
    .S(net10349),
    .X(_06549_));
 sg13g2_buf_2 place9729 (.A(_08209_),
    .X(net9729));
 sg13g2_nor2_1 _24858_ (.A(_03996_),
    .B(_06536_),
    .Y(_06551_));
 sg13g2_nor2_1 _24859_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[13] ),
    .B(_06517_),
    .Y(_06552_));
 sg13g2_xnor2_1 _24860_ (.Y(_06553_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12] ),
    .B(_06489_));
 sg13g2_and2_1 _24861_ (.A(_11651_),
    .B(_06532_),
    .X(_06554_));
 sg13g2_buf_2 place9740 (.A(net9739),
    .X(net9740));
 sg13g2_xnor2_1 _24863_ (.Y(_06556_),
    .A(_03998_),
    .B(_06554_));
 sg13g2_or4_1 _24864_ (.A(_06551_),
    .B(_06552_),
    .C(_06553_),
    .D(_06556_),
    .X(_06557_));
 sg13g2_buf_16 clkbuf_leaf_398_clk (.X(clknet_leaf_398_clk),
    .A(clknet_8_108_0_clk));
 sg13g2_nand2_1 _24866_ (.Y(_06559_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[8] ),
    .B(net10259));
 sg13g2_nand2b_1 _24867_ (.Y(_06560_),
    .B(_06491_),
    .A_N(_06404_));
 sg13g2_a21oi_2 _24868_ (.B1(_06496_),
    .Y(_06561_),
    .A2(_06560_),
    .A1(_06559_));
 sg13g2_nand2_1 _24869_ (.Y(_06562_),
    .A(_10107_),
    .B(net10350));
 sg13g2_and2_1 _24870_ (.A(_11781_),
    .B(_06562_),
    .X(_06563_));
 sg13g2_nor2_1 _24871_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[7] ),
    .B(_06405_),
    .Y(_06564_));
 sg13g2_or3_1 _24872_ (.A(_06443_),
    .B(_06564_),
    .C(_06496_),
    .X(_06565_));
 sg13g2_a221oi_1 _24873_ (.B2(_06440_),
    .C1(_06565_),
    .B1(_06432_),
    .A1(_04008_),
    .Y(_06566_),
    .A2(_06563_));
 sg13g2_a21oi_1 _24874_ (.A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[9] ),
    .A2(_06474_),
    .Y(_06567_),
    .B1(_06462_));
 sg13g2_nand3_1 _24875_ (.B(_06462_),
    .C(_06474_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[9] ),
    .Y(_06568_));
 sg13g2_o21ai_1 _24876_ (.B1(_06568_),
    .Y(_06569_),
    .A1(_03994_),
    .A2(_06567_));
 sg13g2_and2_1 _24877_ (.A(_06494_),
    .B(_06569_),
    .X(_06570_));
 sg13g2_nor3_1 _24878_ (.A(_06561_),
    .B(_06566_),
    .C(_06570_),
    .Y(_06571_));
 sg13g2_nor2_1 _24879_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12] ),
    .B(_06489_),
    .Y(_06572_));
 sg13g2_a22oi_1 _24880_ (.Y(_06573_),
    .B1(_06489_),
    .B2(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12] ),
    .A2(_06483_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11] ));
 sg13g2_nor3_1 _24881_ (.A(_06552_),
    .B(_06572_),
    .C(_06573_),
    .Y(_06574_));
 sg13g2_nor3_1 _24882_ (.A(_06533_),
    .B(_06551_),
    .C(_06574_),
    .Y(_06575_));
 sg13g2_o21ai_1 _24883_ (.B1(_06533_),
    .Y(_06576_),
    .A1(_06551_),
    .A2(_06574_));
 sg13g2_o21ai_1 _24884_ (.B1(_06576_),
    .Y(_06577_),
    .A1(_03998_),
    .A2(_06575_));
 sg13g2_inv_1 _24885_ (.Y(_06578_),
    .A(_06577_));
 sg13g2_o21ai_1 _24886_ (.B1(_06578_),
    .Y(_06579_),
    .A1(_06557_),
    .A2(_06571_));
 sg13g2_buf_2 place9721 (.A(_09947_),
    .X(net9721));
 sg13g2_xnor2_1 _24888_ (.Y(_06581_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15] ),
    .B(_06579_));
 sg13g2_nor2_1 _24889_ (.A(net10362),
    .B(_06581_),
    .Y(_06582_));
 sg13g2_nand3_1 _24890_ (.B(_06489_),
    .C(_06517_),
    .A(_06483_),
    .Y(_06583_));
 sg13g2_or4_1 _24891_ (.A(_06458_),
    .B(_06476_),
    .C(_06554_),
    .D(_06583_),
    .X(_06584_));
 sg13g2_buf_2 place9728 (.A(net9726),
    .X(net9728));
 sg13g2_nor2_1 _24893_ (.A(net10652),
    .B(_06584_),
    .Y(_06586_));
 sg13g2_o21ai_1 _24894_ (.B1(net10660),
    .Y(_06587_),
    .A1(_06582_),
    .A2(_06586_));
 sg13g2_xnor2_1 _24895_ (.Y(_06588_),
    .A(net10257),
    .B(_06587_));
 sg13g2_buf_2 place9769 (.A(net9766),
    .X(net9769));
 sg13g2_nor2b_1 _24897_ (.A(net10723),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[15] ),
    .Y(_06590_));
 sg13g2_a21oi_1 _24898_ (.A1(net10723),
    .A2(_06588_),
    .Y(_06591_),
    .B1(_06590_));
 sg13g2_nor2_1 _24899_ (.A(net11034),
    .B(_06591_),
    .Y(_01869_));
 sg13g2_mux2_1 _24900_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[16] ),
    .A1(_09915_),
    .S(net10349),
    .X(_06592_));
 sg13g2_buf_2 place9724 (.A(net9723),
    .X(net9724));
 sg13g2_nand2_1 _24902_ (.Y(_06594_),
    .A(net10257),
    .B(_06579_));
 sg13g2_o21ai_1 _24903_ (.B1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15] ),
    .Y(_06595_),
    .A1(net10257),
    .A2(_06579_));
 sg13g2_a21oi_1 _24904_ (.A1(_06594_),
    .A2(_06595_),
    .Y(_06596_),
    .B1(_08500_));
 sg13g2_nand3_1 _24905_ (.B(_06594_),
    .C(_06595_),
    .A(_08500_),
    .Y(_06597_));
 sg13g2_nand3b_1 _24906_ (.B(net10652),
    .C(_06597_),
    .Y(_06598_),
    .A_N(_06596_));
 sg13g2_nand3b_1 _24907_ (.B(net10257),
    .C(net10362),
    .Y(_06599_),
    .A_N(_06584_));
 sg13g2_a21oi_1 _24908_ (.A1(_06598_),
    .A2(_06599_),
    .Y(_06600_),
    .B1(net10380));
 sg13g2_xnor2_1 _24909_ (.Y(_06601_),
    .A(_06592_),
    .B(_06600_));
 sg13g2_o21ai_1 _24910_ (.B1(net11054),
    .Y(_06602_),
    .A1(net10724),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[16] ));
 sg13g2_a21oi_1 _24911_ (.A1(net10724),
    .A2(_06601_),
    .Y(_01870_),
    .B1(_06602_));
 sg13g2_or2_1 _24912_ (.X(_06603_),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[17] ),
    .A(net10723));
 sg13g2_mux2_1 _24913_ (.A0(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[17] ),
    .A1(_09923_),
    .S(net10345),
    .X(_06604_));
 sg13g2_buf_2 place9776 (.A(net9775),
    .X(net9776));
 sg13g2_xnor2_1 _24915_ (.Y(_06606_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[16] ),
    .B(_06592_));
 sg13g2_xnor2_1 _24916_ (.Y(_06607_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15] ),
    .B(_06549_));
 sg13g2_nor2_1 _24917_ (.A(_06606_),
    .B(_06607_),
    .Y(_06608_));
 sg13g2_a21oi_1 _24918_ (.A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15] ),
    .A2(_06549_),
    .Y(_06609_),
    .B1(_06592_));
 sg13g2_nand3_1 _24919_ (.B(_06549_),
    .C(_06592_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15] ),
    .Y(_06610_));
 sg13g2_o21ai_1 _24920_ (.B1(_06610_),
    .Y(_06611_),
    .A1(_08500_),
    .A2(_06609_));
 sg13g2_a21oi_1 _24921_ (.A1(_06579_),
    .A2(_06608_),
    .Y(_06612_),
    .B1(_06611_));
 sg13g2_xnor2_1 _24922_ (.Y(_06613_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17] ),
    .B(_06612_));
 sg13g2_and2_1 _24923_ (.A(_06549_),
    .B(_06592_),
    .X(_06614_));
 sg13g2_nor2b_2 _24924_ (.A(_06584_),
    .B_N(_06614_),
    .Y(_06615_));
 sg13g2_and2_1 _24925_ (.A(net10362),
    .B(_06615_),
    .X(_06616_));
 sg13g2_a21oi_2 _24926_ (.B1(_06616_),
    .Y(_06617_),
    .A2(_06613_),
    .A1(net10657));
 sg13g2_nor3_1 _24927_ (.A(net10380),
    .B(_06604_),
    .C(_06617_),
    .Y(_06618_));
 sg13g2_o21ai_1 _24928_ (.B1(_06604_),
    .Y(_06619_),
    .A1(net10380),
    .A2(_06617_));
 sg13g2_nand3b_1 _24929_ (.B(net10723),
    .C(_06619_),
    .Y(_06620_),
    .A_N(_06618_));
 sg13g2_and3_1 _24930_ (.X(_01871_),
    .A(net11054),
    .B(_06603_),
    .C(_06620_));
 sg13g2_nand2_1 _24931_ (.Y(_06621_),
    .A(_09933_),
    .B(net10345));
 sg13g2_nand2_2 _24932_ (.Y(_06622_),
    .A(_11671_),
    .B(_06621_));
 sg13g2_buf_2 place9723 (.A(net9722),
    .X(net9723));
 sg13g2_nor2_1 _24934_ (.A(net10382),
    .B(\u_ac_controller_soc_inst.u_picorv32.decoder_trigger ),
    .Y(_06624_));
 sg13g2_a22oi_1 _24935_ (.Y(_06625_),
    .B1(_06622_),
    .B2(_06624_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[18] ),
    .A1(net10382));
 sg13g2_or2_1 _24936_ (.X(_06626_),
    .B(_06622_),
    .A(_06145_));
 sg13g2_nand2_1 _24937_ (.Y(_06627_),
    .A(net10715),
    .B(_06622_));
 sg13g2_nor2_1 _24938_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17] ),
    .B(net10256),
    .Y(_06628_));
 sg13g2_nand2_1 _24939_ (.Y(_06629_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17] ),
    .B(net10256));
 sg13g2_o21ai_1 _24940_ (.B1(_06629_),
    .Y(_06630_),
    .A1(_06612_),
    .A2(_06628_));
 sg13g2_xor2_1 _24941_ (.B(_06630_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18] ),
    .X(_06631_));
 sg13g2_and2_1 _24942_ (.A(_11501_),
    .B(net10256),
    .X(_06632_));
 sg13g2_a22oi_1 _24943_ (.Y(_06633_),
    .B1(_06632_),
    .B2(_06615_),
    .A2(_06631_),
    .A1(net10657));
 sg13g2_mux2_1 _24944_ (.A0(_06626_),
    .A1(_06627_),
    .S(_06633_),
    .X(_06634_));
 sg13g2_buf_2 place9722 (.A(net9721),
    .X(net9722));
 sg13g2_a21oi_1 _24946_ (.A1(_06625_),
    .A2(_06634_),
    .Y(_01872_),
    .B1(net11019));
 sg13g2_buf_2 place9718 (.A(net9717),
    .X(net9718));
 sg13g2_nand2_2 _24948_ (.Y(_06637_),
    .A(_09943_),
    .B(net10345));
 sg13g2_and2_1 _24949_ (.A(_11676_),
    .B(_06637_),
    .X(_06638_));
 sg13g2_buf_2 place9871 (.A(net9870),
    .X(net9871));
 sg13g2_nand2_1 _24951_ (.Y(_06640_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18] ),
    .B(_06622_));
 sg13g2_nand2_1 _24952_ (.Y(_06641_),
    .A(net10256),
    .B(_06611_));
 sg13g2_o21ai_1 _24953_ (.B1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17] ),
    .Y(_06642_),
    .A1(net10256),
    .A2(_06611_));
 sg13g2_nand3_1 _24954_ (.B(_06641_),
    .C(_06642_),
    .A(_06640_),
    .Y(_06643_));
 sg13g2_o21ai_1 _24955_ (.B1(_06643_),
    .Y(_06644_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18] ),
    .A2(_06622_));
 sg13g2_xor2_1 _24956_ (.B(_06622_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18] ),
    .X(_06645_));
 sg13g2_nor2b_1 _24957_ (.A(_06628_),
    .B_N(_06629_),
    .Y(_06646_));
 sg13g2_and3_2 _24958_ (.X(_06647_),
    .A(_06608_),
    .B(_06645_),
    .C(_06646_));
 sg13g2_nor2b_1 _24959_ (.A(_06557_),
    .B_N(_06647_),
    .Y(_06648_));
 sg13g2_o21ai_1 _24960_ (.B1(_06648_),
    .Y(_06649_),
    .A1(_06561_),
    .A2(_06566_));
 sg13g2_nand2_1 _24961_ (.Y(_06650_),
    .A(_06494_),
    .B(_06569_));
 sg13g2_nor2_1 _24962_ (.A(_06557_),
    .B(_06650_),
    .Y(_06651_));
 sg13g2_o21ai_1 _24963_ (.B1(_06647_),
    .Y(_06652_),
    .A1(_06577_),
    .A2(_06651_));
 sg13g2_nand3_1 _24964_ (.B(_06649_),
    .C(_06652_),
    .A(_06644_),
    .Y(_06653_));
 sg13g2_buf_2 place9717 (.A(net9716),
    .X(net9717));
 sg13g2_xnor2_1 _24966_ (.Y(_06655_),
    .A(_00132_),
    .B(_06653_));
 sg13g2_nand2_1 _24967_ (.Y(_06656_),
    .A(net10657),
    .B(_06655_));
 sg13g2_nand3_1 _24968_ (.B(_06622_),
    .C(_06632_),
    .A(_06615_),
    .Y(_06657_));
 sg13g2_a21oi_1 _24969_ (.A1(_06656_),
    .A2(_06657_),
    .Y(_06658_),
    .B1(net10380));
 sg13g2_xnor2_1 _24970_ (.Y(_06659_),
    .A(_06638_),
    .B(_06658_));
 sg13g2_nor2b_1 _24971_ (.A(net10715),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[19] ),
    .Y(_06660_));
 sg13g2_a21oi_1 _24972_ (.A1(net10715),
    .A2(_06659_),
    .Y(_06661_),
    .B1(_06660_));
 sg13g2_nor2_1 _24973_ (.A(net11019),
    .B(_06661_),
    .Y(_01873_));
 sg13g2_nor2_1 _24974_ (.A(net10730),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[1] ),
    .Y(_06662_));
 sg13g2_nand2_1 _24975_ (.Y(_06663_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1] ),
    .B(_06468_));
 sg13g2_xnor2_1 _24976_ (.Y(_06664_),
    .A(_06411_),
    .B(_06663_));
 sg13g2_nor2_1 _24977_ (.A(net10383),
    .B(_06664_),
    .Y(_06665_));
 sg13g2_nor3_1 _24978_ (.A(net11003),
    .B(_06662_),
    .C(_06665_),
    .Y(_01874_));
 sg13g2_buf_2 place9720 (.A(net9716),
    .X(net9720));
 sg13g2_buf_2 place9719 (.A(net9718),
    .X(net9719));
 sg13g2_buf_2 place9749 (.A(net9748),
    .X(net9749));
 sg13g2_nand4_1 _24982_ (.B(_06644_),
    .C(_06649_),
    .A(_08518_),
    .Y(_06669_),
    .D(_06652_));
 sg13g2_buf_16 clkbuf_leaf_399_clk (.X(clknet_leaf_399_clk),
    .A(clknet_8_114_0_clk));
 sg13g2_nor2_1 _24984_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[19] ),
    .B(_00132_),
    .Y(_06671_));
 sg13g2_nor2_2 _24985_ (.A(_06638_),
    .B(_06671_),
    .Y(_06672_));
 sg13g2_nand2_2 _24986_ (.Y(_06673_),
    .A(_11676_),
    .B(_06637_));
 sg13g2_nor2_1 _24987_ (.A(_00132_),
    .B(_06673_),
    .Y(_06674_));
 sg13g2_a22oi_1 _24988_ (.Y(_06675_),
    .B1(_06674_),
    .B2(_06653_),
    .A2(_06672_),
    .A1(_06669_));
 sg13g2_buf_2 place9712 (.A(_09972_),
    .X(net9712));
 sg13g2_xnor2_1 _24990_ (.Y(_06677_),
    .A(_00133_),
    .B(_06675_));
 sg13g2_nand4_1 _24991_ (.B(_06614_),
    .C(_06622_),
    .A(net10256),
    .Y(_06678_),
    .D(_06673_));
 sg13g2_nor2_2 _24992_ (.A(_06584_),
    .B(_06678_),
    .Y(_06679_));
 sg13g2_nor2_1 _24993_ (.A(net10658),
    .B(_06679_),
    .Y(_06680_));
 sg13g2_a21oi_1 _24994_ (.A1(net10658),
    .A2(_06677_),
    .Y(_06681_),
    .B1(_06680_));
 sg13g2_nand2_1 _24995_ (.Y(_06682_),
    .A(net10661),
    .B(_06681_));
 sg13g2_nand2_1 _24996_ (.Y(_06683_),
    .A(_09959_),
    .B(net10348));
 sg13g2_and2_1 _24997_ (.A(_11683_),
    .B(_06683_),
    .X(_06684_));
 sg13g2_buf_2 place9715 (.A(net9712),
    .X(net9715));
 sg13g2_xnor2_1 _24999_ (.Y(_06686_),
    .A(_06682_),
    .B(_06684_));
 sg13g2_o21ai_1 _25000_ (.B1(net11054),
    .Y(_06687_),
    .A1(net10716),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[20] ));
 sg13g2_a21oi_1 _25001_ (.A1(net10716),
    .A2(_06686_),
    .Y(_01875_),
    .B1(_06687_));
 sg13g2_nand2_2 _25002_ (.Y(_06688_),
    .A(_11683_),
    .B(_06683_));
 sg13g2_buf_2 place9714 (.A(net9713),
    .X(net9714));
 sg13g2_nor2_1 _25004_ (.A(_00133_),
    .B(net10196),
    .Y(_06690_));
 sg13g2_nand2_1 _25005_ (.Y(_06691_),
    .A(_06675_),
    .B(_06690_));
 sg13g2_inv_2 _25006_ (.Y(_06692_),
    .A(net10666));
 sg13g2_buf_2 place9711 (.A(net9710),
    .X(net9711));
 sg13g2_nor2_2 _25008_ (.A(_04001_),
    .B(net10309),
    .Y(_06694_));
 sg13g2_a21oi_1 _25009_ (.A1(_00133_),
    .A2(_06675_),
    .Y(_06695_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20] ));
 sg13g2_o21ai_1 _25010_ (.B1(net10196),
    .Y(_06696_),
    .A1(_06694_),
    .A2(_06695_));
 sg13g2_a21o_1 _25011_ (.A2(_06696_),
    .A1(_06691_),
    .B1(net10364),
    .X(_06697_));
 sg13g2_nor4_2 _25012_ (.A(_06536_),
    .B(_06525_),
    .C(_06554_),
    .Y(_06698_),
    .D(_06678_));
 sg13g2_nand3_1 _25013_ (.B(_06698_),
    .C(net10196),
    .A(net10364),
    .Y(_06699_));
 sg13g2_nand2_1 _25014_ (.Y(_06700_),
    .A(_09967_),
    .B(net10345));
 sg13g2_and2_1 _25015_ (.A(_11690_),
    .B(_06700_),
    .X(_06701_));
 sg13g2_buf_2 place9716 (.A(_09963_),
    .X(net9716));
 sg13g2_nand3_1 _25017_ (.B(_09848_),
    .C(_06701_),
    .A(net10661),
    .Y(_06703_));
 sg13g2_a21o_1 _25018_ (.A2(_06699_),
    .A1(_06697_),
    .B1(_06703_),
    .X(_06704_));
 sg13g2_nand2_2 _25019_ (.Y(_06705_),
    .A(_11690_),
    .B(_06700_));
 sg13g2_buf_16 clkbuf_leaf_400_clk (.X(clknet_leaf_400_clk),
    .A(clknet_8_114_0_clk));
 sg13g2_nand4_1 _25021_ (.B(_06705_),
    .C(_06697_),
    .A(_09848_),
    .Y(_06707_),
    .D(_06699_));
 sg13g2_a22oi_1 _25022_ (.Y(_06708_),
    .B1(_06547_),
    .B2(_06705_),
    .A2(_06486_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[21] ));
 sg13g2_nand3_1 _25023_ (.B(_06707_),
    .C(_06708_),
    .A(_06704_),
    .Y(_01876_));
 sg13g2_nand3_1 _25024_ (.B(_06701_),
    .C(_06690_),
    .A(_06675_),
    .Y(_06709_));
 sg13g2_a21oi_1 _25025_ (.A1(_06705_),
    .A2(_06694_),
    .Y(_06710_),
    .B1(net10364));
 sg13g2_nand2_1 _25026_ (.Y(_06711_),
    .A(_06709_),
    .B(_06710_));
 sg13g2_o21ai_1 _25027_ (.B1(net10309),
    .Y(_06712_),
    .A1(net10196),
    .A2(_06705_));
 sg13g2_nor2_2 _25028_ (.A(_06684_),
    .B(_06701_),
    .Y(_06713_));
 sg13g2_nand2b_1 _25029_ (.Y(_06714_),
    .B(_06713_),
    .A_N(_06675_));
 sg13g2_a21oi_1 _25030_ (.A1(_06712_),
    .A2(_06714_),
    .Y(_06715_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20] ));
 sg13g2_a21oi_1 _25031_ (.A1(_06698_),
    .A2(_06713_),
    .Y(_06716_),
    .B1(net10659));
 sg13g2_nor2_1 _25032_ (.A(net10380),
    .B(_06716_),
    .Y(_06717_));
 sg13g2_o21ai_1 _25033_ (.B1(_06717_),
    .Y(_06718_),
    .A1(_06711_),
    .A2(_06715_));
 sg13g2_nand2_1 _25034_ (.Y(_06719_),
    .A(_09976_),
    .B(net10348));
 sg13g2_nand2_2 _25035_ (.Y(_06720_),
    .A(_11696_),
    .B(_06719_));
 sg13g2_buf_2 place9700 (.A(_08490_),
    .X(net9700));
 sg13g2_xor2_1 _25037_ (.B(net10195),
    .A(_06718_),
    .X(_06722_));
 sg13g2_o21ai_1 _25038_ (.B1(net11054),
    .Y(_06723_),
    .A1(net10716),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[22] ));
 sg13g2_a21oi_1 _25039_ (.A1(net10716),
    .A2(_06722_),
    .Y(_01877_),
    .B1(_06723_));
 sg13g2_nand2_1 _25040_ (.Y(_06724_),
    .A(_09984_),
    .B(net10348));
 sg13g2_and2_1 _25041_ (.A(_11701_),
    .B(_06724_),
    .X(_06725_));
 sg13g2_buf_2 place9710 (.A(_04607_),
    .X(net9710));
 sg13g2_nand3_1 _25043_ (.B(_06705_),
    .C(_06720_),
    .A(net10664),
    .Y(_06727_));
 sg13g2_buf_2 place9709 (.A(net9708),
    .X(net9709));
 sg13g2_nor2_1 _25045_ (.A(_06684_),
    .B(_06727_),
    .Y(_06729_));
 sg13g2_nand3_1 _25046_ (.B(_06672_),
    .C(_06729_),
    .A(_06669_),
    .Y(_06730_));
 sg13g2_buf_2 place9713 (.A(net9712),
    .X(net9713));
 sg13g2_or2_1 _25048_ (.X(_06732_),
    .B(_06720_),
    .A(_06705_));
 sg13g2_buf_2 place9780 (.A(_04813_),
    .X(net9780));
 sg13g2_o21ai_1 _25050_ (.B1(_06727_),
    .Y(_06734_),
    .A1(_00133_),
    .A2(_06732_));
 sg13g2_and2_1 _25051_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20] ),
    .B(_06734_),
    .X(_06735_));
 sg13g2_nor4_1 _25052_ (.A(_00132_),
    .B(_06673_),
    .C(_06684_),
    .D(_06727_),
    .Y(_06736_));
 sg13g2_a22oi_1 _25053_ (.Y(_06737_),
    .B1(_06736_),
    .B2(_06653_),
    .A2(_06735_),
    .A1(net10196));
 sg13g2_buf_2 place9702 (.A(net9700),
    .X(net9702));
 sg13g2_nand4_1 _25055_ (.B(_06644_),
    .C(_06649_),
    .A(_06638_),
    .Y(_06739_),
    .D(_06652_));
 sg13g2_buf_16 clkbuf_leaf_401_clk (.X(clknet_leaf_401_clk),
    .A(clknet_8_115_0_clk));
 sg13g2_mux2_1 _25057_ (.A0(_00132_),
    .A1(_06671_),
    .S(_06673_),
    .X(_06741_));
 sg13g2_nor4_1 _25058_ (.A(net10664),
    .B(_06688_),
    .C(_06732_),
    .D(_06741_),
    .Y(_06742_));
 sg13g2_nand3_1 _25059_ (.B(_06739_),
    .C(_06742_),
    .A(_06669_),
    .Y(_06743_));
 sg13g2_buf_2 place9701 (.A(net9700),
    .X(net9701));
 sg13g2_and3_2 _25061_ (.X(_06745_),
    .A(_06730_),
    .B(_06737_),
    .C(_06743_));
 sg13g2_buf_2 place9706 (.A(net9705),
    .X(net9706));
 sg13g2_nand2_1 _25063_ (.Y(_06747_),
    .A(net10667),
    .B(_06732_));
 sg13g2_a21o_1 _25064_ (.A2(_06747_),
    .A1(_06745_),
    .B1(_00133_),
    .X(_06748_));
 sg13g2_a21oi_1 _25065_ (.A1(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20] ),
    .A2(_06720_),
    .Y(_06749_),
    .B1(net10309));
 sg13g2_a21oi_1 _25066_ (.A1(_06745_),
    .A2(_06749_),
    .Y(_06750_),
    .B1(_06378_));
 sg13g2_nand3_1 _25067_ (.B(_06713_),
    .C(_06720_),
    .A(_06679_),
    .Y(_06751_));
 sg13g2_buf_2 place9693 (.A(_09980_),
    .X(net9693));
 sg13g2_nor2_1 _25069_ (.A(_04739_),
    .B(_06751_),
    .Y(_06753_));
 sg13g2_a21oi_1 _25070_ (.A1(_06748_),
    .A2(_06750_),
    .Y(_06754_),
    .B1(_06753_));
 sg13g2_xnor2_1 _25071_ (.Y(_06755_),
    .A(_06725_),
    .B(_06754_));
 sg13g2_nand2_1 _25072_ (.Y(_06756_),
    .A(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[23] ),
    .B(_06486_));
 sg13g2_o21ai_1 _25073_ (.B1(_06756_),
    .Y(_01878_),
    .A1(_08332_),
    .A2(_06755_));
 sg13g2_nand2_1 _25074_ (.Y(_06757_),
    .A(_09992_),
    .B(net10348));
 sg13g2_and2_1 _25075_ (.A(_11706_),
    .B(_06757_),
    .X(_06758_));
 sg13g2_buf_2 place9705 (.A(_08222_),
    .X(net9705));
 sg13g2_nor3_1 _25077_ (.A(net10664),
    .B(_06688_),
    .C(_06705_),
    .Y(_06760_));
 sg13g2_a21oi_1 _25078_ (.A1(net10664),
    .A2(_06713_),
    .Y(_06761_),
    .B1(_06760_));
 sg13g2_nor2_2 _25079_ (.A(_06741_),
    .B(_06761_),
    .Y(_06762_));
 sg13g2_nand2_2 _25080_ (.Y(_06763_),
    .A(_11701_),
    .B(_06724_));
 sg13g2_and2_1 _25081_ (.A(net10195),
    .B(_06763_),
    .X(_06764_));
 sg13g2_nand4_1 _25082_ (.B(_06739_),
    .C(_06762_),
    .A(_06669_),
    .Y(_06765_),
    .D(_06764_));
 sg13g2_a21oi_1 _25083_ (.A1(net10667),
    .A2(_06763_),
    .Y(_06766_),
    .B1(net10309));
 sg13g2_nor2_1 _25084_ (.A(net10195),
    .B(_06763_),
    .Y(_06767_));
 sg13g2_and3_1 _25085_ (.X(_06768_),
    .A(_06669_),
    .B(_06739_),
    .C(_06762_));
 sg13g2_nand2_1 _25086_ (.Y(_06769_),
    .A(net10667),
    .B(net10309));
 sg13g2_nor3_1 _25087_ (.A(_06688_),
    .B(_06763_),
    .C(_06732_),
    .Y(_06770_));
 sg13g2_o21ai_1 _25088_ (.B1(net10659),
    .Y(_06771_),
    .A1(_06769_),
    .A2(_06770_));
 sg13g2_a221oi_1 _25089_ (.B2(_06768_),
    .C1(_06771_),
    .B1(_06767_),
    .A1(_06765_),
    .Y(_06772_),
    .A2(_06766_));
 sg13g2_nor3_1 _25090_ (.A(net10659),
    .B(_06725_),
    .C(_06751_),
    .Y(_06773_));
 sg13g2_o21ai_1 _25091_ (.B1(net10662),
    .Y(_06774_),
    .A1(_06772_),
    .A2(_06773_));
 sg13g2_xnor2_1 _25092_ (.Y(_06775_),
    .A(_06758_),
    .B(_06774_));
 sg13g2_nor2_1 _25093_ (.A(net10719),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[24] ),
    .Y(_06776_));
 sg13g2_a21oi_1 _25094_ (.A1(net10719),
    .A2(_06775_),
    .Y(_06777_),
    .B1(_06776_));
 sg13g2_and2_1 _25095_ (.A(net11055),
    .B(_06777_),
    .X(_01879_));
 sg13g2_or2_1 _25096_ (.X(_06778_),
    .B(_06758_),
    .A(_06725_));
 sg13g2_buf_2 place9699 (.A(_08581_),
    .X(net9699));
 sg13g2_o21ai_1 _25098_ (.B1(net10364),
    .Y(_06780_),
    .A1(_06751_),
    .A2(_06778_));
 sg13g2_nand2_1 _25099_ (.Y(_06781_),
    .A(net10662),
    .B(_06780_));
 sg13g2_nand2_1 _25100_ (.Y(_06782_),
    .A(_10001_),
    .B(net10348));
 sg13g2_nand2_1 _25101_ (.Y(_06783_),
    .A(_11711_),
    .B(_06782_));
 sg13g2_buf_2 place9704 (.A(net9702),
    .X(net9704));
 sg13g2_nand2_1 _25103_ (.Y(_06785_),
    .A(net10721),
    .B(net10194));
 sg13g2_nor2_1 _25104_ (.A(_06781_),
    .B(_06785_),
    .Y(_06786_));
 sg13g2_nor2_1 _25105_ (.A(net10382),
    .B(net10194),
    .Y(_06787_));
 sg13g2_nand2_2 _25106_ (.Y(_06788_),
    .A(_06725_),
    .B(_06758_));
 sg13g2_buf_2 place9697 (.A(_09450_),
    .X(net9697));
 sg13g2_nor3_1 _25108_ (.A(net10665),
    .B(_06732_),
    .C(_06788_),
    .Y(_06790_));
 sg13g2_a21oi_1 _25109_ (.A1(_06730_),
    .A2(_06737_),
    .Y(_06791_),
    .B1(_06788_));
 sg13g2_and3_1 _25110_ (.X(_06792_),
    .A(net10664),
    .B(_06730_),
    .C(_06737_));
 sg13g2_o21ai_1 _25111_ (.B1(net10664),
    .Y(_06793_),
    .A1(_06725_),
    .A2(_06758_));
 sg13g2_o21ai_1 _25112_ (.B1(_06793_),
    .Y(_06794_),
    .A1(_06743_),
    .A2(_06788_));
 sg13g2_nor3_1 _25113_ (.A(_06791_),
    .B(_06792_),
    .C(_06794_),
    .Y(_06795_));
 sg13g2_nand2_1 _25114_ (.Y(_06796_),
    .A(net10667),
    .B(net10665));
 sg13g2_o21ai_1 _25115_ (.B1(net10659),
    .Y(_06797_),
    .A1(_06796_),
    .A2(_06758_));
 sg13g2_a221oi_1 _25116_ (.B2(_04001_),
    .C1(_06797_),
    .B1(_06795_),
    .A1(_06745_),
    .Y(_06798_),
    .A2(_06790_));
 sg13g2_mux2_1 _25117_ (.A0(_06786_),
    .A1(_06787_),
    .S(_06798_),
    .X(_06799_));
 sg13g2_o21ai_1 _25118_ (.B1(net11055),
    .Y(_06800_),
    .A1(net10721),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[25] ));
 sg13g2_a21oi_1 _25119_ (.A1(_06787_),
    .A2(_06781_),
    .Y(_06801_),
    .B1(_06800_));
 sg13g2_nor2b_1 _25120_ (.A(_06799_),
    .B_N(_06801_),
    .Y(_01880_));
 sg13g2_nand3_1 _25121_ (.B(_06713_),
    .C(_06720_),
    .A(_06698_),
    .Y(_06802_));
 sg13g2_buf_2 place9698 (.A(net9697),
    .X(net9698));
 sg13g2_nand2_1 _25123_ (.Y(_06804_),
    .A(net10364),
    .B(net10194));
 sg13g2_nor3_1 _25124_ (.A(_06802_),
    .B(_06778_),
    .C(_06804_),
    .Y(_06805_));
 sg13g2_nand2_1 _25125_ (.Y(_06806_),
    .A(net10662),
    .B(_06805_));
 sg13g2_nand3_1 _25126_ (.B(net10195),
    .C(_06783_),
    .A(net10666),
    .Y(_06807_));
 sg13g2_or4_1 _25127_ (.A(net10666),
    .B(net10195),
    .C(net10194),
    .D(_06788_),
    .X(_06808_));
 sg13g2_o21ai_1 _25128_ (.B1(_06808_),
    .Y(_06809_),
    .A1(_06778_),
    .A2(_06807_));
 sg13g2_nand4_1 _25129_ (.B(_06739_),
    .C(_06762_),
    .A(_06669_),
    .Y(_06810_),
    .D(_06809_));
 sg13g2_nor2_1 _25130_ (.A(_06732_),
    .B(_06788_),
    .Y(_06811_));
 sg13g2_a21oi_1 _25131_ (.A1(_06684_),
    .A2(_06811_),
    .Y(_06812_),
    .B1(net10665));
 sg13g2_o21ai_1 _25132_ (.B1(net10667),
    .Y(_06813_),
    .A1(net10194),
    .A2(_06812_));
 sg13g2_nor2_2 _25133_ (.A(_00133_),
    .B(_06378_),
    .Y(_06814_));
 sg13g2_nand3_1 _25134_ (.B(_06813_),
    .C(_06814_),
    .A(_06810_),
    .Y(_06815_));
 sg13g2_nand2_1 _25135_ (.Y(_06816_),
    .A(net10665),
    .B(_06468_));
 sg13g2_a21o_1 _25136_ (.A2(_06813_),
    .A1(_06810_),
    .B1(_06816_),
    .X(_06817_));
 sg13g2_nand3_1 _25137_ (.B(_06815_),
    .C(_06817_),
    .A(_06806_),
    .Y(_06818_));
 sg13g2_o21ai_1 _25138_ (.B1(_11716_),
    .Y(_06819_),
    .A1(_10012_),
    .A2(net10343));
 sg13g2_buf_2 place9707 (.A(net9705),
    .X(net9707));
 sg13g2_xor2_1 _25140_ (.B(_06819_),
    .A(_06818_),
    .X(_06821_));
 sg13g2_nor2b_1 _25141_ (.A(net10721),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[26] ),
    .Y(_06822_));
 sg13g2_a21oi_1 _25142_ (.A1(net10721),
    .A2(_06821_),
    .Y(_06823_),
    .B1(_06822_));
 sg13g2_nor2_1 _25143_ (.A(net11036),
    .B(_06823_),
    .Y(_01881_));
 sg13g2_nand2_2 _25144_ (.Y(_06824_),
    .A(_10019_),
    .B(net10348));
 sg13g2_nand2_2 _25145_ (.Y(_06825_),
    .A(_11721_),
    .B(_06824_));
 sg13g2_buf_16 clkbuf_leaf_410_clk (.X(clknet_leaf_410_clk),
    .A(clknet_8_101_0_clk));
 sg13g2_nor2_1 _25147_ (.A(_08332_),
    .B(_06825_),
    .Y(_06827_));
 sg13g2_a21oi_1 _25148_ (.A1(_11721_),
    .A2(_06824_),
    .Y(_06828_),
    .B1(_08332_));
 sg13g2_nor2_1 _25149_ (.A(net10194),
    .B(_06819_),
    .Y(_06829_));
 sg13g2_nand2_1 _25150_ (.Y(_06830_),
    .A(_06811_),
    .B(_06829_));
 sg13g2_nand2_1 _25151_ (.Y(_06831_),
    .A(net10667),
    .B(_06830_));
 sg13g2_and2_1 _25152_ (.A(_06814_),
    .B(_06831_),
    .X(_06832_));
 sg13g2_nand2_1 _25153_ (.Y(_06833_),
    .A(net10194),
    .B(_06819_));
 sg13g2_nor2_2 _25154_ (.A(_06778_),
    .B(_06833_),
    .Y(_06834_));
 sg13g2_nor2b_1 _25155_ (.A(_06788_),
    .B_N(_06829_),
    .Y(_06835_));
 sg13g2_mux2_1 _25156_ (.A0(_06834_),
    .A1(_06835_),
    .S(net10309),
    .X(_06836_));
 sg13g2_buf_2 place9786 (.A(_04813_),
    .X(net9786));
 sg13g2_nand2b_1 _25158_ (.Y(_06838_),
    .B(_06836_),
    .A_N(_06745_));
 sg13g2_nand3_1 _25159_ (.B(_06468_),
    .C(_06834_),
    .A(net10665),
    .Y(_06839_));
 sg13g2_nor2_1 _25160_ (.A(net10364),
    .B(_06796_),
    .Y(_06840_));
 sg13g2_and2_1 _25161_ (.A(net10662),
    .B(_06819_),
    .X(_06841_));
 sg13g2_o21ai_1 _25162_ (.B1(_06841_),
    .Y(_06842_),
    .A1(_06805_),
    .A2(_06840_));
 sg13g2_o21ai_1 _25163_ (.B1(_06842_),
    .Y(_06843_),
    .A1(_06745_),
    .A2(_06839_));
 sg13g2_a21oi_2 _25164_ (.B1(_06843_),
    .Y(_06844_),
    .A2(_06838_),
    .A1(_06832_));
 sg13g2_mux2_1 _25165_ (.A0(_06827_),
    .A1(_06828_),
    .S(_06844_),
    .X(_06845_));
 sg13g2_a21o_1 _25166_ (.A2(_06486_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[27] ),
    .B1(_06845_),
    .X(_01882_));
 sg13g2_nand2_1 _25167_ (.Y(_06846_),
    .A(_10028_),
    .B(net10348));
 sg13g2_nand2_1 _25168_ (.Y(_06847_),
    .A(_11726_),
    .B(_06846_));
 sg13g2_buf_2 place9684 (.A(_09997_),
    .X(net9684));
 sg13g2_nand3_1 _25170_ (.B(_06819_),
    .C(_06825_),
    .A(net10194),
    .Y(_06849_));
 sg13g2_or4_1 _25171_ (.A(_04739_),
    .B(_06802_),
    .C(_06778_),
    .D(_06849_),
    .X(_06850_));
 sg13g2_or2_1 _25172_ (.X(_06851_),
    .B(net10193),
    .A(_06819_));
 sg13g2_nand3_1 _25173_ (.B(_06819_),
    .C(net10193),
    .A(net10666),
    .Y(_06852_));
 sg13g2_o21ai_1 _25174_ (.B1(_06852_),
    .Y(_06853_),
    .A1(net10666),
    .A2(_06851_));
 sg13g2_and2_1 _25175_ (.A(_06809_),
    .B(_06853_),
    .X(_06854_));
 sg13g2_nand4_1 _25176_ (.B(_06739_),
    .C(_06762_),
    .A(_06669_),
    .Y(_06855_),
    .D(_06854_));
 sg13g2_buf_2 place9696 (.A(net9693),
    .X(net9696));
 sg13g2_nor2_1 _25178_ (.A(_06688_),
    .B(_06732_),
    .Y(_06857_));
 sg13g2_a21oi_1 _25179_ (.A1(_06857_),
    .A2(_06835_),
    .Y(_06858_),
    .B1(net10665));
 sg13g2_o21ai_1 _25180_ (.B1(net10667),
    .Y(_06859_),
    .A1(_06825_),
    .A2(_06858_));
 sg13g2_nand3_1 _25181_ (.B(_06855_),
    .C(_06859_),
    .A(_06814_),
    .Y(_06860_));
 sg13g2_a21o_1 _25182_ (.A2(_06859_),
    .A1(_06855_),
    .B1(_06816_),
    .X(_06861_));
 sg13g2_nand3_1 _25183_ (.B(_06860_),
    .C(_06861_),
    .A(_06850_),
    .Y(_06862_));
 sg13g2_xnor2_1 _25184_ (.Y(_06863_),
    .A(net10192),
    .B(_06862_));
 sg13g2_o21ai_1 _25185_ (.B1(net11055),
    .Y(_06864_),
    .A1(net10721),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[28] ));
 sg13g2_a21oi_1 _25186_ (.A1(net10721),
    .A2(_06863_),
    .Y(_01883_),
    .B1(_06864_));
 sg13g2_nand2_2 _25187_ (.Y(_06865_),
    .A(_10037_),
    .B(net10348));
 sg13g2_nand2_2 _25188_ (.Y(_06866_),
    .A(_11731_),
    .B(_06865_));
 sg13g2_buf_2 place9695 (.A(net9694),
    .X(net9695));
 sg13g2_buf_16 clkbuf_leaf_409_clk (.X(clknet_leaf_409_clk),
    .A(clknet_8_100_0_clk));
 sg13g2_nor2_1 _25191_ (.A(net10382),
    .B(_06866_),
    .Y(_06869_));
 sg13g2_a21oi_1 _25192_ (.A1(_11731_),
    .A2(_06865_),
    .Y(_06870_),
    .B1(_06145_));
 sg13g2_nand2_1 _25193_ (.Y(_06871_),
    .A(_06730_),
    .B(_06737_));
 sg13g2_inv_1 _25194_ (.Y(_06872_),
    .A(net10192));
 sg13g2_o21ai_1 _25195_ (.B1(_06692_),
    .Y(_06873_),
    .A1(_06830_),
    .A2(net10193));
 sg13g2_a21oi_2 _25196_ (.B1(_04001_),
    .Y(_06874_),
    .A2(_06873_),
    .A1(_06872_));
 sg13g2_nor3_1 _25197_ (.A(net10309),
    .B(_06871_),
    .C(_06874_),
    .Y(_06875_));
 sg13g2_nor3_1 _25198_ (.A(net10666),
    .B(net10193),
    .C(net10192),
    .Y(_06876_));
 sg13g2_nand2_2 _25199_ (.Y(_06877_),
    .A(_06836_),
    .B(_06876_));
 sg13g2_a21oi_1 _25200_ (.A1(_06730_),
    .A2(_06737_),
    .Y(_06878_),
    .B1(_06877_));
 sg13g2_and2_1 _25201_ (.A(net10193),
    .B(net10192),
    .X(_06879_));
 sg13g2_a21o_2 _25202_ (.A2(_06879_),
    .A1(net10666),
    .B1(_06876_),
    .X(_06880_));
 sg13g2_buf_16 clkbuf_leaf_408_clk (.X(clknet_leaf_408_clk),
    .A(clknet_8_100_0_clk));
 sg13g2_a221oi_1 _25204_ (.B2(_06834_),
    .C1(net10309),
    .B1(_06880_),
    .A1(net10667),
    .Y(_06882_),
    .A2(net10192));
 sg13g2_a21oi_1 _25205_ (.A1(_06692_),
    .A2(_06874_),
    .Y(_06883_),
    .B1(_06882_));
 sg13g2_o21ai_1 _25206_ (.B1(_06883_),
    .Y(_06884_),
    .A1(_06743_),
    .A2(_06877_));
 sg13g2_nor3_1 _25207_ (.A(_06875_),
    .B(_06878_),
    .C(_06884_),
    .Y(_06885_));
 sg13g2_mux2_1 _25208_ (.A0(_06869_),
    .A1(_06870_),
    .S(_06885_),
    .X(_06886_));
 sg13g2_nand2_1 _25209_ (.Y(_06887_),
    .A(net10662),
    .B(_06866_));
 sg13g2_nand2_2 _25210_ (.Y(_06888_),
    .A(_06834_),
    .B(_06879_));
 sg13g2_or2_1 _25211_ (.X(_06889_),
    .B(_06888_),
    .A(_06751_));
 sg13g2_mux2_1 _25212_ (.A0(_06887_),
    .A1(_06866_),
    .S(_06889_),
    .X(_06890_));
 sg13g2_nand3_1 _25213_ (.B(_11731_),
    .C(_06865_),
    .A(net10380),
    .Y(_06891_));
 sg13g2_o21ai_1 _25214_ (.B1(_06891_),
    .Y(_06892_),
    .A1(net10659),
    .A2(_06890_));
 sg13g2_o21ai_1 _25215_ (.B1(net11055),
    .Y(_06893_),
    .A1(net10716),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[29] ));
 sg13g2_a221oi_1 _25216_ (.B2(net10716),
    .C1(_06893_),
    .B1(_06892_),
    .A1(net10659),
    .Y(_01884_),
    .A2(_06886_));
 sg13g2_nand2_1 _25217_ (.Y(_06894_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1] ),
    .B(_06411_));
 sg13g2_xor2_1 _25218_ (.B(_06894_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2] ),
    .X(_06895_));
 sg13g2_a21oi_1 _25219_ (.A1(net10655),
    .A2(_06895_),
    .Y(_06896_),
    .B1(net10379));
 sg13g2_xnor2_1 _25220_ (.Y(_06897_),
    .A(_06408_),
    .B(_06896_));
 sg13g2_nand2_1 _25221_ (.Y(_06898_),
    .A(net10730),
    .B(_06897_));
 sg13g2_o21ai_1 _25222_ (.B1(_06898_),
    .Y(_06899_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[2] ),
    .A2(net10730));
 sg13g2_nor2_1 _25223_ (.A(net11003),
    .B(_06899_),
    .Y(_01885_));
 sg13g2_inv_1 _25224_ (.Y(_06900_),
    .A(_06859_));
 sg13g2_nor4_1 _25225_ (.A(net10665),
    .B(net10192),
    .C(_06900_),
    .D(net10191),
    .Y(_06901_));
 sg13g2_nand2_1 _25226_ (.Y(_06902_),
    .A(net10364),
    .B(net10191));
 sg13g2_nor3_1 _25227_ (.A(_06802_),
    .B(_06888_),
    .C(_06902_),
    .Y(_06903_));
 sg13g2_a221oi_1 _25228_ (.B2(_06855_),
    .C1(_06903_),
    .B1(_06901_),
    .A1(_06694_),
    .Y(_06904_),
    .A2(net10191));
 sg13g2_nand2_1 _25229_ (.Y(_06905_),
    .A(net10192),
    .B(net10191));
 sg13g2_o21ai_1 _25230_ (.B1(_06692_),
    .Y(_06906_),
    .A1(net10192),
    .A2(net10191));
 sg13g2_o21ai_1 _25231_ (.B1(_06906_),
    .Y(_06907_),
    .A1(_06855_),
    .A2(_06905_));
 sg13g2_nand2_1 _25232_ (.Y(_06908_),
    .A(_04001_),
    .B(_06907_));
 sg13g2_o21ai_1 _25233_ (.B1(net10662),
    .Y(_06909_),
    .A1(net10659),
    .A2(_06903_));
 sg13g2_a21oi_1 _25234_ (.A1(_06904_),
    .A2(_06908_),
    .Y(_06910_),
    .B1(_06909_));
 sg13g2_o21ai_1 _25235_ (.B1(_11745_),
    .Y(_06911_),
    .A1(_10054_),
    .A2(net10343));
 sg13g2_buf_16 clkbuf_leaf_407_clk (.X(clknet_leaf_407_clk),
    .A(clknet_8_112_0_clk));
 sg13g2_xnor2_1 _25237_ (.Y(_06913_),
    .A(_06910_),
    .B(_06911_));
 sg13g2_o21ai_1 _25238_ (.B1(net11055),
    .Y(_06914_),
    .A1(net10721),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[30] ));
 sg13g2_a21oi_1 _25239_ (.A1(net10721),
    .A2(_06913_),
    .Y(_01886_),
    .B1(_06914_));
 sg13g2_nand2_1 _25240_ (.Y(_06915_),
    .A(net10658),
    .B(_09848_));
 sg13g2_nor2_1 _25241_ (.A(_10063_),
    .B(net10342),
    .Y(_06916_));
 sg13g2_a21oi_2 _25242_ (.B1(_06916_),
    .Y(_06917_),
    .A2(net10341),
    .A1(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[31] ));
 sg13g2_nand2_1 _25243_ (.Y(_06918_),
    .A(net10661),
    .B(_06917_));
 sg13g2_nand4_1 _25244_ (.B(_06880_),
    .C(_06866_),
    .A(_06836_),
    .Y(_06919_),
    .D(_06911_));
 sg13g2_o21ai_1 _25245_ (.B1(_06692_),
    .Y(_06920_),
    .A1(_06866_),
    .A2(_06911_));
 sg13g2_o21ai_1 _25246_ (.B1(_06920_),
    .Y(_06921_),
    .A1(_06745_),
    .A2(_06919_));
 sg13g2_nor4_1 _25247_ (.A(net10665),
    .B(_06874_),
    .C(net10191),
    .D(_06911_),
    .Y(_06922_));
 sg13g2_nand3b_1 _25248_ (.B(_06836_),
    .C(_06880_),
    .Y(_06923_),
    .A_N(_06745_));
 sg13g2_and2_1 _25249_ (.A(_06694_),
    .B(_06911_),
    .X(_06924_));
 sg13g2_a221oi_1 _25250_ (.B2(_06923_),
    .C1(_06924_),
    .B1(_06922_),
    .A1(_04001_),
    .Y(_06925_),
    .A2(_06921_));
 sg13g2_mux2_1 _25251_ (.A0(_06918_),
    .A1(_06917_),
    .S(_06925_),
    .X(_06926_));
 sg13g2_nor2b_1 _25252_ (.A(_06917_),
    .B_N(_06624_),
    .Y(_06927_));
 sg13g2_a21o_1 _25253_ (.A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[31] ),
    .A1(net10382),
    .B1(_06927_),
    .X(_06928_));
 sg13g2_nand2_1 _25254_ (.Y(_06929_),
    .A(_06866_),
    .B(_06911_));
 sg13g2_nor2_2 _25255_ (.A(_06889_),
    .B(_06929_),
    .Y(_06930_));
 sg13g2_xnor2_1 _25256_ (.Y(_06931_),
    .A(_06917_),
    .B(_06930_));
 sg13g2_a22oi_1 _25257_ (.Y(_06932_),
    .B1(_06931_),
    .B2(_04740_),
    .A2(_06928_),
    .A1(net11054));
 sg13g2_o21ai_1 _25258_ (.B1(_06932_),
    .Y(_01887_),
    .A1(_06915_),
    .A2(_06926_));
 sg13g2_nor2_1 _25259_ (.A(net10730),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[3] ),
    .Y(_06933_));
 sg13g2_nor2_1 _25260_ (.A(_11492_),
    .B(_06408_),
    .Y(_06934_));
 sg13g2_o21ai_1 _25261_ (.B1(_06410_),
    .Y(_06935_),
    .A1(_06894_),
    .A2(_06934_));
 sg13g2_nand2_1 _25262_ (.Y(_06936_),
    .A(_08548_),
    .B(_06935_));
 sg13g2_and2_1 _25263_ (.A(_06410_),
    .B(_06415_),
    .X(_06937_));
 sg13g2_a22oi_1 _25264_ (.Y(_06938_),
    .B1(_06937_),
    .B2(_11503_),
    .A2(_06408_),
    .A1(net10363));
 sg13g2_a21oi_1 _25265_ (.A1(_06936_),
    .A2(_06938_),
    .Y(_06939_),
    .B1(net10379));
 sg13g2_xor2_1 _25266_ (.B(_06939_),
    .A(net10258),
    .X(_06940_));
 sg13g2_nor2_1 _25267_ (.A(net10383),
    .B(_06940_),
    .Y(_06941_));
 sg13g2_nor3_1 _25268_ (.A(net11032),
    .B(_06933_),
    .C(_06941_),
    .Y(_01888_));
 sg13g2_o21ai_1 _25269_ (.B1(_06427_),
    .Y(_06942_),
    .A1(_06425_),
    .A2(_06937_));
 sg13g2_xnor2_1 _25270_ (.Y(_06943_),
    .A(_06418_),
    .B(_06942_));
 sg13g2_nand3_1 _25271_ (.B(net10258),
    .C(_06408_),
    .A(net10363),
    .Y(_06944_));
 sg13g2_o21ai_1 _25272_ (.B1(_06944_),
    .Y(_06945_),
    .A1(net10363),
    .A2(_06943_));
 sg13g2_nand2_1 _25273_ (.Y(_06946_),
    .A(net10660),
    .B(_06945_));
 sg13g2_xor2_1 _25274_ (.B(_06946_),
    .A(_06421_),
    .X(_06947_));
 sg13g2_nand2_1 _25275_ (.Y(_06948_),
    .A(net10731),
    .B(_06947_));
 sg13g2_o21ai_1 _25276_ (.B1(_06948_),
    .Y(_06949_),
    .A1(net10731),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[4] ));
 sg13g2_nor2_1 _25277_ (.A(net11003),
    .B(_06949_),
    .Y(_01889_));
 sg13g2_buf_2 place9694 (.A(net9693),
    .X(net9694));
 sg13g2_nand4_1 _25279_ (.B(_06421_),
    .C(net10258),
    .A(net10363),
    .Y(_06951_),
    .D(_06408_));
 sg13g2_xnor2_1 _25280_ (.Y(_06952_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[5] ),
    .B(_06432_));
 sg13g2_nand2_1 _25281_ (.Y(_06953_),
    .A(net10655),
    .B(_06952_));
 sg13g2_a21o_1 _25282_ (.A2(_06953_),
    .A1(_06951_),
    .B1(net10379),
    .X(_06954_));
 sg13g2_xor2_1 _25283_ (.B(_06954_),
    .A(_06437_),
    .X(_06955_));
 sg13g2_nand2_1 _25284_ (.Y(_06956_),
    .A(net10731),
    .B(_06955_));
 sg13g2_o21ai_1 _25285_ (.B1(_06956_),
    .Y(_06957_),
    .A1(net10731),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[5] ));
 sg13g2_nor2_1 _25286_ (.A(_08213_),
    .B(_06957_),
    .Y(_01890_));
 sg13g2_nor2_1 _25287_ (.A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[5] ),
    .B(_06437_),
    .Y(_06958_));
 sg13g2_o21ai_1 _25288_ (.B1(_06439_),
    .Y(_06959_),
    .A1(_06958_),
    .A2(_06432_));
 sg13g2_xor2_1 _25289_ (.B(_06959_),
    .A(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[6] ),
    .X(_06960_));
 sg13g2_mux2_1 _25290_ (.A0(_06455_),
    .A1(_06960_),
    .S(net10655),
    .X(_06961_));
 sg13g2_nand2_2 _25291_ (.Y(_06962_),
    .A(net10660),
    .B(_06961_));
 sg13g2_xor2_1 _25292_ (.B(_06962_),
    .A(_06434_),
    .X(_06963_));
 sg13g2_nand2_1 _25293_ (.Y(_06964_),
    .A(net10731),
    .B(_06963_));
 sg13g2_o21ai_1 _25294_ (.B1(_06964_),
    .Y(_06965_),
    .A1(net10731),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[6] ));
 sg13g2_nor2_1 _25295_ (.A(net11003),
    .B(_06965_),
    .Y(_01891_));
 sg13g2_nand3_1 _25296_ (.B(_06434_),
    .C(_06455_),
    .A(net10362),
    .Y(_06966_));
 sg13g2_a21oi_1 _25297_ (.A1(_06432_),
    .A2(_06440_),
    .Y(_06967_),
    .B1(_06443_));
 sg13g2_xnor2_1 _25298_ (.Y(_06968_),
    .A(_04005_),
    .B(_06967_));
 sg13g2_nand2_1 _25299_ (.Y(_06969_),
    .A(net10656),
    .B(_06968_));
 sg13g2_a21o_1 _25300_ (.A2(_06969_),
    .A1(_06966_),
    .B1(net10379),
    .X(_06970_));
 sg13g2_xnor2_1 _25301_ (.Y(_06971_),
    .A(_06407_),
    .B(_06970_));
 sg13g2_nand2_1 _25302_ (.Y(_06972_),
    .A(net10726),
    .B(_06971_));
 sg13g2_o21ai_1 _25303_ (.B1(_06972_),
    .Y(_06973_),
    .A1(net10726),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[7] ));
 sg13g2_nor2_1 _25304_ (.A(net11003),
    .B(_06973_),
    .Y(_01892_));
 sg13g2_nor2_1 _25305_ (.A(_06444_),
    .B(_06491_),
    .Y(_06974_));
 sg13g2_xnor2_1 _25306_ (.Y(_06975_),
    .A(net10663),
    .B(_06974_));
 sg13g2_nor2_1 _25307_ (.A(net10656),
    .B(_06457_),
    .Y(_06976_));
 sg13g2_a21oi_1 _25308_ (.A1(net10656),
    .A2(_06975_),
    .Y(_06977_),
    .B1(_06976_));
 sg13g2_o21ai_1 _25309_ (.B1(_06402_),
    .Y(_06978_),
    .A1(net10379),
    .A2(_06977_));
 sg13g2_nand3b_1 _25310_ (.B(_06563_),
    .C(net10660),
    .Y(_06979_),
    .A_N(_06977_));
 sg13g2_nand3_1 _25311_ (.B(_06978_),
    .C(_06979_),
    .A(net10726),
    .Y(_06980_));
 sg13g2_o21ai_1 _25312_ (.B1(_06980_),
    .Y(_06981_),
    .A1(net10726),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[8] ));
 sg13g2_nor2_1 _25313_ (.A(net11004),
    .B(_06981_),
    .Y(_01893_));
 sg13g2_nor2_1 _25314_ (.A(_06404_),
    .B(_06446_),
    .Y(_06982_));
 sg13g2_xnor2_1 _25315_ (.Y(_06983_),
    .A(_04011_),
    .B(_06982_));
 sg13g2_nor2_1 _25316_ (.A(net10656),
    .B(_06458_),
    .Y(_06984_));
 sg13g2_a21oi_1 _25317_ (.A1(net10656),
    .A2(_06983_),
    .Y(_06985_),
    .B1(_06984_));
 sg13g2_nor2_1 _25318_ (.A(net10379),
    .B(_06985_),
    .Y(_06986_));
 sg13g2_xnor2_1 _25319_ (.Y(_06987_),
    .A(_06474_),
    .B(_06986_));
 sg13g2_o21ai_1 _25320_ (.B1(net11037),
    .Y(_06988_),
    .A1(net10726),
    .A2(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[9] ));
 sg13g2_a21oi_1 _25321_ (.A1(net10726),
    .A2(_06987_),
    .Y(_01894_),
    .B1(_06988_));
 sg13g2_nor2b_1 _25322_ (.A(net10728),
    .B_N(net10498),
    .Y(_06989_));
 sg13g2_a21oi_1 _25323_ (.A1(net10728),
    .A2(_06462_),
    .Y(_06990_),
    .B1(_06989_));
 sg13g2_nor2_1 _25324_ (.A(net11033),
    .B(_06990_),
    .Y(_01959_));
 sg13g2_buf_16 clkbuf_leaf_406_clk (.X(clknet_leaf_406_clk),
    .A(clknet_8_112_0_clk));
 sg13g2_nor2b_1 _25326_ (.A(net10727),
    .B_N(net10497),
    .Y(_06992_));
 sg13g2_a21oi_1 _25327_ (.A1(net10727),
    .A2(_06483_),
    .Y(_06993_),
    .B1(_06992_));
 sg13g2_nor2_1 _25328_ (.A(net11033),
    .B(_06993_),
    .Y(_01960_));
 sg13g2_nor2b_1 _25329_ (.A(net10727),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[12] ),
    .Y(_06994_));
 sg13g2_a21oi_1 _25330_ (.A1(net10727),
    .A2(_06489_),
    .Y(_06995_),
    .B1(_06994_));
 sg13g2_nor2_1 _25331_ (.A(net11033),
    .B(_06995_),
    .Y(_01961_));
 sg13g2_nor2b_1 _25332_ (.A(net10727),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[13] ),
    .Y(_06996_));
 sg13g2_a21oi_1 _25333_ (.A1(net10727),
    .A2(_06517_),
    .Y(_06997_),
    .B1(_06996_));
 sg13g2_nor2_1 _25334_ (.A(net11033),
    .B(_06997_),
    .Y(_01962_));
 sg13g2_nor2b_1 _25335_ (.A(net10727),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[14] ),
    .Y(_06998_));
 sg13g2_a21oi_1 _25336_ (.A1(net10727),
    .A2(_06533_),
    .Y(_06999_),
    .B1(_06998_));
 sg13g2_nor2_1 _25337_ (.A(net11034),
    .B(_06999_),
    .Y(_01963_));
 sg13g2_nor2b_1 _25338_ (.A(net10724),
    .B_N(net10496),
    .Y(_07000_));
 sg13g2_a21oi_1 _25339_ (.A1(net10724),
    .A2(net10257),
    .Y(_07001_),
    .B1(_07000_));
 sg13g2_nor2_2 _25340_ (.A(net11034),
    .B(_07001_),
    .Y(_01964_));
 sg13g2_buf_16 clkbuf_leaf_404_clk (.X(clknet_leaf_404_clk),
    .A(clknet_8_114_0_clk));
 sg13g2_nor2b_1 _25342_ (.A(net10724),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[16] ),
    .Y(_07003_));
 sg13g2_a21oi_1 _25343_ (.A1(net10724),
    .A2(_06592_),
    .Y(_07004_),
    .B1(_07003_));
 sg13g2_nor2_1 _25344_ (.A(net11034),
    .B(_07004_),
    .Y(_01965_));
 sg13g2_nor2b_1 _25345_ (.A(net10724),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[17] ),
    .Y(_07005_));
 sg13g2_a21oi_1 _25346_ (.A1(net10724),
    .A2(_06604_),
    .Y(_07006_),
    .B1(_07005_));
 sg13g2_nor2_1 _25347_ (.A(net11034),
    .B(_07006_),
    .Y(_01966_));
 sg13g2_nand2_1 _25348_ (.Y(_07007_),
    .A(_09847_),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[18] ));
 sg13g2_a21oi_1 _25349_ (.A1(_06627_),
    .A2(_07007_),
    .Y(_01967_),
    .B1(net11019));
 sg13g2_buf_16 clkbuf_leaf_403_clk (.X(clknet_leaf_403_clk),
    .A(clknet_8_114_0_clk));
 sg13g2_nor2b_1 _25351_ (.A(net10718),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[19] ),
    .Y(_07009_));
 sg13g2_a21oi_1 _25352_ (.A1(net10718),
    .A2(_06673_),
    .Y(_07010_),
    .B1(_07009_));
 sg13g2_nor2_1 _25353_ (.A(net11035),
    .B(_07010_),
    .Y(_01968_));
 sg13g2_nor2b_1 _25354_ (.A(net10731),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[1] ),
    .Y(_07011_));
 sg13g2_a21oi_1 _25355_ (.A1(net10731),
    .A2(_06411_),
    .Y(_07012_),
    .B1(_07011_));
 sg13g2_nor2_1 _25356_ (.A(net11003),
    .B(_07012_),
    .Y(_01969_));
 sg13g2_nor2b_1 _25357_ (.A(net10717),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[20] ),
    .Y(_07013_));
 sg13g2_a21oi_1 _25358_ (.A1(net10717),
    .A2(_06688_),
    .Y(_07014_),
    .B1(_07013_));
 sg13g2_nor2_1 _25359_ (.A(net11035),
    .B(_07014_),
    .Y(_01970_));
 sg13g2_buf_2 place9683 (.A(_03959_),
    .X(net9683));
 sg13g2_nor2b_1 _25361_ (.A(net10717),
    .B_N(net10495),
    .Y(_07016_));
 sg13g2_a21oi_1 _25362_ (.A1(net10717),
    .A2(_06705_),
    .Y(_07017_),
    .B1(_07016_));
 sg13g2_nor2_1 _25363_ (.A(net11035),
    .B(_07017_),
    .Y(_01971_));
 sg13g2_nor2b_1 _25364_ (.A(net10717),
    .B_N(net10494),
    .Y(_07018_));
 sg13g2_a21oi_1 _25365_ (.A1(net10717),
    .A2(net10195),
    .Y(_07019_),
    .B1(_07018_));
 sg13g2_nor2_1 _25366_ (.A(net11035),
    .B(_07019_),
    .Y(_01972_));
 sg13g2_nor2b_1 _25367_ (.A(net10718),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[23] ),
    .Y(_07020_));
 sg13g2_a21oi_1 _25368_ (.A1(net10718),
    .A2(_06763_),
    .Y(_07021_),
    .B1(_07020_));
 sg13g2_nor2_1 _25369_ (.A(net11035),
    .B(_07021_),
    .Y(_01973_));
 sg13g2_mux2_1 _25370_ (.A0(_09993_),
    .A1(_06758_),
    .S(net10718),
    .X(_07022_));
 sg13g2_nor2_1 _25371_ (.A(net11036),
    .B(_07022_),
    .Y(_01974_));
 sg13g2_nand2_1 _25372_ (.Y(_07023_),
    .A(net10382),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[25] ));
 sg13g2_a21oi_1 _25373_ (.A1(_06785_),
    .A2(_07023_),
    .Y(_01975_),
    .B1(net11036));
 sg13g2_nor2b_1 _25374_ (.A(net10718),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[26] ),
    .Y(_07024_));
 sg13g2_a21oi_1 _25375_ (.A1(net10718),
    .A2(_06819_),
    .Y(_07025_),
    .B1(_07024_));
 sg13g2_nor2_1 _25376_ (.A(net11036),
    .B(_07025_),
    .Y(_01976_));
 sg13g2_buf_2 place10945 (.A(net10944),
    .X(net10945));
 sg13g2_nor2b_1 _25378_ (.A(net10720),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[27] ),
    .Y(_07027_));
 sg13g2_a21oi_1 _25379_ (.A1(net10720),
    .A2(net10193),
    .Y(_07028_),
    .B1(_07027_));
 sg13g2_nor2_1 _25380_ (.A(net11036),
    .B(_07028_),
    .Y(_01977_));
 sg13g2_nor2_1 _25381_ (.A(net10720),
    .B(_10029_),
    .Y(_07029_));
 sg13g2_a21oi_1 _25382_ (.A1(net10720),
    .A2(_06847_),
    .Y(_07030_),
    .B1(_07029_));
 sg13g2_nor2_1 _25383_ (.A(net11036),
    .B(_07030_),
    .Y(_01978_));
 sg13g2_nor2b_1 _25384_ (.A(net10720),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[29] ),
    .Y(_07031_));
 sg13g2_a21oi_1 _25385_ (.A1(net10720),
    .A2(_06866_),
    .Y(_07032_),
    .B1(_07031_));
 sg13g2_nor2_1 _25386_ (.A(net11036),
    .B(_07032_),
    .Y(_01979_));
 sg13g2_nor2b_1 _25387_ (.A(net10729),
    .B_N(net10491),
    .Y(_07033_));
 sg13g2_a21oi_1 _25388_ (.A1(net10729),
    .A2(_06408_),
    .Y(_07034_),
    .B1(_07033_));
 sg13g2_nor2_1 _25389_ (.A(net11032),
    .B(_07034_),
    .Y(_01980_));
 sg13g2_nor2b_1 _25390_ (.A(net10720),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[30] ),
    .Y(_07035_));
 sg13g2_a21oi_1 _25391_ (.A1(net10719),
    .A2(_06911_),
    .Y(_07036_),
    .B1(_07035_));
 sg13g2_nor2_1 _25392_ (.A(net11036),
    .B(_07036_),
    .Y(_01981_));
 sg13g2_nand2_1 _25393_ (.Y(_07037_),
    .A(net10382),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[31] ));
 sg13g2_o21ai_1 _25394_ (.B1(_07037_),
    .Y(_07038_),
    .A1(net10382),
    .A2(_06917_));
 sg13g2_and2_1 _25395_ (.A(net11054),
    .B(_07038_),
    .X(_01982_));
 sg13g2_nor2b_1 _25396_ (.A(net10729),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[3] ),
    .Y(_07039_));
 sg13g2_a21oi_1 _25397_ (.A1(net10729),
    .A2(net10258),
    .Y(_07040_),
    .B1(_07039_));
 sg13g2_nor2_1 _25398_ (.A(net11032),
    .B(_07040_),
    .Y(_01983_));
 sg13g2_nand2_1 _25399_ (.Y(_07041_),
    .A(net10729),
    .B(_06421_));
 sg13g2_nand2_1 _25400_ (.Y(_07042_),
    .A(net10383),
    .B(\u_ac_controller_soc_inst.u_picorv32.reg_pc[4] ));
 sg13g2_a21oi_1 _25401_ (.A1(_07041_),
    .A2(_07042_),
    .Y(_01984_),
    .B1(net11032));
 sg13g2_nor2b_1 _25402_ (.A(net10729),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[5] ),
    .Y(_07043_));
 sg13g2_a21oi_1 _25403_ (.A1(net10725),
    .A2(_06437_),
    .Y(_07044_),
    .B1(_07043_));
 sg13g2_nor2_1 _25404_ (.A(net11032),
    .B(_07044_),
    .Y(_01985_));
 sg13g2_nor2_1 _25405_ (.A(net10729),
    .B(_09285_),
    .Y(_07045_));
 sg13g2_a21oi_1 _25406_ (.A1(net10729),
    .A2(_06434_),
    .Y(_07046_),
    .B1(_07045_));
 sg13g2_nor2_1 _25407_ (.A(net11032),
    .B(_07046_),
    .Y(_01986_));
 sg13g2_nor2_1 _25408_ (.A(net10728),
    .B(_09861_),
    .Y(_07047_));
 sg13g2_a21oi_1 _25409_ (.A1(net10728),
    .A2(_06405_),
    .Y(_07048_),
    .B1(_07047_));
 sg13g2_nor2_1 _25410_ (.A(net11033),
    .B(_07048_),
    .Y(_01987_));
 sg13g2_nor2b_1 _25411_ (.A(net10728),
    .B_N(net10488),
    .Y(_07049_));
 sg13g2_a21oi_1 _25412_ (.A1(net10728),
    .A2(_06402_),
    .Y(_07050_),
    .B1(_07049_));
 sg13g2_nor2_1 _25413_ (.A(net11032),
    .B(_07050_),
    .Y(_01988_));
 sg13g2_buf_2 place10896 (.A(net10894),
    .X(net10896));
 sg13g2_nor2b_1 _25415_ (.A(net10728),
    .B_N(\u_ac_controller_soc_inst.u_picorv32.reg_pc[9] ),
    .Y(_07052_));
 sg13g2_a21oi_1 _25416_ (.A1(net10728),
    .A2(_06474_),
    .Y(_07053_),
    .B1(_07052_));
 sg13g2_nor2_1 _25417_ (.A(net11033),
    .B(_07053_),
    .Y(_01989_));
 sg13g2_and2_1 _25418_ (.A(net11050),
    .B(\u_ac_controller_soc_inst.u_picorv32.cpu_state[0] ),
    .X(_01992_));
 sg13g2_nor4_2 _25419_ (.A(_07744_),
    .B(_07890_),
    .C(_07892_),
    .Y(_07054_),
    .D(_04552_));
 sg13g2_buf_2 place10882 (.A(_00008_),
    .X(net10882));
 sg13g2_nand2b_2 _25421_ (.Y(_07056_),
    .B(net9986),
    .A_N(_00106_));
 sg13g2_buf_16 clkbuf_leaf_411_clk (.X(clknet_leaf_411_clk),
    .A(clknet_8_100_0_clk));
 sg13g2_nor2b_2 _25423_ (.A(_00106_),
    .B_N(_07054_),
    .Y(_07058_));
 sg13g2_buf_2 place9692 (.A(net9691),
    .X(net9692));
 sg13g2_and3_2 _25425_ (.X(_07060_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[4] ),
    .B(net10298),
    .C(_07058_));
 sg13g2_a21oi_1 _25426_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.config_clk ),
    .A2(_07056_),
    .Y(_07061_),
    .B1(_07060_));
 sg13g2_nor2_1 _25427_ (.A(net10978),
    .B(_07061_),
    .Y(_02017_));
 sg13g2_buf_2 place9774 (.A(net9773),
    .X(net9774));
 sg13g2_nand3_1 _25429_ (.B(\u_ac_controller_soc_inst.cbus_wdata[20] ),
    .C(net9986),
    .A(net10600),
    .Y(_07063_));
 sg13g2_nand2_2 _25430_ (.Y(_07064_),
    .A(net10600),
    .B(net9986));
 sg13g2_buf_2 place9685 (.A(net9684),
    .X(net9685));
 sg13g2_nand2_1 _25432_ (.Y(_07066_),
    .A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[20] ),
    .B(_07064_));
 sg13g2_a21oi_1 _25433_ (.A1(_07063_),
    .A2(_07066_),
    .Y(_02018_),
    .B1(net10976));
 sg13g2_and3_2 _25434_ (.X(_07067_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[5] ),
    .B(net10298),
    .C(_07058_));
 sg13g2_a21oi_1 _25435_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.config_csb ),
    .A2(_07056_),
    .Y(_07068_),
    .B1(_07067_));
 sg13g2_nor2_1 _25436_ (.A(net10978),
    .B(_07068_),
    .Y(_02019_));
 sg13g2_nand3_1 _25437_ (.B(\u_ac_controller_soc_inst.cbus_wdata[22] ),
    .C(net9986),
    .A(net10600),
    .Y(_07069_));
 sg13g2_nand2_1 _25438_ (.Y(_07070_),
    .A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[22] ),
    .B(_07064_));
 sg13g2_a21oi_1 _25439_ (.A1(_07069_),
    .A2(_07070_),
    .Y(_02020_),
    .B1(net10977));
 sg13g2_and3_2 _25440_ (.X(_07071_),
    .A(net10605),
    .B(net10298),
    .C(_07058_));
 sg13g2_a21oi_1 _25441_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[0] ),
    .A2(_07056_),
    .Y(_07072_),
    .B1(_07071_));
 sg13g2_nor2_1 _25442_ (.A(net10978),
    .B(_07072_),
    .Y(_02021_));
 sg13g2_and3_2 _25443_ (.X(_07073_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[1] ),
    .B(net10298),
    .C(_07058_));
 sg13g2_a21oi_1 _25444_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[1] ),
    .A2(_07056_),
    .Y(_07074_),
    .B1(_07073_));
 sg13g2_nor2_1 _25445_ (.A(net10978),
    .B(_07074_),
    .Y(_02022_));
 sg13g2_and3_2 _25446_ (.X(_07075_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[2] ),
    .B(net10297),
    .C(_07058_));
 sg13g2_a21oi_1 _25447_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[2] ),
    .A2(_07056_),
    .Y(_07076_),
    .B1(_07075_));
 sg13g2_nor2_1 _25448_ (.A(net10977),
    .B(_07076_),
    .Y(_02023_));
 sg13g2_and3_2 _25449_ (.X(_07077_),
    .A(\u_ac_controller_soc_inst.cbus_wdata[3] ),
    .B(net10297),
    .C(_07058_));
 sg13g2_a21oi_1 _25450_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[3] ),
    .A2(_07056_),
    .Y(_07078_),
    .B1(_07077_));
 sg13g2_nor2_1 _25451_ (.A(net10977),
    .B(_07078_),
    .Y(_02024_));
 sg13g2_nand3_1 _25452_ (.B(\u_ac_controller_soc_inst.cbus_wdata[16] ),
    .C(net9986),
    .A(net10600),
    .Y(_07079_));
 sg13g2_nand2_1 _25453_ (.Y(_07080_),
    .A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[16] ),
    .B(_07064_));
 sg13g2_a21oi_1 _25454_ (.A1(_07079_),
    .A2(_07080_),
    .Y(_02025_),
    .B1(net10977));
 sg13g2_nand3_1 _25455_ (.B(\u_ac_controller_soc_inst.cbus_wdata[17] ),
    .C(net9986),
    .A(net10600),
    .Y(_07081_));
 sg13g2_nand2_1 _25456_ (.Y(_07082_),
    .A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[17] ),
    .B(_07064_));
 sg13g2_a21oi_1 _25457_ (.A1(_07081_),
    .A2(_07082_),
    .Y(_02026_),
    .B1(net10977));
 sg13g2_nand3_1 _25458_ (.B(\u_ac_controller_soc_inst.cbus_wdata[18] ),
    .C(net9986),
    .A(net10600),
    .Y(_07083_));
 sg13g2_nand2_1 _25459_ (.Y(_07084_),
    .A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[18] ),
    .B(_07064_));
 sg13g2_a21oi_1 _25460_ (.A1(_07083_),
    .A2(_07084_),
    .Y(_02027_),
    .B1(net10976));
 sg13g2_nand2_1 _25461_ (.Y(_07085_),
    .A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[19] ),
    .B(_07064_));
 sg13g2_nand3_1 _25462_ (.B(\u_ac_controller_soc_inst.cbus_wdata[19] ),
    .C(_07054_),
    .A(net10600),
    .Y(_07086_));
 sg13g2_nand3_1 _25463_ (.B(_07085_),
    .C(_07086_),
    .A(net11041),
    .Y(_02028_));
 sg13g2_a21oi_1 _25464_ (.A1(\u_ac_controller_soc_inst.cbus_wstrb[3] ),
    .A2(_07054_),
    .Y(_07087_),
    .B1(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[31] ));
 sg13g2_nand2_1 _25465_ (.Y(_07088_),
    .A(\u_ac_controller_soc_inst.cbus_wstrb[3] ),
    .B(_07054_));
 sg13g2_a21oi_1 _25466_ (.A1(\u_ac_controller_soc_inst.cbus_wdata[31] ),
    .A2(net10298),
    .Y(_07089_),
    .B1(_07088_));
 sg13g2_o21ai_1 _25467_ (.B1(net11041),
    .Y(_02029_),
    .A1(_07087_),
    .A2(_07089_));
 sg13g2_nand2_2 _25468_ (.Y(_07090_),
    .A(\u_ac_controller_soc_inst.cbus_wstrb[1] ),
    .B(_07054_));
 sg13g2_buf_2 place9690 (.A(_09988_),
    .X(net9690));
 sg13g2_nor3_1 _25470_ (.A(_05878_),
    .B(net10302),
    .C(_07090_),
    .Y(_07092_));
 sg13g2_a21oi_1 _25471_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[0] ),
    .A2(_07090_),
    .Y(_07093_),
    .B1(_07092_));
 sg13g2_nor2_1 _25472_ (.A(net10978),
    .B(_07093_),
    .Y(_02030_));
 sg13g2_nor3_1 _25473_ (.A(_05881_),
    .B(net10302),
    .C(_07090_),
    .Y(_07094_));
 sg13g2_a21oi_1 _25474_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[1] ),
    .A2(_07090_),
    .Y(_07095_),
    .B1(_07094_));
 sg13g2_nor2_1 _25475_ (.A(net10978),
    .B(_07095_),
    .Y(_02031_));
 sg13g2_nor3_1 _25476_ (.A(_05840_),
    .B(net10302),
    .C(_07090_),
    .Y(_07096_));
 sg13g2_a21oi_1 _25477_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[2] ),
    .A2(_07090_),
    .Y(_07097_),
    .B1(_07096_));
 sg13g2_nor2_1 _25478_ (.A(net10977),
    .B(_07097_),
    .Y(_02032_));
 sg13g2_nor3_1 _25479_ (.A(_05843_),
    .B(net10302),
    .C(_07090_),
    .Y(_07098_));
 sg13g2_a21oi_1 _25480_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[3] ),
    .A2(_07090_),
    .Y(_07099_),
    .B1(_07098_));
 sg13g2_nor2_1 _25481_ (.A(net10978),
    .B(_07099_),
    .Y(_02033_));
 sg13g2_nand3_1 _25482_ (.B(\u_ac_controller_soc_inst.cbus_wdata[21] ),
    .C(net9986),
    .A(net10600),
    .Y(_07100_));
 sg13g2_nand2_1 _25483_ (.Y(_07101_),
    .A(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[21] ),
    .B(_07064_));
 sg13g2_a21oi_1 _25484_ (.A1(_07100_),
    .A2(_07101_),
    .Y(_02034_),
    .B1(net10976));
 sg13g2_nand2_1 _25485_ (.Y(_07102_),
    .A(_04802_),
    .B(_07054_));
 sg13g2_nand3b_1 _25486_ (.B(_07102_),
    .C(net11041),
    .Y(_02107_),
    .A_N(_00120_));
 sg13g2_nand2_1 _25487_ (.Y(_07103_),
    .A(_00093_),
    .B(_08163_));
 sg13g2_xnor2_1 _25488_ (.Y(_07104_),
    .A(_00092_),
    .B(_07103_));
 sg13g2_nand2b_1 _25489_ (.Y(_07105_),
    .B(net10260),
    .A_N(_08177_));
 sg13g2_nand2b_1 _25490_ (.Y(_07106_),
    .B(net10457),
    .A_N(_08190_));
 sg13g2_nand3_1 _25491_ (.B(_07105_),
    .C(_07106_),
    .A(_00092_),
    .Y(_07107_));
 sg13g2_a22oi_1 _25492_ (.Y(_07108_),
    .B1(net10260),
    .B2(_08177_),
    .A2(net10457),
    .A1(_08190_));
 sg13g2_nand2b_1 _25493_ (.Y(_07109_),
    .B(_07108_),
    .A_N(_00092_));
 sg13g2_a221oi_1 _25494_ (.B2(_07109_),
    .C1(_04779_),
    .B1(_07107_),
    .A1(net10464),
    .Y(_07110_),
    .A2(_07104_));
 sg13g2_a21oi_1 _25495_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[3] ),
    .A2(_04779_),
    .Y(_07111_),
    .B1(_07110_));
 sg13g2_a21o_1 _25496_ (.A2(_07111_),
    .A1(_08221_),
    .B1(_08220_),
    .X(_07112_));
 sg13g2_inv_1 _25497_ (.Y(_02111_),
    .A(_07112_));
 sg13g2_and2_1 _25498_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_rd ),
    .B(net9747),
    .X(_07113_));
 sg13g2_buf_2 place9687 (.A(net9686),
    .X(net9687));
 sg13g2_xor2_1 _25500_ (.B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk ),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[0] ),
    .X(_07115_));
 sg13g2_a22oi_1 _25501_ (.Y(_07116_),
    .B1(_07115_),
    .B2(_08204_),
    .A2(_07113_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[0] ));
 sg13g2_nor2_1 _25502_ (.A(_08220_),
    .B(_07116_),
    .Y(_02112_));
 sg13g2_nand2b_1 _25503_ (.Y(_07117_),
    .B(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk ),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[0] ));
 sg13g2_xnor2_1 _25504_ (.Y(_07118_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[1] ),
    .B(_07117_));
 sg13g2_a22oi_1 _25505_ (.Y(_07119_),
    .B1(_07118_),
    .B2(_08204_),
    .A2(_07113_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[1] ));
 sg13g2_nor2_1 _25506_ (.A(_08220_),
    .B(_07119_),
    .Y(_02113_));
 sg13g2_nor2_1 _25507_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[1] ),
    .B(_07117_),
    .Y(_07120_));
 sg13g2_xor2_1 _25508_ (.B(_07120_),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[2] ),
    .X(_07121_));
 sg13g2_a22oi_1 _25509_ (.Y(_07122_),
    .B1(_07121_),
    .B2(_08204_),
    .A2(_07113_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[2] ));
 sg13g2_nor2_1 _25510_ (.A(_08220_),
    .B(_07122_),
    .Y(_02114_));
 sg13g2_nand2b_1 _25511_ (.Y(_07123_),
    .B(_07120_),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[2] ));
 sg13g2_a22oi_1 _25512_ (.Y(_07124_),
    .B1(_07123_),
    .B2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[3] ),
    .A2(_07113_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[3] ));
 sg13g2_nor2_1 _25513_ (.A(_08220_),
    .B(_07124_),
    .Y(_02115_));
 sg13g2_nand2b_1 _25514_ (.Y(_02116_),
    .B(net10461),
    .A_N(_08206_));
 sg13g2_a21o_1 _25515_ (.A2(_08221_),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_csb ),
    .B1(_08220_),
    .X(_02118_));
 sg13g2_nand3b_1 _25516_ (.B(net10466),
    .C(net10461),
    .Y(_02127_),
    .A_N(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.fetch ));
 sg13g2_nand2_1 _25517_ (.Y(_07125_),
    .A(net10466),
    .B(_08221_));
 sg13g2_nand3_1 _25518_ (.B(\u_ac_controller_soc_inst.u_spi_flash_mem.din_qspi ),
    .C(net9747),
    .A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_ddr ),
    .Y(_07126_));
 sg13g2_a21oi_1 _25519_ (.A1(_07125_),
    .A2(_07126_),
    .Y(_02136_),
    .B1(_08220_));
 sg13g2_nor2b_1 _25520_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.din_qspi ),
    .B_N(\u_ac_controller_soc_inst.u_spi_flash_mem.din_ddr ),
    .Y(_07127_));
 sg13g2_mux2_1 _25521_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi ),
    .A1(_07127_),
    .S(net9747),
    .X(_07128_));
 sg13g2_and2_1 _25522_ (.A(net10461),
    .B(_07128_),
    .X(_02137_));
 sg13g2_mux2_1 _25523_ (.A0(net10462),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_qspi ),
    .S(net9747),
    .X(_07129_));
 sg13g2_and2_1 _25524_ (.A(net10461),
    .B(_07129_),
    .X(_02138_));
 sg13g2_a21oi_1 _25525_ (.A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_rd ),
    .A2(_08221_),
    .Y(_07130_),
    .B1(_07113_));
 sg13g2_nor2b_1 _25526_ (.A(_07130_),
    .B_N(net10461),
    .Y(_02139_));
 sg13g2_mux2_1 _25527_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[0] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[0] ),
    .S(_08207_),
    .X(_07131_));
 sg13g2_and2_1 _25528_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.resetn ),
    .B(_07131_),
    .X(_02140_));
 sg13g2_mux2_1 _25529_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[1] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[1] ),
    .S(_08207_),
    .X(_07132_));
 sg13g2_and2_1 _25530_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.resetn ),
    .B(_07132_),
    .X(_02141_));
 sg13g2_mux2_1 _25531_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[2] ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[2] ),
    .S(_08207_),
    .X(_07133_));
 sg13g2_and2_1 _25532_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.resetn ),
    .B(_07133_),
    .X(_02142_));
 sg13g2_nor2b_2 _25533_ (.A(net10487),
    .B_N(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io0_do ),
    .Y(_07134_));
 sg13g2_a21oi_2 _25534_ (.B1(_07134_),
    .Y(_07135_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io0_90 ),
    .A1(net10487));
 sg13g2_nor2_1 _25535_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[0] ),
    .B(net10486),
    .Y(_07136_));
 sg13g2_a21oi_2 _25536_ (.B1(_07136_),
    .Y(spi_flash_io0_do),
    .A2(_07135_),
    .A1(net10486));
 sg13g2_nor3_1 _25537_ (.A(net10487),
    .B(_08564_),
    .C(_08567_),
    .Y(_07137_));
 sg13g2_a21oi_2 _25538_ (.B1(_07137_),
    .Y(_07138_),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io1_90 ),
    .A1(net10487));
 sg13g2_nor2_1 _25539_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[1] ),
    .B(net10486),
    .Y(_07139_));
 sg13g2_a21oi_2 _25540_ (.B1(_07139_),
    .Y(spi_flash_io1_do),
    .A2(_07138_),
    .A1(net10486));
 sg13g2_mux2_1 _25541_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io2_do ),
    .A1(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io2_90 ),
    .S(net10487),
    .X(_07140_));
 sg13g2_mux2_1 _25542_ (.A0(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[2] ),
    .A1(_07140_),
    .S(net10485),
    .X(spi_flash_io2_do));
 sg13g2_nor3_1 _25543_ (.A(net10487),
    .B(_00124_),
    .C(_08569_),
    .Y(_07141_));
 sg13g2_a21oi_1 _25544_ (.A1(net10487),
    .A2(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io3_90 ),
    .Y(_07142_),
    .B1(_07141_));
 sg13g2_nor2_1 _25545_ (.A(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[3] ),
    .B(net10485),
    .Y(_07143_));
 sg13g2_a21oi_2 _25546_ (.B1(_07143_),
    .Y(spi_flash_io3_do),
    .A2(_07142_),
    .A1(net10485));
 sg13g2_a21oi_1 _25547_ (.A1(_07886_),
    .A2(_04554_),
    .Y(_07144_),
    .B1(_05425_));
 sg13g2_nor2b_2 _25548_ (.A(_07144_),
    .B_N(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[39] ),
    .Y(spi_sensor_mosi));
 sg13g2_nor2_1 _25549_ (.A(_00138_),
    .B(_08865_),
    .Y(_07145_));
 sg13g2_buf_2 place9689 (.A(_09988_),
    .X(net9689));
 sg13g2_buf_2 place9783 (.A(net9782),
    .X(net9783));
 sg13g2_or2_1 _25552_ (.X(_07148_),
    .B(\u_ac_controller_soc_inst.u_picorv32.instr_xori ),
    .A(\u_ac_controller_soc_inst.u_picorv32.instr_xor ));
 sg13g2_buf_2 place9782 (.A(net9781),
    .X(net9782));
 sg13g2_a21oi_2 _25554_ (.B1(net10306),
    .Y(_07150_),
    .A2(net10447),
    .A1(_00138_));
 sg13g2_mux2_1 _25555_ (.A0(net10448),
    .A1(_07150_),
    .S(_08845_),
    .X(_07151_));
 sg13g2_a21oi_2 _25556_ (.B1(_08844_),
    .Y(_07152_),
    .A2(_07151_),
    .A1(net10453));
 sg13g2_a21o_1 _25557_ (.A2(_07145_),
    .A1(_08859_),
    .B1(_07152_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[0] ));
 sg13g2_and3_2 _25558_ (.X(_07153_),
    .A(_00138_),
    .B(_08295_),
    .C(_08297_));
 sg13g2_buf_2 place10881 (.A(_00008_),
    .X(net10881));
 sg13g2_buf_2 place10732 (.A(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[0] ),
    .X(net10732));
 sg13g2_buf_2 place9772 (.A(_04955_),
    .X(net9772));
 sg13g2_nor2_1 _25562_ (.A(net10500),
    .B(net10523),
    .Y(_07157_));
 sg13g2_a22oi_1 _25563_ (.Y(_07158_),
    .B1(net10500),
    .B2(net10523),
    .A2(net10524),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[7] ));
 sg13g2_nor2_2 _25564_ (.A(_07157_),
    .B(_07158_),
    .Y(_07159_));
 sg13g2_nor3_1 _25565_ (.A(net10531),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[2] ),
    .C(net10539),
    .Y(_07160_));
 sg13g2_nor3_1 _25566_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[3] ),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[2] ),
    .C(net10539),
    .Y(_07161_));
 sg13g2_nor2_1 _25567_ (.A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[3] ),
    .B(net10531),
    .Y(_07162_));
 sg13g2_or3_1 _25568_ (.A(_07160_),
    .B(_07161_),
    .C(_07162_),
    .X(_07163_));
 sg13g2_buf_2 place9773 (.A(net9772),
    .X(net9773));
 sg13g2_a21o_1 _25570_ (.A2(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[0] ),
    .A1(net10599),
    .B1(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[1] ),
    .X(_07165_));
 sg13g2_a21o_1 _25571_ (.A2(net10539),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[2] ),
    .B1(net10532),
    .X(_07166_));
 sg13g2_a21o_1 _25572_ (.A2(net10539),
    .A1(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[2] ),
    .B1(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[3] ),
    .X(_07167_));
 sg13g2_and3_1 _25573_ (.X(_07168_),
    .A(net10599),
    .B(net10520),
    .C(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[1] ));
 sg13g2_a221oi_1 _25574_ (.B2(_07167_),
    .C1(_07168_),
    .B1(_07166_),
    .A1(net10572),
    .Y(_07169_),
    .A2(_07165_));
 sg13g2_buf_2 place9680 (.A(_10005_),
    .X(net9680));
 sg13g2_and2_1 _25576_ (.A(net10502),
    .B(net10527),
    .X(_07171_));
 sg13g2_buf_2 place9765 (.A(net9764),
    .X(net9765));
 sg13g2_nor3_1 _25578_ (.A(net10503),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[4] ),
    .C(_07171_),
    .Y(_07173_));
 sg13g2_o21ai_1 _25579_ (.B1(_07173_),
    .Y(_07174_),
    .A1(_07163_),
    .A2(_07169_));
 sg13g2_nor3_1 _25580_ (.A(net10529),
    .B(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[4] ),
    .C(_07171_),
    .Y(_07175_));
 sg13g2_o21ai_1 _25581_ (.B1(_07175_),
    .Y(_07176_),
    .A1(_07163_),
    .A2(_07169_));
 sg13g2_nor3_1 _25582_ (.A(net10529),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[4] ),
    .C(_07171_),
    .Y(_07177_));
 sg13g2_o21ai_1 _25583_ (.B1(_07177_),
    .Y(_07178_),
    .A1(_07163_),
    .A2(_07169_));
 sg13g2_or2_1 _25584_ (.X(_07179_),
    .B(net10527),
    .A(net10502));
 sg13g2_nand4_1 _25585_ (.B(_07176_),
    .C(_07178_),
    .A(_07174_),
    .Y(_07180_),
    .D(_07179_));
 sg13g2_o21ai_1 _25586_ (.B1(_08701_),
    .Y(_07181_),
    .A1(_07173_),
    .A2(_07175_));
 sg13g2_nor2_1 _25587_ (.A(net10503),
    .B(net10529),
    .Y(_07182_));
 sg13g2_nand2b_1 _25588_ (.Y(_07183_),
    .B(_07182_),
    .A_N(_07171_));
 sg13g2_nor3_1 _25589_ (.A(net10503),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[4] ),
    .C(_07171_),
    .Y(_07184_));
 sg13g2_o21ai_1 _25590_ (.B1(_07184_),
    .Y(_07185_),
    .A1(_07163_),
    .A2(_07169_));
 sg13g2_nand3_1 _25591_ (.B(_07183_),
    .C(_07185_),
    .A(_07181_),
    .Y(_07186_));
 sg13g2_a21oi_1 _25592_ (.A1(_03677_),
    .A2(_08716_),
    .Y(_07187_),
    .B1(_07157_));
 sg13g2_inv_1 _25593_ (.Y(_07188_),
    .A(_07187_));
 sg13g2_nor3_2 _25594_ (.A(_07180_),
    .B(_07186_),
    .C(_07188_),
    .Y(_07189_));
 sg13g2_o21ai_1 _25595_ (.B1(net10521),
    .Y(_07190_),
    .A1(_07159_),
    .A2(_07189_));
 sg13g2_nor3_1 _25596_ (.A(net10521),
    .B(_07159_),
    .C(_07189_),
    .Y(_07191_));
 sg13g2_a21oi_2 _25597_ (.B1(_07191_),
    .Y(_07192_),
    .A2(_07190_),
    .A1(_08779_));
 sg13g2_inv_4 _25598_ (.A(net10633),
    .Y(_07193_));
 sg13g2_buf_2 place9790 (.A(net9788),
    .X(net9790));
 sg13g2_nor2_1 _25600_ (.A(_08779_),
    .B(net10521),
    .Y(_07195_));
 sg13g2_nand2_1 _25601_ (.Y(_07196_),
    .A(_08712_),
    .B(_08723_));
 sg13g2_or4_1 _25602_ (.A(_08698_),
    .B(_08706_),
    .C(_08776_),
    .D(_08777_),
    .X(_07197_));
 sg13g2_a22oi_1 _25603_ (.Y(_07198_),
    .B1(_07196_),
    .B2(_07197_),
    .A2(net10522),
    .A1(_08779_));
 sg13g2_or3_1 _25604_ (.A(net10304),
    .B(_07195_),
    .C(_07198_),
    .X(_07199_));
 sg13g2_o21ai_1 _25605_ (.B1(_07199_),
    .Y(_07200_),
    .A1(net10636),
    .A2(_07192_));
 sg13g2_xnor2_1 _25606_ (.Y(_07201_),
    .A(_08740_),
    .B(_07200_));
 sg13g2_buf_2 place9681 (.A(_10005_),
    .X(net9681));
 sg13g2_buf_2 place9768 (.A(net9766),
    .X(net9768));
 sg13g2_buf_2 place9676 (.A(net9675),
    .X(net9676));
 sg13g2_nand3_1 _25610_ (.B(net10594),
    .C(net10447),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[10] ),
    .Y(_07205_));
 sg13g2_o21ai_1 _25611_ (.B1(_07205_),
    .Y(_07206_),
    .A1(net10594),
    .A2(net10307));
 sg13g2_nand2_2 _25612_ (.Y(_07207_),
    .A(_08292_),
    .B(_08294_));
 sg13g2_buf_2 place9767 (.A(net9766),
    .X(net9767));
 sg13g2_buf_2 place9766 (.A(net9761),
    .X(net9766));
 sg13g2_nand2_1 _25615_ (.Y(_07210_),
    .A(net10594),
    .B(net10254));
 sg13g2_a22oi_1 _25616_ (.Y(_07211_),
    .B1(_07210_),
    .B2(_03279_),
    .A2(_07206_),
    .A1(net10453));
 sg13g2_a21o_1 _25617_ (.A2(_07201_),
    .A1(net10189),
    .B1(_07211_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[10] ));
 sg13g2_nor2_1 _25618_ (.A(net10594),
    .B(_07192_),
    .Y(_07212_));
 sg13g2_a21oi_1 _25619_ (.A1(net10594),
    .A2(_07192_),
    .Y(_07213_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[10] ));
 sg13g2_nor2_1 _25620_ (.A(_07212_),
    .B(_07213_),
    .Y(_07214_));
 sg13g2_nor3_1 _25621_ (.A(_12002_),
    .B(_07195_),
    .C(_07198_),
    .Y(_07215_));
 sg13g2_o21ai_1 _25622_ (.B1(_12002_),
    .Y(_07216_),
    .A1(_07195_),
    .A2(_07198_));
 sg13g2_nand2_1 _25623_ (.Y(_07217_),
    .A(_03279_),
    .B(_07216_));
 sg13g2_nand2b_1 _25624_ (.Y(_07218_),
    .B(_07217_),
    .A_N(_07215_));
 sg13g2_nand2_1 _25625_ (.Y(_07219_),
    .A(net10635),
    .B(_07218_));
 sg13g2_o21ai_1 _25626_ (.B1(_07219_),
    .Y(_07220_),
    .A1(net10635),
    .A2(_07214_));
 sg13g2_xnor2_1 _25627_ (.Y(_07221_),
    .A(_08743_),
    .B(_07220_));
 sg13g2_buf_2 place9781 (.A(net9780),
    .X(net9781));
 sg13g2_nand3_1 _25629_ (.B(net10592),
    .C(net10448),
    .A(net10519),
    .Y(_07223_));
 sg13g2_o21ai_1 _25630_ (.B1(_07223_),
    .Y(_07224_),
    .A1(net10592),
    .A2(net10307));
 sg13g2_buf_2 place9677 (.A(net9675),
    .X(net9677));
 sg13g2_a21oi_1 _25632_ (.A1(net10592),
    .A2(net10253),
    .Y(_07226_),
    .B1(net10519));
 sg13g2_a21oi_1 _25633_ (.A1(net10453),
    .A2(_07224_),
    .Y(_07227_),
    .B1(_07226_));
 sg13g2_a21o_1 _25634_ (.A2(_07221_),
    .A1(net10188),
    .B1(_07227_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[11] ));
 sg13g2_nand2_1 _25635_ (.Y(_07228_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[11] ),
    .B(_08754_));
 sg13g2_nand2_1 _25636_ (.Y(_07229_),
    .A(_07228_),
    .B(_07218_));
 sg13g2_o21ai_1 _25637_ (.B1(_07229_),
    .Y(_07230_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[11] ),
    .A2(_08754_));
 sg13g2_nor2_1 _25638_ (.A(net10519),
    .B(net10592),
    .Y(_07231_));
 sg13g2_nand2b_1 _25639_ (.Y(_07232_),
    .B(_07214_),
    .A_N(_07231_));
 sg13g2_buf_2 place9672 (.A(net9671),
    .X(net9672));
 sg13g2_a21oi_1 _25641_ (.A1(net10519),
    .A2(net10592),
    .Y(_07234_),
    .B1(net10635));
 sg13g2_a22oi_1 _25642_ (.Y(_07235_),
    .B1(_07232_),
    .B2(_07234_),
    .A2(_07230_),
    .A1(net10635));
 sg13g2_xor2_1 _25643_ (.B(_07235_),
    .A(_08746_),
    .X(_07236_));
 sg13g2_nand3_1 _25644_ (.B(net10589),
    .C(net10447),
    .A(net10518),
    .Y(_07237_));
 sg13g2_o21ai_1 _25645_ (.B1(_07237_),
    .Y(_07238_),
    .A1(net10589),
    .A2(net10307));
 sg13g2_nand2_1 _25646_ (.Y(_07239_),
    .A(net10589),
    .B(net10254));
 sg13g2_a22oi_1 _25647_ (.Y(_07240_),
    .B1(_07239_),
    .B2(_03352_),
    .A2(_07238_),
    .A1(net10453));
 sg13g2_a21o_2 _25648_ (.A2(_07236_),
    .A1(net10189),
    .B1(_07240_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[12] ));
 sg13g2_o21ai_1 _25649_ (.B1(_08758_),
    .Y(_07241_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[11] ),
    .A2(_08754_));
 sg13g2_o21ai_1 _25650_ (.B1(net10518),
    .Y(_07242_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[11] ),
    .A2(_08754_));
 sg13g2_a221oi_1 _25651_ (.B2(_07242_),
    .C1(_07215_),
    .B1(_07241_),
    .A1(_03279_),
    .Y(_07243_),
    .A2(_07216_));
 sg13g2_a21oi_1 _25652_ (.A1(_03352_),
    .A2(net10590),
    .Y(_07244_),
    .B1(_07228_));
 sg13g2_or3_1 _25653_ (.A(_08762_),
    .B(_07243_),
    .C(_07244_),
    .X(_07245_));
 sg13g2_buf_2 place9675 (.A(_10014_),
    .X(net9675));
 sg13g2_nor2_2 _25655_ (.A(_07159_),
    .B(_07189_),
    .Y(_07247_));
 sg13g2_nand4_1 _25656_ (.B(_08743_),
    .C(_08746_),
    .A(_08740_),
    .Y(_07248_),
    .D(_08830_));
 sg13g2_a21oi_1 _25657_ (.A1(net10499),
    .A2(net10521),
    .Y(_07249_),
    .B1(net10593));
 sg13g2_nand3_1 _25658_ (.B(net10499),
    .C(net10521),
    .A(net10593),
    .Y(_07250_));
 sg13g2_o21ai_1 _25659_ (.B1(_07250_),
    .Y(_07251_),
    .A1(_03279_),
    .A2(_07249_));
 sg13g2_a21oi_1 _25660_ (.A1(net10519),
    .A2(net10592),
    .Y(_07252_),
    .B1(_07251_));
 sg13g2_o21ai_1 _25661_ (.B1(_08758_),
    .Y(_07253_),
    .A1(_07231_),
    .A2(_07252_));
 sg13g2_nor3_1 _25662_ (.A(_08758_),
    .B(_07231_),
    .C(_07252_),
    .Y(_07254_));
 sg13g2_a21o_2 _25663_ (.A2(_07253_),
    .A1(net10518),
    .B1(_07254_),
    .X(_07255_));
 sg13g2_inv_1 _25664_ (.Y(_07256_),
    .A(_07255_));
 sg13g2_o21ai_1 _25665_ (.B1(_07256_),
    .Y(_07257_),
    .A1(_07247_),
    .A2(_07248_));
 sg13g2_buf_2 place9674 (.A(_10014_),
    .X(net9674));
 sg13g2_buf_2 place9686 (.A(net9685),
    .X(net9686));
 sg13g2_mux2_1 _25668_ (.A0(_07245_),
    .A1(_07257_),
    .S(net10304),
    .X(_07260_));
 sg13g2_xnor2_1 _25669_ (.Y(_07261_),
    .A(_08727_),
    .B(_07260_));
 sg13g2_buf_2 place9682 (.A(_06265_),
    .X(net9682));
 sg13g2_nand3_1 _25671_ (.B(net10587),
    .C(net10448),
    .A(net10517),
    .Y(_07263_));
 sg13g2_o21ai_1 _25672_ (.B1(_07263_),
    .Y(_07264_),
    .A1(net10587),
    .A2(net10307));
 sg13g2_nand2_1 _25673_ (.Y(_07265_),
    .A(net10587),
    .B(net10253));
 sg13g2_a22oi_1 _25674_ (.Y(_07266_),
    .B1(_07265_),
    .B2(_08752_),
    .A2(_07264_),
    .A1(net10453));
 sg13g2_a21o_1 _25675_ (.A2(_07261_),
    .A1(net10188),
    .B1(_07266_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[13] ));
 sg13g2_o21ai_1 _25676_ (.B1(net10517),
    .Y(_07267_),
    .A1(net10587),
    .A2(_07257_));
 sg13g2_inv_1 _25677_ (.Y(_07268_),
    .A(_07267_));
 sg13g2_a21oi_1 _25678_ (.A1(net10587),
    .A2(_07257_),
    .Y(_07269_),
    .B1(_07268_));
 sg13g2_nand2b_1 _25679_ (.Y(_07270_),
    .B(net10587),
    .A_N(_07245_));
 sg13g2_a21o_1 _25680_ (.A2(_07245_),
    .A1(_08761_),
    .B1(net10517),
    .X(_07271_));
 sg13g2_a21oi_1 _25681_ (.A1(_07270_),
    .A2(_07271_),
    .Y(_07272_),
    .B1(net10304));
 sg13g2_a21o_1 _25682_ (.A2(_07269_),
    .A1(net10304),
    .B1(_07272_),
    .X(_07273_));
 sg13g2_xor2_1 _25683_ (.B(_07273_),
    .A(_08733_),
    .X(_07274_));
 sg13g2_nand3_1 _25684_ (.B(net10585),
    .C(net10448),
    .A(net10516),
    .Y(_07275_));
 sg13g2_o21ai_1 _25685_ (.B1(_07275_),
    .Y(_07276_),
    .A1(net10585),
    .A2(net10307));
 sg13g2_a21oi_1 _25686_ (.A1(net10585),
    .A2(net10253),
    .Y(_07277_),
    .B1(net10516));
 sg13g2_a21oi_1 _25687_ (.A1(net10452),
    .A2(_07276_),
    .Y(_07278_),
    .B1(_07277_));
 sg13g2_a21o_1 _25688_ (.A2(_07274_),
    .A1(net10188),
    .B1(_07278_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[14] ));
 sg13g2_nand2_1 _25689_ (.Y(_07279_),
    .A(net10635),
    .B(_08730_));
 sg13g2_a22oi_1 _25690_ (.Y(_07280_),
    .B1(_07270_),
    .B2(_07271_),
    .A2(_02354_),
    .A1(net10516));
 sg13g2_a21o_1 _25691_ (.A2(net10586),
    .A1(net10517),
    .B1(net10585),
    .X(_07281_));
 sg13g2_nor2_1 _25692_ (.A(_08727_),
    .B(_08733_),
    .Y(_07282_));
 sg13g2_and3_1 _25693_ (.X(_07283_),
    .A(net10585),
    .B(net10517),
    .C(net10586));
 sg13g2_a221oi_1 _25694_ (.B2(_07257_),
    .C1(_07283_),
    .B1(_07282_),
    .A1(net10516),
    .Y(_07284_),
    .A2(_07281_));
 sg13g2_or2_1 _25695_ (.X(_07285_),
    .B(_07284_),
    .A(net10635));
 sg13g2_o21ai_1 _25696_ (.B1(_07285_),
    .Y(_07286_),
    .A1(_07279_),
    .A2(_07280_));
 sg13g2_xor2_1 _25697_ (.B(_07286_),
    .A(_08737_),
    .X(_07287_));
 sg13g2_buf_2 place9671 (.A(_11943_),
    .X(net9671));
 sg13g2_nand3_1 _25699_ (.B(net10583),
    .C(net10448),
    .A(net10515),
    .Y(_07289_));
 sg13g2_o21ai_1 _25700_ (.B1(_07289_),
    .Y(_07290_),
    .A1(net10583),
    .A2(net10307));
 sg13g2_nand2_1 _25701_ (.Y(_07291_),
    .A(net10583),
    .B(net10253));
 sg13g2_a22oi_1 _25702_ (.Y(_07292_),
    .B1(_07291_),
    .B2(_08770_),
    .A2(_07290_),
    .A1(net10452));
 sg13g2_a21o_1 _25703_ (.A2(_07287_),
    .A1(net10188),
    .B1(_07292_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[15] ));
 sg13g2_nand2_1 _25704_ (.Y(_07293_),
    .A(net10515),
    .B(net10583));
 sg13g2_nor2_1 _25705_ (.A(net10515),
    .B(net10583),
    .Y(_07294_));
 sg13g2_a21oi_2 _25706_ (.B1(_07294_),
    .Y(_07295_),
    .A2(_07293_),
    .A1(_07284_));
 sg13g2_nand2_1 _25707_ (.Y(_07296_),
    .A(net10635),
    .B(_08784_));
 sg13g2_o21ai_1 _25708_ (.B1(_07296_),
    .Y(_07297_),
    .A1(net10634),
    .A2(_07295_));
 sg13g2_xnor2_1 _25709_ (.Y(_07298_),
    .A(_08668_),
    .B(_07297_));
 sg13g2_buf_2 place9669 (.A(net9668),
    .X(net9669));
 sg13g2_nand3_1 _25711_ (.B(net10581),
    .C(net10446),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[16] ),
    .Y(_07300_));
 sg13g2_o21ai_1 _25712_ (.B1(_07300_),
    .Y(_07301_),
    .A1(net10581),
    .A2(net10306));
 sg13g2_nand2_1 _25713_ (.Y(_07302_),
    .A(net10581),
    .B(net10253));
 sg13g2_a22oi_1 _25714_ (.Y(_07303_),
    .B1(_07302_),
    .B2(_11840_),
    .A2(_07301_),
    .A1(net10452));
 sg13g2_a21o_1 _25715_ (.A2(_07298_),
    .A1(net10188),
    .B1(_07303_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[16] ));
 sg13g2_nor2_1 _25716_ (.A(net10581),
    .B(_07295_),
    .Y(_07304_));
 sg13g2_nand2_1 _25717_ (.Y(_07305_),
    .A(net10581),
    .B(_07295_));
 sg13g2_o21ai_1 _25718_ (.B1(_07305_),
    .Y(_07306_),
    .A1(_11840_),
    .A2(_07304_));
 sg13g2_nand2_1 _25719_ (.Y(_07307_),
    .A(net10580),
    .B(_08784_));
 sg13g2_o21ai_1 _25720_ (.B1(_11840_),
    .Y(_07308_),
    .A1(net10581),
    .A2(_08784_));
 sg13g2_nand2_1 _25721_ (.Y(_07309_),
    .A(_07307_),
    .B(_07308_));
 sg13g2_nand2_1 _25722_ (.Y(_07310_),
    .A(net10634),
    .B(_07309_));
 sg13g2_o21ai_1 _25723_ (.B1(_07310_),
    .Y(_07311_),
    .A1(net10634),
    .A2(_07306_));
 sg13g2_xnor2_1 _25724_ (.Y(_07312_),
    .A(_08655_),
    .B(_07311_));
 sg13g2_nand3_1 _25725_ (.B(net10578),
    .C(net10446),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[17] ),
    .Y(_07313_));
 sg13g2_o21ai_1 _25726_ (.B1(_07313_),
    .Y(_07314_),
    .A1(net10578),
    .A2(net10306));
 sg13g2_nand2_1 _25727_ (.Y(_07315_),
    .A(net10578),
    .B(net10253));
 sg13g2_a22oi_1 _25728_ (.Y(_07316_),
    .B1(_07315_),
    .B2(_11845_),
    .A2(_07314_),
    .A1(net10452));
 sg13g2_a21o_1 _25729_ (.A2(_07312_),
    .A1(net10188),
    .B1(_07316_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[17] ));
 sg13g2_o21ai_1 _25730_ (.B1(_08654_),
    .Y(_07317_),
    .A1(_08652_),
    .A2(_07309_));
 sg13g2_nand2_1 _25731_ (.Y(_07318_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[17] ),
    .B(net10578));
 sg13g2_a21oi_1 _25732_ (.A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[17] ),
    .A2(net10578),
    .Y(_07319_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[16] ));
 sg13g2_a22oi_1 _25733_ (.Y(_07320_),
    .B1(_07319_),
    .B2(_07305_),
    .A2(_07304_),
    .A1(_07318_));
 sg13g2_a21oi_1 _25734_ (.A1(_11845_),
    .A2(_08653_),
    .Y(_07321_),
    .B1(net10634));
 sg13g2_a22oi_1 _25735_ (.Y(_07322_),
    .B1(_07320_),
    .B2(_07321_),
    .A2(_07317_),
    .A1(net10634));
 sg13g2_xnor2_1 _25736_ (.Y(_07323_),
    .A(_08664_),
    .B(_07322_));
 sg13g2_nand3_1 _25737_ (.B(net10576),
    .C(net10446),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[18] ),
    .Y(_07324_));
 sg13g2_o21ai_1 _25738_ (.B1(_07324_),
    .Y(_07325_),
    .A1(net10576),
    .A2(net10306));
 sg13g2_nand2_1 _25739_ (.Y(_07326_),
    .A(net10576),
    .B(net10253));
 sg13g2_a22oi_1 _25740_ (.Y(_07327_),
    .B1(_07326_),
    .B2(_08786_),
    .A2(_07325_),
    .A1(net10452));
 sg13g2_a21o_1 _25741_ (.A2(_07323_),
    .A1(net10188),
    .B1(_07327_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[18] ));
 sg13g2_or2_1 _25742_ (.X(_07328_),
    .B(_08733_),
    .A(_08727_));
 sg13g2_nand4_1 _25743_ (.B(_08664_),
    .C(_08668_),
    .A(_08655_),
    .Y(_07329_),
    .D(_08737_));
 sg13g2_nor2_1 _25744_ (.A(_07328_),
    .B(_07329_),
    .Y(_07330_));
 sg13g2_inv_1 _25745_ (.Y(_07331_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[18] ));
 sg13g2_a221oi_1 _25746_ (.B2(_07281_),
    .C1(_07283_),
    .B1(net10516),
    .A1(net10515),
    .Y(_07332_),
    .A2(net10583));
 sg13g2_nor2_1 _25747_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[16] ),
    .B(net10580),
    .Y(_07333_));
 sg13g2_or2_1 _25748_ (.X(_07334_),
    .B(_07333_),
    .A(_07294_));
 sg13g2_nand2_1 _25749_ (.Y(_07335_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[16] ),
    .B(net10580));
 sg13g2_o21ai_1 _25750_ (.B1(_07335_),
    .Y(_07336_),
    .A1(_07332_),
    .A2(_07334_));
 sg13g2_nand2_1 _25751_ (.Y(_07337_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[17] ),
    .B(_07336_));
 sg13g2_o21ai_1 _25752_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[17] ),
    .Y(_07338_),
    .A1(net10578),
    .A2(_07336_));
 sg13g2_a22oi_1 _25753_ (.Y(_07339_),
    .B1(_07337_),
    .B2(_07338_),
    .A2(_07331_),
    .A1(_08786_));
 sg13g2_a221oi_1 _25754_ (.B2(_07330_),
    .C1(_07339_),
    .B1(_07255_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[18] ),
    .Y(_07340_),
    .A2(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[18] ));
 sg13g2_buf_2 place9663 (.A(_03812_),
    .X(net9663));
 sg13g2_nor3_1 _25756_ (.A(_07248_),
    .B(_07328_),
    .C(_07329_),
    .Y(_07342_));
 sg13g2_o21ai_1 _25757_ (.B1(_07342_),
    .Y(_07343_),
    .A1(_07159_),
    .A2(_07189_));
 sg13g2_buf_2 place9654 (.A(_03822_),
    .X(net9654));
 sg13g2_and2_1 _25759_ (.A(_07340_),
    .B(_07343_),
    .X(_07345_));
 sg13g2_a21oi_1 _25760_ (.A1(_08792_),
    .A2(_07317_),
    .Y(_07346_),
    .B1(_08787_));
 sg13g2_mux2_1 _25761_ (.A0(_07345_),
    .A1(_07346_),
    .S(net10634),
    .X(_07347_));
 sg13g2_xnor2_1 _25762_ (.Y(_07348_),
    .A(_08661_),
    .B(_07347_));
 sg13g2_nand3_1 _25763_ (.B(net10574),
    .C(net10446),
    .A(net10514),
    .Y(_07349_));
 sg13g2_o21ai_1 _25764_ (.B1(_07349_),
    .Y(_07350_),
    .A1(net10574),
    .A2(_07148_));
 sg13g2_a21oi_1 _25765_ (.A1(net10574),
    .A2(_07207_),
    .Y(_07351_),
    .B1(net10514));
 sg13g2_a21oi_1 _25766_ (.A1(net10452),
    .A2(_07350_),
    .Y(_07352_),
    .B1(_07351_));
 sg13g2_a21o_2 _25767_ (.A2(_07348_),
    .A1(_07153_),
    .B1(_07352_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[19] ));
 sg13g2_buf_16 clkbuf_leaf_412_clk (.X(clknet_leaf_412_clk),
    .A(clknet_8_91_0_clk));
 sg13g2_nor2b_1 _25769_ (.A(net10636),
    .B_N(net10599),
    .Y(_07354_));
 sg13g2_nor2_1 _25770_ (.A(net10599),
    .B(net10304),
    .Y(_07355_));
 sg13g2_o21ai_1 _25771_ (.B1(net10520),
    .Y(_07356_),
    .A1(_07354_),
    .A2(_07355_));
 sg13g2_xnor2_1 _25772_ (.Y(_07357_),
    .A(_08832_),
    .B(_07356_));
 sg13g2_nand3_1 _25773_ (.B(net10513),
    .C(net10449),
    .A(net10572),
    .Y(_07358_));
 sg13g2_o21ai_1 _25774_ (.B1(_07358_),
    .Y(_07359_),
    .A1(net10513),
    .A2(net10308));
 sg13g2_nand2_1 _25775_ (.Y(_07360_),
    .A(net10513),
    .B(net10255));
 sg13g2_a22oi_1 _25776_ (.Y(_07361_),
    .B1(_07360_),
    .B2(net10400),
    .A2(_07359_),
    .A1(net10454));
 sg13g2_a21o_1 _25777_ (.A2(_07357_),
    .A1(net10190),
    .B1(_07361_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[1] ));
 sg13g2_a21oi_2 _25778_ (.B1(_08796_),
    .Y(_07362_),
    .A2(_08784_),
    .A1(_08669_));
 sg13g2_and2_1 _25779_ (.A(_02611_),
    .B(_07345_),
    .X(_07363_));
 sg13g2_a21oi_1 _25780_ (.A1(_07340_),
    .A2(_07343_),
    .Y(_07364_),
    .B1(_02611_));
 sg13g2_nor2_1 _25781_ (.A(net10514),
    .B(_07364_),
    .Y(_07365_));
 sg13g2_o21ai_1 _25782_ (.B1(_07193_),
    .Y(_07366_),
    .A1(_07363_),
    .A2(_07365_));
 sg13g2_o21ai_1 _25783_ (.B1(_07366_),
    .Y(_07367_),
    .A1(_07193_),
    .A2(_07362_));
 sg13g2_xor2_1 _25784_ (.B(_07367_),
    .A(_08641_),
    .X(_07368_));
 sg13g2_nor2_1 _25785_ (.A(_11862_),
    .B(_02650_),
    .Y(_07369_));
 sg13g2_nand2_1 _25786_ (.Y(_07370_),
    .A(net10446),
    .B(_07369_));
 sg13g2_o21ai_1 _25787_ (.B1(_07370_),
    .Y(_07371_),
    .A1(net10567),
    .A2(_07148_));
 sg13g2_nand2_1 _25788_ (.Y(_07372_),
    .A(net10567),
    .B(_07207_));
 sg13g2_a22oi_1 _25789_ (.Y(_07373_),
    .B1(_07372_),
    .B2(_11862_),
    .A2(_07371_),
    .A1(net10452));
 sg13g2_a21o_2 _25790_ (.A2(_07368_),
    .A1(_07153_),
    .B1(_07373_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[20] ));
 sg13g2_a21oi_1 _25791_ (.A1(_02650_),
    .A2(_07362_),
    .Y(_07374_),
    .B1(net10512));
 sg13g2_a21oi_1 _25792_ (.A1(net10567),
    .A2(_08797_),
    .Y(_07375_),
    .B1(_07374_));
 sg13g2_a221oi_1 _25793_ (.B2(_07343_),
    .C1(_02611_),
    .B1(_07340_),
    .A1(_11862_),
    .Y(_07376_),
    .A2(_02650_));
 sg13g2_nand2_1 _25794_ (.Y(_07377_),
    .A(net10567),
    .B(net10514));
 sg13g2_nand2_1 _25795_ (.Y(_07378_),
    .A(net10512),
    .B(net10514));
 sg13g2_a22oi_1 _25796_ (.Y(_07379_),
    .B1(_07377_),
    .B2(_07378_),
    .A2(_07343_),
    .A1(_07340_));
 sg13g2_a21oi_1 _25797_ (.A1(_07377_),
    .A2(_07378_),
    .Y(_07380_),
    .B1(_02611_));
 sg13g2_nor4_1 _25798_ (.A(_07369_),
    .B(_07376_),
    .C(_07379_),
    .D(_07380_),
    .Y(_07381_));
 sg13g2_nand2_1 _25799_ (.Y(_07382_),
    .A(_07193_),
    .B(_07381_));
 sg13g2_o21ai_1 _25800_ (.B1(_07382_),
    .Y(_07383_),
    .A1(_07193_),
    .A2(_07375_));
 sg13g2_xor2_1 _25801_ (.B(_07383_),
    .A(_08631_),
    .X(_07384_));
 sg13g2_nand3_1 _25802_ (.B(net10565),
    .C(net10446),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[21] ),
    .Y(_07385_));
 sg13g2_o21ai_1 _25803_ (.B1(_07385_),
    .Y(_07386_),
    .A1(net10565),
    .A2(_07148_));
 sg13g2_nand2_1 _25804_ (.Y(_07387_),
    .A(net10565),
    .B(_07207_));
 sg13g2_a22oi_1 _25805_ (.Y(_07388_),
    .B1(_07387_),
    .B2(_08801_),
    .A2(_07386_),
    .A1(_08292_));
 sg13g2_a21o_2 _25806_ (.A2(_07384_),
    .A1(_07153_),
    .B1(_07388_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[21] ));
 sg13g2_nand2_1 _25807_ (.Y(_07389_),
    .A(_08801_),
    .B(net10565));
 sg13g2_nor2_1 _25808_ (.A(_08801_),
    .B(net10565),
    .Y(_07390_));
 sg13g2_a21oi_1 _25809_ (.A1(_07389_),
    .A2(_07375_),
    .Y(_07391_),
    .B1(_07390_));
 sg13g2_nor2_1 _25810_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[21] ),
    .B(net10565),
    .Y(_07392_));
 sg13g2_nand2_1 _25811_ (.Y(_07393_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[21] ),
    .B(net10564));
 sg13g2_o21ai_1 _25812_ (.B1(_07393_),
    .Y(_07394_),
    .A1(_07381_),
    .A2(_07392_));
 sg13g2_buf_2 place9655 (.A(net9654),
    .X(net9655));
 sg13g2_nand2_1 _25814_ (.Y(_07396_),
    .A(_07193_),
    .B(_07394_));
 sg13g2_o21ai_1 _25815_ (.B1(_07396_),
    .Y(_07397_),
    .A1(_07193_),
    .A2(_07391_));
 sg13g2_xnor2_1 _25816_ (.Y(_07398_),
    .A(_08638_),
    .B(_07397_));
 sg13g2_and2_1 _25817_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[22] ),
    .B(net10561),
    .X(_07399_));
 sg13g2_buf_2 place9653 (.A(_08228_),
    .X(net9653));
 sg13g2_nand2_1 _25819_ (.Y(_07401_),
    .A(_08297_),
    .B(_07399_));
 sg13g2_o21ai_1 _25820_ (.B1(_07401_),
    .Y(_07402_),
    .A1(net10561),
    .A2(_07148_));
 sg13g2_a21oi_1 _25821_ (.A1(net10561),
    .A2(_07207_),
    .Y(_07403_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[22] ));
 sg13g2_a21oi_1 _25822_ (.A1(_08292_),
    .A2(_07402_),
    .Y(_07404_),
    .B1(_07403_));
 sg13g2_a21o_2 _25823_ (.A2(_07398_),
    .A1(_07153_),
    .B1(_07404_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[22] ));
 sg13g2_or2_1 _25824_ (.X(_07405_),
    .B(net10561),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[22] ));
 sg13g2_a21oi_2 _25825_ (.B1(_07399_),
    .Y(_07406_),
    .A2(_07405_),
    .A1(_07394_));
 sg13g2_nor2_1 _25826_ (.A(net10638),
    .B(_07406_),
    .Y(_07407_));
 sg13g2_nand2_1 _25827_ (.Y(_07408_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[18] ),
    .B(_08652_));
 sg13g2_o21ai_1 _25828_ (.B1(_08786_),
    .Y(_07409_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[18] ),
    .A2(_08652_));
 sg13g2_a221oi_1 _25829_ (.B2(_07409_),
    .C1(_08659_),
    .B1(_07408_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[20] ),
    .Y(_07410_),
    .A2(_02650_));
 sg13g2_a21oi_1 _25830_ (.A1(net10512),
    .A2(_02650_),
    .Y(_07411_),
    .B1(_08660_));
 sg13g2_or2_1 _25831_ (.X(_07412_),
    .B(_08634_),
    .A(net10564));
 sg13g2_nor4_1 _25832_ (.A(_08799_),
    .B(_07410_),
    .C(_07411_),
    .D(_07412_),
    .Y(_07413_));
 sg13g2_nand2b_1 _25833_ (.Y(_07414_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[21] ),
    .A_N(_08634_));
 sg13g2_nor4_1 _25834_ (.A(_08799_),
    .B(_07410_),
    .C(_07411_),
    .D(_07414_),
    .Y(_07415_));
 sg13g2_nor3_1 _25835_ (.A(_08801_),
    .B(net10564),
    .C(_08634_),
    .Y(_07416_));
 sg13g2_or4_1 _25836_ (.A(_08636_),
    .B(_07413_),
    .C(_07415_),
    .D(_07416_),
    .X(_07417_));
 sg13g2_buf_2 place9657 (.A(net9656),
    .X(net9657));
 sg13g2_nand3b_1 _25838_ (.B(_08773_),
    .C(_07417_),
    .Y(_07419_),
    .A_N(net10579));
 sg13g2_nand3_1 _25839_ (.B(_08773_),
    .C(_07417_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[16] ),
    .Y(_07420_));
 sg13g2_nand2_1 _25840_ (.Y(_07421_),
    .A(_08751_),
    .B(_08783_));
 sg13g2_a21o_2 _25841_ (.A2(_07420_),
    .A1(_07419_),
    .B1(_07421_),
    .X(_07422_));
 sg13g2_buf_2 place9656 (.A(_03822_),
    .X(net9656));
 sg13g2_nor2_1 _25843_ (.A(_11840_),
    .B(net10580),
    .Y(_07424_));
 sg13g2_or4_1 _25844_ (.A(_08642_),
    .B(_08655_),
    .C(_08661_),
    .D(_08664_),
    .X(_07425_));
 sg13g2_o21ai_1 _25845_ (.B1(_07417_),
    .Y(_07426_),
    .A1(_07424_),
    .A2(_07425_));
 sg13g2_and2_1 _25846_ (.A(_07422_),
    .B(_07426_),
    .X(_07427_));
 sg13g2_buf_16 clkbuf_leaf_416_clk (.X(clknet_leaf_416_clk),
    .A(clknet_8_90_0_clk));
 sg13g2_nor2_1 _25848_ (.A(net10303),
    .B(_07427_),
    .Y(_07429_));
 sg13g2_nor2_1 _25849_ (.A(_07407_),
    .B(_07429_),
    .Y(_07430_));
 sg13g2_xor2_1 _25850_ (.B(_07430_),
    .A(_08627_),
    .X(_07431_));
 sg13g2_nand3_1 _25851_ (.B(net10559),
    .C(_08297_),
    .A(net10511),
    .Y(_07432_));
 sg13g2_o21ai_1 _25852_ (.B1(_07432_),
    .Y(_07433_),
    .A1(net10559),
    .A2(_07148_));
 sg13g2_nand2_1 _25853_ (.Y(_07434_),
    .A(net10559),
    .B(_07207_));
 sg13g2_a22oi_1 _25854_ (.Y(_07435_),
    .B1(_07434_),
    .B2(_11875_),
    .A2(_07433_),
    .A1(_08292_));
 sg13g2_a21o_2 _25855_ (.A2(_07431_),
    .A1(net10187),
    .B1(_07435_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[23] ));
 sg13g2_a21oi_1 _25856_ (.A1(net10559),
    .A2(_07427_),
    .Y(_07436_),
    .B1(_11875_));
 sg13g2_nor2_1 _25857_ (.A(net10559),
    .B(_07427_),
    .Y(_07437_));
 sg13g2_nor2_1 _25858_ (.A(_07436_),
    .B(_07437_),
    .Y(_07438_));
 sg13g2_nor2_1 _25859_ (.A(_08627_),
    .B(_08638_),
    .Y(_07439_));
 sg13g2_nor4_2 _25860_ (.A(_08631_),
    .B(_08641_),
    .C(_07363_),
    .Y(_07440_),
    .D(_07365_));
 sg13g2_a21oi_1 _25861_ (.A1(net10512),
    .A2(net10567),
    .Y(_07441_),
    .B1(net10564));
 sg13g2_nand3_1 _25862_ (.B(net10512),
    .C(net10567),
    .A(net10564),
    .Y(_07442_));
 sg13g2_o21ai_1 _25863_ (.B1(_07442_),
    .Y(_07443_),
    .A1(_08801_),
    .A2(_07441_));
 sg13g2_nor2_1 _25864_ (.A(net10558),
    .B(_07399_),
    .Y(_07444_));
 sg13g2_a21oi_1 _25865_ (.A1(net10558),
    .A2(_07399_),
    .Y(_07445_),
    .B1(net10511));
 sg13g2_nor2_1 _25866_ (.A(_07444_),
    .B(_07445_),
    .Y(_07446_));
 sg13g2_a21o_1 _25867_ (.A2(_07443_),
    .A1(_07439_),
    .B1(_07446_),
    .X(_07447_));
 sg13g2_buf_16 clkbuf_leaf_414_clk (.X(clknet_leaf_414_clk),
    .A(clknet_8_91_0_clk));
 sg13g2_nand2b_1 _25869_ (.Y(_07449_),
    .B(net10303),
    .A_N(_07447_));
 sg13g2_a21oi_2 _25870_ (.B1(_07449_),
    .Y(_07450_),
    .A2(_07440_),
    .A1(_07439_));
 sg13g2_a21oi_1 _25871_ (.A1(net10633),
    .A2(_07438_),
    .Y(_07451_),
    .B1(_07450_));
 sg13g2_xor2_1 _25872_ (.B(_07451_),
    .A(_08622_),
    .X(_07452_));
 sg13g2_nand3_1 _25873_ (.B(net10556),
    .C(net10450),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[24] ),
    .Y(_07453_));
 sg13g2_o21ai_1 _25874_ (.B1(_07453_),
    .Y(_07454_),
    .A1(net10556),
    .A2(net10305));
 sg13g2_nand2_1 _25875_ (.Y(_07455_),
    .A(net10556),
    .B(net10252));
 sg13g2_a22oi_1 _25876_ (.Y(_07456_),
    .B1(_07455_),
    .B2(_08620_),
    .A2(_07454_),
    .A1(net10451));
 sg13g2_a21o_2 _25877_ (.A2(_07452_),
    .A1(_07153_),
    .B1(_07456_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[24] ));
 sg13g2_inv_1 _25878_ (.Y(_07457_),
    .A(_07450_));
 sg13g2_o21ai_1 _25879_ (.B1(net10633),
    .Y(_07458_),
    .A1(_07436_),
    .A2(_07437_));
 sg13g2_a21oi_1 _25880_ (.A1(_08620_),
    .A2(_07458_),
    .Y(_07459_),
    .B1(net10556));
 sg13g2_nor2_1 _25881_ (.A(_08620_),
    .B(_07438_),
    .Y(_07460_));
 sg13g2_nand2_1 _25882_ (.Y(_07461_),
    .A(net10303),
    .B(net10556));
 sg13g2_a21oi_1 _25883_ (.A1(_08620_),
    .A2(_07450_),
    .Y(_07462_),
    .B1(_07461_));
 sg13g2_a221oi_1 _25884_ (.B2(net10556),
    .C1(_07462_),
    .B1(_07460_),
    .A1(_07457_),
    .Y(_07463_),
    .A2(_07459_));
 sg13g2_xnor2_1 _25885_ (.Y(_07464_),
    .A(_08615_),
    .B(_07463_));
 sg13g2_nand3_1 _25886_ (.B(net10553),
    .C(net10450),
    .A(net10510),
    .Y(_07465_));
 sg13g2_o21ai_1 _25887_ (.B1(_07465_),
    .Y(_07466_),
    .A1(net10553),
    .A2(net10305));
 sg13g2_a21oi_1 _25888_ (.A1(net10553),
    .A2(net10252),
    .Y(_07467_),
    .B1(net10510));
 sg13g2_a21oi_1 _25889_ (.A1(net10451),
    .A2(_07466_),
    .Y(_07468_),
    .B1(_07467_));
 sg13g2_a21o_2 _25890_ (.A2(_07464_),
    .A1(net10187),
    .B1(_07468_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[25] ));
 sg13g2_nor2b_2 _25891_ (.A(_08606_),
    .B_N(_08607_),
    .Y(_07469_));
 sg13g2_or2_1 _25892_ (.X(_07470_),
    .B(net10558),
    .A(net10555));
 sg13g2_nand2b_1 _25893_ (.Y(_07471_),
    .B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[24] ),
    .A_N(net10558));
 sg13g2_a22oi_1 _25894_ (.Y(_07472_),
    .B1(_07470_),
    .B2(_07471_),
    .A2(_07426_),
    .A1(_07422_));
 sg13g2_nand2b_1 _25895_ (.Y(_07473_),
    .B(net10511),
    .A_N(net10555));
 sg13g2_nand2_1 _25896_ (.Y(_07474_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[24] ),
    .B(net10511));
 sg13g2_a22oi_1 _25897_ (.Y(_07475_),
    .B1(_07473_),
    .B2(_07474_),
    .A2(_07426_),
    .A1(_07422_));
 sg13g2_a21oi_1 _25898_ (.A1(_07473_),
    .A2(_07474_),
    .Y(_07476_),
    .B1(net10558));
 sg13g2_nor4_2 _25899_ (.A(_08621_),
    .B(_07472_),
    .C(_07475_),
    .Y(_07477_),
    .D(_07476_));
 sg13g2_a21oi_1 _25900_ (.A1(_08614_),
    .A2(_07477_),
    .Y(_07478_),
    .B1(_08611_));
 sg13g2_nand2_1 _25901_ (.Y(_07479_),
    .A(_08615_),
    .B(_08622_));
 sg13g2_or2_1 _25902_ (.X(_07480_),
    .B(_07479_),
    .A(_08627_));
 sg13g2_or2_1 _25903_ (.X(_07481_),
    .B(_08636_),
    .A(_08634_));
 sg13g2_nand2_2 _25904_ (.Y(_07482_),
    .A(_07481_),
    .B(_07394_));
 sg13g2_nor2_1 _25905_ (.A(net10510),
    .B(net10553),
    .Y(_07483_));
 sg13g2_nand2_1 _25906_ (.Y(_07484_),
    .A(net10510),
    .B(net10553));
 sg13g2_nand2_1 _25907_ (.Y(_07485_),
    .A(net10555),
    .B(_07446_));
 sg13g2_o21ai_1 _25908_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[24] ),
    .Y(_07486_),
    .A1(net10555),
    .A2(_07446_));
 sg13g2_nand3_1 _25909_ (.B(_07485_),
    .C(_07486_),
    .A(_07484_),
    .Y(_07487_));
 sg13g2_nand2b_2 _25910_ (.Y(_07488_),
    .B(_07487_),
    .A_N(_07483_));
 sg13g2_o21ai_1 _25911_ (.B1(_07488_),
    .Y(_07489_),
    .A1(_07480_),
    .A2(_07482_));
 sg13g2_mux2_1 _25912_ (.A0(_07478_),
    .A1(_07489_),
    .S(net10303),
    .X(_07490_));
 sg13g2_xnor2_1 _25913_ (.Y(_07491_),
    .A(_07469_),
    .B(_07490_));
 sg13g2_nand3_1 _25914_ (.B(net10550),
    .C(net10450),
    .A(net10509),
    .Y(_07492_));
 sg13g2_o21ai_1 _25915_ (.B1(_07492_),
    .Y(_07493_),
    .A1(net10550),
    .A2(net10305));
 sg13g2_buf_2 place9652 (.A(net9650),
    .X(net9652));
 sg13g2_a21oi_1 _25917_ (.A1(net10550),
    .A2(net10252),
    .Y(_07495_),
    .B1(net10509));
 sg13g2_a21oi_1 _25918_ (.A1(net10451),
    .A2(_07493_),
    .Y(_07496_),
    .B1(_07495_));
 sg13g2_a21o_2 _25919_ (.A2(_07491_),
    .A1(net10187),
    .B1(_07496_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[26] ));
 sg13g2_nor2_2 _25920_ (.A(_07469_),
    .B(_07480_),
    .Y(_07497_));
 sg13g2_nand2_1 _25921_ (.Y(_07498_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[26] ),
    .B(net10549));
 sg13g2_a21oi_1 _25922_ (.A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[23] ),
    .A2(net10557),
    .Y(_07499_),
    .B1(net10554));
 sg13g2_nand3_1 _25923_ (.B(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[23] ),
    .C(net10557),
    .A(net10554),
    .Y(_07500_));
 sg13g2_o21ai_1 _25924_ (.B1(_07500_),
    .Y(_07501_),
    .A1(_08620_),
    .A2(_07499_));
 sg13g2_nand2_1 _25925_ (.Y(_07502_),
    .A(net10552),
    .B(_07501_));
 sg13g2_o21ai_1 _25926_ (.B1(net10510),
    .Y(_07503_),
    .A1(net10552),
    .A2(_07501_));
 sg13g2_nand3_1 _25927_ (.B(_07502_),
    .C(_07503_),
    .A(_07498_),
    .Y(_07504_));
 sg13g2_o21ai_1 _25928_ (.B1(_07504_),
    .Y(_07505_),
    .A1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[26] ),
    .A2(net10549));
 sg13g2_nand2b_1 _25929_ (.Y(_07506_),
    .B(_07427_),
    .A_N(_08628_));
 sg13g2_nor2b_1 _25930_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[23] ),
    .B_N(net10557),
    .Y(_07507_));
 sg13g2_nor2_1 _25931_ (.A(net10554),
    .B(_07507_),
    .Y(_07508_));
 sg13g2_a21oi_1 _25932_ (.A1(net10554),
    .A2(_07507_),
    .Y(_07509_),
    .B1(_08620_));
 sg13g2_nor2_1 _25933_ (.A(_07508_),
    .B(_07509_),
    .Y(_07510_));
 sg13g2_a21o_1 _25934_ (.A2(_07510_),
    .A1(_08614_),
    .B1(_08611_),
    .X(_07511_));
 sg13g2_nand2_1 _25935_ (.Y(_07512_),
    .A(net10549),
    .B(_07511_));
 sg13g2_nand2_1 _25936_ (.Y(_07513_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[26] ),
    .B(_07512_));
 sg13g2_o21ai_1 _25937_ (.B1(_07513_),
    .Y(_07514_),
    .A1(net10549),
    .A2(_07511_));
 sg13g2_a21oi_1 _25938_ (.A1(_07506_),
    .A2(_07514_),
    .Y(_07515_),
    .B1(net10303));
 sg13g2_a21oi_1 _25939_ (.A1(net10303),
    .A2(_07505_),
    .Y(_07516_),
    .B1(_07515_));
 sg13g2_a21oi_1 _25940_ (.A1(_07407_),
    .A2(_07497_),
    .Y(_07517_),
    .B1(_07516_));
 sg13g2_xnor2_1 _25941_ (.Y(_07518_),
    .A(_08647_),
    .B(_07517_));
 sg13g2_nand3_1 _25942_ (.B(net10547),
    .C(net10450),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[27] ),
    .Y(_07519_));
 sg13g2_o21ai_1 _25943_ (.B1(_07519_),
    .Y(_07520_),
    .A1(net10547),
    .A2(net10305));
 sg13g2_a21oi_1 _25944_ (.A1(net10547),
    .A2(net10252),
    .Y(_07521_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[27] ));
 sg13g2_a21oi_1 _25945_ (.A1(net10451),
    .A2(_07520_),
    .Y(_07522_),
    .B1(_07521_));
 sg13g2_a21o_2 _25946_ (.A2(_07518_),
    .A1(net10187),
    .B1(_07522_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[27] ));
 sg13g2_nand4_1 _25947_ (.B(_08647_),
    .C(_07440_),
    .A(_07481_),
    .Y(_07523_),
    .D(_07497_));
 sg13g2_a21o_1 _25948_ (.A2(_07447_),
    .A1(net10555),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[24] ),
    .X(_07524_));
 sg13g2_o21ai_1 _25949_ (.B1(_07524_),
    .Y(_07525_),
    .A1(net10555),
    .A2(_07447_));
 sg13g2_o21ai_1 _25950_ (.B1(_07484_),
    .Y(_07526_),
    .A1(_07483_),
    .A2(_07525_));
 sg13g2_nand2_1 _25951_ (.Y(_07527_),
    .A(net10550),
    .B(_07526_));
 sg13g2_o21ai_1 _25952_ (.B1(net10509),
    .Y(_07528_),
    .A1(net10549),
    .A2(_07526_));
 sg13g2_nor2_1 _25953_ (.A(net10508),
    .B(net10547),
    .Y(_07529_));
 sg13g2_a21oi_1 _25954_ (.A1(_07527_),
    .A2(_07528_),
    .Y(_07530_),
    .B1(_07529_));
 sg13g2_a21oi_1 _25955_ (.A1(net10508),
    .A2(net10547),
    .Y(_07531_),
    .B1(_07530_));
 sg13g2_a21oi_1 _25956_ (.A1(_07523_),
    .A2(_07531_),
    .Y(_07532_),
    .B1(net10633));
 sg13g2_a21oi_1 _25957_ (.A1(net10633),
    .A2(_08815_),
    .Y(_07533_),
    .B1(_07532_));
 sg13g2_xnor2_1 _25958_ (.Y(_07534_),
    .A(_08597_),
    .B(_07533_));
 sg13g2_nand3_1 _25959_ (.B(net10545),
    .C(net10450),
    .A(net10507),
    .Y(_07535_));
 sg13g2_o21ai_1 _25960_ (.B1(_07535_),
    .Y(_07536_),
    .A1(net10545),
    .A2(net10305));
 sg13g2_a21oi_1 _25961_ (.A1(net10545),
    .A2(net10252),
    .Y(_07537_),
    .B1(net10507));
 sg13g2_a21oi_1 _25962_ (.A1(net10451),
    .A2(_07536_),
    .Y(_07538_),
    .B1(_07537_));
 sg13g2_a21o_1 _25963_ (.A2(_07534_),
    .A1(net10187),
    .B1(_07538_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[28] ));
 sg13g2_buf_2 place9651 (.A(net9650),
    .X(net9651));
 sg13g2_nand3_1 _25965_ (.B(_08647_),
    .C(_07497_),
    .A(_08597_),
    .Y(_07540_));
 sg13g2_buf_2 place9650 (.A(_10023_),
    .X(net9650));
 sg13g2_nor2_1 _25967_ (.A(net10507),
    .B(net10544),
    .Y(_07542_));
 sg13g2_nand2_1 _25968_ (.Y(_07543_),
    .A(_08798_),
    .B(_07505_));
 sg13g2_nor2_1 _25969_ (.A(_08798_),
    .B(_07505_),
    .Y(_07544_));
 sg13g2_a221oi_1 _25970_ (.B2(_07543_),
    .C1(_07544_),
    .B1(net10508),
    .A1(net10507),
    .Y(_07545_),
    .A2(net10544));
 sg13g2_nor2_2 _25971_ (.A(_07542_),
    .B(_07545_),
    .Y(_07546_));
 sg13g2_inv_1 _25972_ (.Y(_07547_),
    .A(_07546_));
 sg13g2_o21ai_1 _25973_ (.B1(_07547_),
    .Y(_07548_),
    .A1(_07406_),
    .A2(_07540_));
 sg13g2_nor3_2 _25974_ (.A(_08597_),
    .B(_08608_),
    .C(_08647_),
    .Y(_07549_));
 sg13g2_nor2b_1 _25975_ (.A(_08615_),
    .B_N(_07549_),
    .Y(_07550_));
 sg13g2_nand2_1 _25976_ (.Y(_07551_),
    .A(net10550),
    .B(_08611_));
 sg13g2_nand2_1 _25977_ (.Y(_07552_),
    .A(net10509),
    .B(_07551_));
 sg13g2_o21ai_1 _25978_ (.B1(_07552_),
    .Y(_07553_),
    .A1(net10550),
    .A2(_08611_));
 sg13g2_a21oi_1 _25979_ (.A1(_08646_),
    .A2(_07553_),
    .Y(_07554_),
    .B1(_08645_));
 sg13g2_nand2_1 _25980_ (.Y(_07555_),
    .A(net10545),
    .B(_07554_));
 sg13g2_nand2_1 _25981_ (.Y(_07556_),
    .A(net10507),
    .B(_07555_));
 sg13g2_or2_1 _25982_ (.X(_07557_),
    .B(_07554_),
    .A(net10545));
 sg13g2_a221oi_1 _25983_ (.B2(_07557_),
    .C1(net10303),
    .B1(_07556_),
    .A1(_07477_),
    .Y(_07558_),
    .A2(_07550_));
 sg13g2_a21oi_1 _25984_ (.A1(net10303),
    .A2(_07548_),
    .Y(_07559_),
    .B1(_07558_));
 sg13g2_xnor2_1 _25985_ (.Y(_07560_),
    .A(_08600_),
    .B(_07559_));
 sg13g2_nand3_1 _25986_ (.B(net10543),
    .C(net10450),
    .A(net10506),
    .Y(_07561_));
 sg13g2_o21ai_1 _25987_ (.B1(_07561_),
    .Y(_07562_),
    .A1(net10543),
    .A2(net10305));
 sg13g2_a21oi_1 _25988_ (.A1(net10543),
    .A2(net10252),
    .Y(_07563_),
    .B1(net10506));
 sg13g2_a21oi_1 _25989_ (.A1(net10451),
    .A2(_07562_),
    .Y(_07564_),
    .B1(_07563_));
 sg13g2_a21o_1 _25990_ (.A2(_07560_),
    .A1(net10187),
    .B1(_07564_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[29] ));
 sg13g2_a21oi_1 _25991_ (.A1(net10599),
    .A2(net10513),
    .Y(_07565_),
    .B1(_07355_));
 sg13g2_nor2_1 _25992_ (.A(net10599),
    .B(_08682_),
    .Y(_07566_));
 sg13g2_nor3_1 _25993_ (.A(net10400),
    .B(_07566_),
    .C(_07354_),
    .Y(_07567_));
 sg13g2_a21oi_1 _25994_ (.A1(net10400),
    .A2(_07565_),
    .Y(_07568_),
    .B1(_07567_));
 sg13g2_xor2_1 _25995_ (.B(net10636),
    .A(net10572),
    .X(_07569_));
 sg13g2_a22oi_1 _25996_ (.Y(_07570_),
    .B1(_07569_),
    .B2(net10513),
    .A2(_07568_),
    .A1(net10520));
 sg13g2_xor2_1 _25997_ (.B(_07570_),
    .A(_08842_),
    .X(_07571_));
 sg13g2_nand3_1 _25998_ (.B(net10540),
    .C(net10449),
    .A(net10505),
    .Y(_07572_));
 sg13g2_o21ai_1 _25999_ (.B1(_07572_),
    .Y(_07573_),
    .A1(net10540),
    .A2(net10308));
 sg13g2_a21oi_1 _26000_ (.A1(net10540),
    .A2(net10255),
    .Y(_07574_),
    .B1(net10505));
 sg13g2_a21oi_1 _26001_ (.A1(net10454),
    .A2(_07573_),
    .Y(_07575_),
    .B1(_07574_));
 sg13g2_a21o_1 _26002_ (.A2(_07571_),
    .A1(net10190),
    .B1(_07575_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[2] ));
 sg13g2_inv_1 _26003_ (.Y(_07576_),
    .A(_07482_));
 sg13g2_nor2_1 _26004_ (.A(net10506),
    .B(net10543),
    .Y(_07577_));
 sg13g2_nor3_1 _26005_ (.A(net10638),
    .B(_07540_),
    .C(_07577_),
    .Y(_07578_));
 sg13g2_nand2b_2 _26006_ (.Y(_07579_),
    .B(net10506),
    .A_N(net10542));
 sg13g2_buf_2 place9649 (.A(_10023_),
    .X(net9649));
 sg13g2_nand3b_1 _26008_ (.B(_07549_),
    .C(_07579_),
    .Y(_07581_),
    .A_N(_07478_));
 sg13g2_nor2b_1 _26009_ (.A(net10506),
    .B_N(net10542),
    .Y(_07582_));
 sg13g2_nand2_1 _26010_ (.Y(_07583_),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[27] ),
    .B(_08606_));
 sg13g2_nor2_1 _26011_ (.A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[27] ),
    .B(_08606_),
    .Y(_07584_));
 sg13g2_a21oi_1 _26012_ (.A1(net10508),
    .A2(_07583_),
    .Y(_07585_),
    .B1(_07584_));
 sg13g2_nor2_1 _26013_ (.A(_08817_),
    .B(_07585_),
    .Y(_07586_));
 sg13g2_a21oi_1 _26014_ (.A1(net10507),
    .A2(_02952_),
    .Y(_07587_),
    .B1(_07586_));
 sg13g2_o21ai_1 _26015_ (.B1(_07579_),
    .Y(_07588_),
    .A1(_07582_),
    .A2(_07587_));
 sg13g2_and2_1 _26016_ (.A(net10638),
    .B(_07588_),
    .X(_07589_));
 sg13g2_nand2_1 _26017_ (.Y(_07590_),
    .A(_08605_),
    .B(_07488_));
 sg13g2_nor2_1 _26018_ (.A(_08605_),
    .B(_07488_),
    .Y(_07591_));
 sg13g2_a221oi_1 _26019_ (.B2(_07590_),
    .C1(_07591_),
    .B1(net10509),
    .A1(net10508),
    .Y(_07592_),
    .A2(net10547));
 sg13g2_nor3_1 _26020_ (.A(_07529_),
    .B(_07542_),
    .C(_07592_),
    .Y(_07593_));
 sg13g2_a221oi_1 _26021_ (.B2(net10545),
    .C1(_07593_),
    .B1(net10507),
    .A1(net10506),
    .Y(_07594_),
    .A2(net10542));
 sg13g2_nor3_1 _26022_ (.A(net10638),
    .B(_07577_),
    .C(_07594_),
    .Y(_07595_));
 sg13g2_a221oi_1 _26023_ (.B2(_07589_),
    .C1(_07595_),
    .B1(_07581_),
    .A1(_07576_),
    .Y(_07596_),
    .A2(_07578_));
 sg13g2_xnor2_1 _26024_ (.Y(_07597_),
    .A(_08591_),
    .B(_07596_));
 sg13g2_nand3_1 _26025_ (.B(net10537),
    .C(net10450),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[30] ),
    .Y(_07598_));
 sg13g2_o21ai_1 _26026_ (.B1(_07598_),
    .Y(_07599_),
    .A1(net10537),
    .A2(net10305));
 sg13g2_a21oi_1 _26027_ (.A1(net10537),
    .A2(net10252),
    .Y(_07600_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[30] ));
 sg13g2_a21oi_1 _26028_ (.A1(net10451),
    .A2(_07599_),
    .Y(_07601_),
    .B1(_07600_));
 sg13g2_a21o_1 _26029_ (.A2(_07597_),
    .A1(net10187),
    .B1(_07601_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[30] ));
 sg13g2_nand2_1 _26030_ (.Y(_07602_),
    .A(_08591_),
    .B(_08600_));
 sg13g2_or4_1 _26031_ (.A(net10638),
    .B(_07406_),
    .C(_07540_),
    .D(_07602_),
    .X(_07603_));
 sg13g2_and3_1 _26032_ (.X(_07604_),
    .A(net10552),
    .B(_07579_),
    .C(_07549_));
 sg13g2_nand3b_1 _26033_ (.B(_07579_),
    .C(_07549_),
    .Y(_07605_),
    .A_N(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[25] ));
 sg13g2_inv_1 _26034_ (.Y(_07606_),
    .A(_07605_));
 sg13g2_o21ai_1 _26035_ (.B1(_07477_),
    .Y(_07607_),
    .A1(_07604_),
    .A2(_07606_));
 sg13g2_nand3_1 _26036_ (.B(_08611_),
    .C(_07549_),
    .A(_07579_),
    .Y(_07608_));
 sg13g2_and2_1 _26037_ (.A(_07588_),
    .B(_07608_),
    .X(_07609_));
 sg13g2_nand4_1 _26038_ (.B(_08590_),
    .C(_07607_),
    .A(net10638),
    .Y(_07610_),
    .D(_07609_));
 sg13g2_nor2b_1 _26039_ (.A(net10638),
    .B_N(net10537),
    .Y(_07611_));
 sg13g2_a21oi_1 _26040_ (.A1(net10543),
    .A2(_07546_),
    .Y(_07612_),
    .B1(net10506));
 sg13g2_nor2_1 _26041_ (.A(net10543),
    .B(_07546_),
    .Y(_07613_));
 sg13g2_o21ai_1 _26042_ (.B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[30] ),
    .Y(_07614_),
    .A1(net10638),
    .A2(net10537));
 sg13g2_o21ai_1 _26043_ (.B1(_07614_),
    .Y(_07615_),
    .A1(_07612_),
    .A2(_07613_));
 sg13g2_o21ai_1 _26044_ (.B1(_07615_),
    .Y(_07616_),
    .A1(_08589_),
    .A2(_07611_));
 sg13g2_nand3_1 _26045_ (.B(_07610_),
    .C(_07616_),
    .A(_07603_),
    .Y(_07617_));
 sg13g2_xor2_1 _26046_ (.B(_07617_),
    .A(_08593_),
    .X(_07618_));
 sg13g2_nand3_1 _26047_ (.B(net10534),
    .C(net10450),
    .A(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[31] ),
    .Y(_07619_));
 sg13g2_o21ai_1 _26048_ (.B1(_07619_),
    .Y(_07620_),
    .A1(net10534),
    .A2(net10305));
 sg13g2_a21oi_1 _26049_ (.A1(net10534),
    .A2(net10252),
    .Y(_07621_),
    .B1(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[31] ));
 sg13g2_a21oi_1 _26050_ (.A1(net10451),
    .A2(_07620_),
    .Y(_07622_),
    .B1(_07621_));
 sg13g2_a21o_1 _26051_ (.A2(_07618_),
    .A1(net10187),
    .B1(_07622_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[31] ));
 sg13g2_a21oi_1 _26052_ (.A1(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[0] ),
    .A2(_07566_),
    .Y(_07623_),
    .B1(_08684_));
 sg13g2_o21ai_1 _26053_ (.B1(_08677_),
    .Y(_07624_),
    .A1(_07623_),
    .A2(_08688_));
 sg13g2_nor2_1 _26054_ (.A(net10505),
    .B(net10540),
    .Y(_07625_));
 sg13g2_a221oi_1 _26055_ (.B2(net10572),
    .C1(_07168_),
    .B1(_07165_),
    .A1(net10505),
    .Y(_07626_),
    .A2(net10540));
 sg13g2_nor3_1 _26056_ (.A(net10637),
    .B(_07625_),
    .C(_07626_),
    .Y(_07627_));
 sg13g2_a21oi_1 _26057_ (.A1(net10637),
    .A2(_07624_),
    .Y(_07628_),
    .B1(_07627_));
 sg13g2_xor2_1 _26058_ (.B(_07628_),
    .A(_08840_),
    .X(_07629_));
 sg13g2_nand3_1 _26059_ (.B(net10532),
    .C(net10449),
    .A(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[3] ),
    .Y(_07630_));
 sg13g2_o21ai_1 _26060_ (.B1(_07630_),
    .Y(_07631_),
    .A1(net10532),
    .A2(net10308));
 sg13g2_nand2_1 _26061_ (.Y(_07632_),
    .A(net10532),
    .B(net10255));
 sg13g2_a22oi_1 _26062_ (.Y(_07633_),
    .B1(_07632_),
    .B2(_08680_),
    .A2(_07631_),
    .A1(net10454));
 sg13g2_a21o_1 _26063_ (.A2(_07629_),
    .A1(net10190),
    .B1(_07633_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[3] ));
 sg13g2_nand2_2 _26064_ (.Y(_07634_),
    .A(_08685_),
    .B(_08690_));
 sg13g2_nor2_1 _26065_ (.A(_07163_),
    .B(_07169_),
    .Y(_07635_));
 sg13g2_nor2_1 _26066_ (.A(net10637),
    .B(_07635_),
    .Y(_07636_));
 sg13g2_a21oi_1 _26067_ (.A1(net10637),
    .A2(_07634_),
    .Y(_07637_),
    .B1(_07636_));
 sg13g2_xnor2_1 _26068_ (.Y(_07638_),
    .A(_08839_),
    .B(_07637_));
 sg13g2_nand3_1 _26069_ (.B(net10530),
    .C(net10449),
    .A(net10504),
    .Y(_07639_));
 sg13g2_o21ai_1 _26070_ (.B1(_07639_),
    .Y(_07640_),
    .A1(net10530),
    .A2(net10308));
 sg13g2_a21oi_1 _26071_ (.A1(net10530),
    .A2(net10255),
    .Y(_07641_),
    .B1(net10504));
 sg13g2_a21oi_1 _26072_ (.A1(net10454),
    .A2(_07640_),
    .Y(_07642_),
    .B1(_07641_));
 sg13g2_a21o_1 _26073_ (.A2(_07638_),
    .A1(net10190),
    .B1(_07642_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[4] ));
 sg13g2_inv_1 _26074_ (.Y(_07643_),
    .A(_07634_));
 sg13g2_a21oi_1 _26075_ (.A1(_08701_),
    .A2(_07643_),
    .Y(_07644_),
    .B1(net10504));
 sg13g2_a21oi_1 _26076_ (.A1(net10530),
    .A2(_07634_),
    .Y(_07645_),
    .B1(_07644_));
 sg13g2_a21oi_1 _26077_ (.A1(net10530),
    .A2(_07635_),
    .Y(_07646_),
    .B1(net10504));
 sg13g2_nor2_1 _26078_ (.A(net10530),
    .B(_07635_),
    .Y(_07647_));
 sg13g2_o21ai_1 _26079_ (.B1(net10304),
    .Y(_07648_),
    .A1(_07646_),
    .A2(_07647_));
 sg13g2_o21ai_1 _26080_ (.B1(_07648_),
    .Y(_07649_),
    .A1(net10304),
    .A2(_07645_));
 sg13g2_xor2_1 _26081_ (.B(_07649_),
    .A(_08837_),
    .X(_07650_));
 sg13g2_and2_1 _26082_ (.A(net10503),
    .B(net10529),
    .X(_07651_));
 sg13g2_nand2_1 _26083_ (.Y(_07652_),
    .A(net10449),
    .B(_07651_));
 sg13g2_o21ai_1 _26084_ (.B1(_07652_),
    .Y(_07653_),
    .A1(net10529),
    .A2(net10308));
 sg13g2_a21oi_1 _26085_ (.A1(net10529),
    .A2(net10255),
    .Y(_07654_),
    .B1(net10503));
 sg13g2_a21oi_1 _26086_ (.A1(net10454),
    .A2(_07653_),
    .Y(_07655_),
    .B1(_07654_));
 sg13g2_a21o_1 _26087_ (.A2(_07650_),
    .A1(net10190),
    .B1(_07655_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[5] ));
 sg13g2_nor2_1 _26088_ (.A(_08698_),
    .B(_08706_),
    .Y(_07656_));
 sg13g2_nor2_1 _26089_ (.A(_07646_),
    .B(_07647_),
    .Y(_07657_));
 sg13g2_nor2_1 _26090_ (.A(_07651_),
    .B(_07657_),
    .Y(_07658_));
 sg13g2_nor3_1 _26091_ (.A(net10637),
    .B(_07182_),
    .C(_07658_),
    .Y(_07659_));
 sg13g2_a21oi_1 _26092_ (.A1(net10637),
    .A2(_07656_),
    .Y(_07660_),
    .B1(_07659_));
 sg13g2_xor2_1 _26093_ (.B(_07660_),
    .A(_08836_),
    .X(_07661_));
 sg13g2_nand2_1 _26094_ (.Y(_07662_),
    .A(net10449),
    .B(_07171_));
 sg13g2_o21ai_1 _26095_ (.B1(_07662_),
    .Y(_07663_),
    .A1(net10527),
    .A2(net10308));
 sg13g2_a21oi_1 _26096_ (.A1(net10527),
    .A2(net10255),
    .Y(_07664_),
    .B1(net10502));
 sg13g2_a21oi_1 _26097_ (.A1(net10454),
    .A2(_07663_),
    .Y(_07665_),
    .B1(_07664_));
 sg13g2_a21o_1 _26098_ (.A2(_07661_),
    .A1(net10190),
    .B1(_07665_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[6] ));
 sg13g2_nor2_1 _26099_ (.A(_07180_),
    .B(_07186_),
    .Y(_07666_));
 sg13g2_o21ai_1 _26100_ (.B1(net10527),
    .Y(_07667_),
    .A1(_08698_),
    .A2(_08706_));
 sg13g2_nor3_1 _26101_ (.A(net10527),
    .B(_08698_),
    .C(_08706_),
    .Y(_07668_));
 sg13g2_a21oi_1 _26102_ (.A1(net10502),
    .A2(_07667_),
    .Y(_07669_),
    .B1(_07668_));
 sg13g2_nand2_1 _26103_ (.Y(_07670_),
    .A(net10636),
    .B(_07669_));
 sg13g2_o21ai_1 _26104_ (.B1(_07670_),
    .Y(_07671_),
    .A1(net10637),
    .A2(_07666_));
 sg13g2_xnor2_1 _26105_ (.Y(_07672_),
    .A(_08834_),
    .B(_07671_));
 sg13g2_nand3_1 _26106_ (.B(net10525),
    .C(net10449),
    .A(net10501),
    .Y(_07673_));
 sg13g2_o21ai_1 _26107_ (.B1(_07673_),
    .Y(_07674_),
    .A1(net10525),
    .A2(net10308));
 sg13g2_nand2_1 _26108_ (.Y(_07675_),
    .A(net10525),
    .B(net10255));
 sg13g2_a22oi_1 _26109_ (.Y(_07676_),
    .B1(_07675_),
    .B2(_03677_),
    .A2(_07674_),
    .A1(net10454));
 sg13g2_a21o_1 _26110_ (.A2(_07672_),
    .A1(net10190),
    .B1(_07676_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[7] ));
 sg13g2_a21o_1 _26111_ (.A2(_07669_),
    .A1(net10525),
    .B1(_03677_),
    .X(_07677_));
 sg13g2_o21ai_1 _26112_ (.B1(_07677_),
    .Y(_07678_),
    .A1(net10525),
    .A2(_07669_));
 sg13g2_a21oi_1 _26113_ (.A1(net10525),
    .A2(_07666_),
    .Y(_07679_),
    .B1(net10501));
 sg13g2_nor2_1 _26114_ (.A(net10525),
    .B(_07666_),
    .Y(_07680_));
 sg13g2_nor3_1 _26115_ (.A(net10636),
    .B(_07679_),
    .C(_07680_),
    .Y(_07681_));
 sg13g2_a21oi_1 _26116_ (.A1(net10637),
    .A2(_07678_),
    .Y(_07682_),
    .B1(_07681_));
 sg13g2_xnor2_1 _26117_ (.Y(_07683_),
    .A(_08833_),
    .B(_07682_));
 sg13g2_nand3_1 _26118_ (.B(net10523),
    .C(net10449),
    .A(net10500),
    .Y(_07684_));
 sg13g2_o21ai_1 _26119_ (.B1(_07684_),
    .Y(_07685_),
    .A1(net10523),
    .A2(net10308));
 sg13g2_a21oi_1 _26120_ (.A1(net10523),
    .A2(net10255),
    .Y(_07686_),
    .B1(net10500));
 sg13g2_a21oi_1 _26121_ (.A1(net10454),
    .A2(_07685_),
    .Y(_07687_),
    .B1(_07686_));
 sg13g2_a21o_1 _26122_ (.A2(_07683_),
    .A1(net10190),
    .B1(_07687_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[8] ));
 sg13g2_nand2_1 _26123_ (.Y(_07688_),
    .A(_07196_),
    .B(_07197_));
 sg13g2_nor2_1 _26124_ (.A(net10636),
    .B(_07247_),
    .Y(_07689_));
 sg13g2_a21oi_1 _26125_ (.A1(net10636),
    .A2(_07688_),
    .Y(_07690_),
    .B1(_07689_));
 sg13g2_xnor2_1 _26126_ (.Y(_07691_),
    .A(_08830_),
    .B(_07690_));
 sg13g2_nand3_1 _26127_ (.B(net10522),
    .C(net10447),
    .A(net10499),
    .Y(_07692_));
 sg13g2_o21ai_1 _26128_ (.B1(_07692_),
    .Y(_07693_),
    .A1(net10522),
    .A2(net10307));
 sg13g2_nand2_1 _26129_ (.Y(_07694_),
    .A(net10522),
    .B(net10254));
 sg13g2_a22oi_1 _26130_ (.Y(_07695_),
    .B1(_07694_),
    .B2(_08779_),
    .A2(_07693_),
    .A1(net10453));
 sg13g2_a21o_1 _26131_ (.A2(_07691_),
    .A1(net10189),
    .B1(_07695_),
    .X(\u_ac_controller_soc_inst.u_picorv32.alu_out[9] ));
 sg13g2_dfrbp_1 _26132_ (.CLK(clknet_leaf_953_clk),
    .RESET_B(net1),
    .D(_00038_),
    .Q_N(_14013_),
    .Q(_00005_));
 sg13g2_dfrbp_1 _26133_ (.CLK(clknet_leaf_955_clk),
    .RESET_B(net2),
    .D(_00039_),
    .Q_N(_14014_),
    .Q(_00006_));
 sg13g2_dfrbp_1 _26134_ (.CLK(clknet_8_252_0_clk),
    .RESET_B(net3),
    .D(_00040_),
    .Q_N(_14015_),
    .Q(_00007_));
 sg13g2_dfrbp_1 _26135_ (.CLK(clknet_leaf_952_clk),
    .RESET_B(net4),
    .D(_00041_),
    .Q_N(_14016_),
    .Q(_00008_));
 sg13g2_dfrbp_1 _26136_ (.CLK(clknet_leaf_672_clk),
    .RESET_B(net5),
    .D(_00042_),
    .Q_N(_14017_),
    .Q(_00009_));
 sg13g2_dfrbp_1 _26137_ (.CLK(clknet_leaf_966_clk),
    .RESET_B(net6),
    .D(_00033_),
    .Q_N(_14018_),
    .Q(_00000_));
 sg13g2_dfrbp_1 _26138_ (.CLK(clknet_leaf_965_clk),
    .RESET_B(net7),
    .D(_00034_),
    .Q_N(_14019_),
    .Q(_00001_));
 sg13g2_dfrbp_1 _26139_ (.CLK(clknet_leaf_991_clk),
    .RESET_B(net8),
    .D(_00035_),
    .Q_N(_14020_),
    .Q(_00002_));
 sg13g2_dfrbp_1 _26140_ (.CLK(clknet_8_240_0_clk),
    .RESET_B(net9),
    .D(_00036_),
    .Q_N(_14021_),
    .Q(_00003_));
 sg13g2_dfrbp_1 _26141_ (.CLK(clknet_leaf_991_clk),
    .RESET_B(net10),
    .D(_00037_),
    .Q_N(_14012_),
    .Q(_00004_));
 sg13g2_buf_16 clkbuf_leaf_833_clk (.X(clknet_leaf_833_clk),
    .A(clknet_8_174_0_clk));
 sg13g2_IOPadInOut16mA sg13g2_IOPadInOut16mA_gpio_1_pad_inst (.c2p(gpio_out1),
    .c2p_en(gpio_io1_oe),
    .p2c(gpio_in1),
    .pad(gpio_1_pad));
 sg13g2_IOPadInOut16mA sg13g2_IOPadInOut16mA_gpio_2_pad_inst (.c2p(gpio_out2),
    .c2p_en(gpio_io2_oe),
    .p2c(gpio_in2),
    .pad(gpio_2_pad));
 sg13g2_IOPadInOut16mA sg13g2_IOPadInOut16mA_spi_flash_io0_pad_inst (.c2p(spi_flash_io0_do),
    .c2p_en(spi_flash_io0_oe),
    .p2c(spi_flash_io0_di),
    .pad(spi_flash_io0_pad));
 sg13g2_IOPadInOut16mA sg13g2_IOPadInOut16mA_spi_flash_io1_pad_inst (.c2p(spi_flash_io1_do),
    .c2p_en(spi_flash_io1_oe),
    .p2c(spi_flash_io1_di),
    .pad(spi_flash_io1_pad));
 sg13g2_IOPadInOut16mA sg13g2_IOPadInOut16mA_spi_flash_io2_pad_inst (.c2p(spi_flash_io2_do),
    .c2p_en(spi_flash_io2_oe),
    .p2c(spi_flash_io2_di),
    .pad(spi_flash_io2_pad));
 sg13g2_IOPadInOut16mA sg13g2_IOPadInOut16mA_spi_flash_io3_pad_inst (.c2p(spi_flash_io3_do),
    .c2p_en(spi_flash_io3_oe),
    .p2c(spi_flash_io3_di),
    .pad(spi_flash_io3_pad));
 sg13g2_IOPadIn sg13g2_IOPadIn_clk_pad_inst (.p2c(clk),
    .pad(clk_pad));
 sg13g2_IOPadIn sg13g2_IOPadIn_resetn_pad_inst (.p2c(resetn),
    .pad(resetn_pad));
 sg13g2_IOPadIn sg13g2_IOPadIn_ser_rx_pad_inst (.p2c(ser_rx),
    .pad(ser_rx_pad));
 sg13g2_IOPadIn sg13g2_IOPadIn_spi_sensor_miso_pad_inst (.p2c(spi_sensor_miso),
    .pad(spi_sensor_miso_pad));
 sg13g2_IOPadOut16mA sg13g2_IOPadOut16mA_pwm_out_pad_inst (.c2p(pwm_out),
    .pad(pwm_out_pad));
 sg13g2_IOPadOut16mA sg13g2_IOPadOut16mA_ser_tx_pad_inst (.c2p(ser_tx),
    .pad(ser_tx_pad));
 sg13g2_IOPadOut16mA sg13g2_IOPadOut16mA_spi_flash_clk_pad_inst (.c2p(spi_flash_clk),
    .pad(spi_flash_clk_pad));
 sg13g2_IOPadOut16mA sg13g2_IOPadOut16mA_spi_flash_cs_n_pad_inst (.c2p(spi_flash_cs_n),
    .pad(spi_flash_cs_n_pad));
 sg13g2_IOPadOut16mA sg13g2_IOPadOut16mA_spi_sensor_clk_pad_inst (.c2p(spi_sensor_clk),
    .pad(spi_sensor_clk_pad));
 sg13g2_IOPadOut16mA sg13g2_IOPadOut16mA_spi_sensor_cs_n_pad_inst (.c2p(spi_sensor_cs_n),
    .pad(spi_sensor_cs_n_pad));
 sg13g2_IOPadOut16mA sg13g2_IOPadOut16mA_spi_sensor_mosi_pad_inst (.c2p(spi_sensor_mosi),
    .pad(spi_sensor_mosi_pad));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.sram_wrapper_inst.ready_state$_SDFF_PP0_  (.CLK(clknet_leaf_422_clk),
    .RESET_B(net11),
    .D(_00143_),
    .Q_N(_14011_),
    .Q(\u_ac_controller_soc_inst.sram_ready ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net12),
    .D(_00144_),
    .Q_N(_00139_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10]$_SDFF_PP0_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net13),
    .D(_00145_),
    .Q_N(_14010_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[11]$_SDFF_PP0_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net14),
    .D(_00146_),
    .Q_N(_14009_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[12]$_SDFF_PP0_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net15),
    .D(_00147_),
    .Q_N(_14008_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[13]$_SDFF_PP0_  (.CLK(clknet_8_95_0_clk),
    .RESET_B(net16),
    .D(_00148_),
    .Q_N(_14007_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14]$_SDFF_PP0_  (.CLK(clknet_8_95_0_clk),
    .RESET_B(net17),
    .D(_00149_),
    .Q_N(_14006_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[15]$_SDFF_PP0_  (.CLK(clknet_leaf_343_clk),
    .RESET_B(net18),
    .D(_00150_),
    .Q_N(_14005_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[16]$_SDFF_PP0_  (.CLK(clknet_leaf_343_clk),
    .RESET_B(net19),
    .D(_00151_),
    .Q_N(_14004_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[17]$_SDFF_PP0_  (.CLK(clknet_leaf_344_clk),
    .RESET_B(net20),
    .D(_00152_),
    .Q_N(_14003_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[18]$_SDFF_PP0_  (.CLK(clknet_leaf_344_clk),
    .RESET_B(net21),
    .D(_00153_),
    .Q_N(_14002_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[19]$_SDFF_PP0_  (.CLK(clknet_8_117_0_clk),
    .RESET_B(net22),
    .D(_00154_),
    .Q_N(_14001_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[1]$_SDFF_PP0_  (.CLK(clknet_8_71_0_clk),
    .RESET_B(net23),
    .D(_00155_),
    .Q_N(_14000_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[20]$_SDFF_PP0_  (.CLK(clknet_leaf_346_clk),
    .RESET_B(net24),
    .D(_00156_),
    .Q_N(_13999_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21]$_SDFF_PP0_  (.CLK(clknet_leaf_346_clk),
    .RESET_B(net25),
    .D(_00157_),
    .Q_N(_13998_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22]$_SDFF_PP0_  (.CLK(clknet_leaf_346_clk),
    .RESET_B(net26),
    .D(_00158_),
    .Q_N(_13997_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[23]$_SDFF_PP0_  (.CLK(clknet_8_119_0_clk),
    .RESET_B(net27),
    .D(_00159_),
    .Q_N(_13996_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24]$_SDFF_PP0_  (.CLK(clknet_leaf_348_clk),
    .RESET_B(net28),
    .D(_00160_),
    .Q_N(_13995_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[25]$_SDFF_PP0_  (.CLK(clknet_leaf_348_clk),
    .RESET_B(net29),
    .D(_00161_),
    .Q_N(_13994_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26]$_SDFF_PP0_  (.CLK(clknet_leaf_359_clk),
    .RESET_B(net30),
    .D(_00162_),
    .Q_N(_13993_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[27]$_SDFF_PP0_  (.CLK(clknet_leaf_359_clk),
    .RESET_B(net31),
    .D(_00163_),
    .Q_N(_13992_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[28]$_SDFF_PP0_  (.CLK(clknet_leaf_360_clk),
    .RESET_B(net32),
    .D(_00164_),
    .Q_N(_13991_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[29]$_SDFF_PP0_  (.CLK(clknet_8_125_0_clk),
    .RESET_B(net33),
    .D(_00165_),
    .Q_N(_13990_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net34),
    .D(_00166_),
    .Q_N(_13989_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[30]$_SDFF_PP0_  (.CLK(clknet_leaf_362_clk),
    .RESET_B(net35),
    .D(_00167_),
    .Q_N(_13988_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[31]$_SDFF_PP0_  (.CLK(clknet_leaf_362_clk),
    .RESET_B(net36),
    .D(_00168_),
    .Q_N(_13987_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net37),
    .D(_00169_),
    .Q_N(_13986_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net38),
    .D(_00170_),
    .Q_N(_13985_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[5]$_SDFF_PP0_  (.CLK(clknet_8_81_0_clk),
    .RESET_B(net39),
    .D(_00171_),
    .Q_N(_13984_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[6]$_SDFF_PP0_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net40),
    .D(_00172_),
    .Q_N(_13983_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[7]$_SDFF_PP0_  (.CLK(clknet_8_84_0_clk),
    .RESET_B(net41),
    .D(_00173_),
    .Q_N(_13982_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[8]$_SDFF_PP0_  (.CLK(clknet_8_85_0_clk),
    .RESET_B(net42),
    .D(_00174_),
    .Q_N(_13981_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9]$_SDFF_PP0_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net43),
    .D(_00175_),
    .Q_N(_13980_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_416_clk),
    .RESET_B(net44),
    .D(_00176_),
    .Q_N(_13979_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[10]$_SDFFE_PN0P_  (.CLK(clknet_8_86_0_clk),
    .RESET_B(net45),
    .D(_00177_),
    .Q_N(_13978_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net46),
    .D(_00178_),
    .Q_N(_13977_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net47),
    .D(_00179_),
    .Q_N(_13976_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[13]$_SDFFE_PN0P_  (.CLK(clknet_8_93_0_clk),
    .RESET_B(net48),
    .D(_00180_),
    .Q_N(_13975_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net49),
    .D(_00181_),
    .Q_N(_13974_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net50),
    .D(_00182_),
    .Q_N(_13973_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[16]$_SDFFE_PN0P_  (.CLK(clknet_8_93_0_clk),
    .RESET_B(net51),
    .D(_00183_),
    .Q_N(_13972_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_336_clk),
    .RESET_B(net52),
    .D(_00184_),
    .Q_N(_13971_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net53),
    .D(_00185_),
    .Q_N(_13970_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_336_clk),
    .RESET_B(net54),
    .D(_00186_),
    .Q_N(_13969_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net55),
    .D(_00187_),
    .Q_N(_13968_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_333_clk),
    .RESET_B(net56),
    .D(_00188_),
    .Q_N(_13967_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net57),
    .D(_00189_),
    .Q_N(_13966_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_330_clk),
    .RESET_B(net58),
    .D(_00190_),
    .Q_N(_13965_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net59),
    .D(_00191_),
    .Q_N(_13964_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_352_clk),
    .RESET_B(net60),
    .D(_00192_),
    .Q_N(_13963_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_353_clk),
    .RESET_B(net61),
    .D(_00193_),
    .Q_N(_13962_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_353_clk),
    .RESET_B(net62),
    .D(_00194_),
    .Q_N(_13961_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[27]$_SDFFE_PN0P_  (.CLK(clknet_8_124_0_clk),
    .RESET_B(net63),
    .D(_00195_),
    .Q_N(_13960_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_372_clk),
    .RESET_B(net64),
    .D(_00196_),
    .Q_N(_13959_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_370_clk),
    .RESET_B(net65),
    .D(_00197_),
    .Q_N(_13958_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net66),
    .D(_00198_),
    .Q_N(_13957_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_370_clk),
    .RESET_B(net67),
    .D(_00199_),
    .Q_N(_13956_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_369_clk),
    .RESET_B(net68),
    .D(_00200_),
    .Q_N(_13955_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net69),
    .D(_00201_),
    .Q_N(_13954_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net70),
    .D(_00202_),
    .Q_N(_13953_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_8_83_0_clk),
    .RESET_B(net71),
    .D(_00203_),
    .Q_N(_13952_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[6]$_SDFFE_PN0P_  (.CLK(clknet_8_86_0_clk),
    .RESET_B(net72),
    .D(_00204_),
    .Q_N(_13951_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net73),
    .D(_00205_),
    .Q_N(_13950_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[8]$_SDFFE_PN0P_  (.CLK(clknet_8_84_0_clk),
    .RESET_B(net74),
    .D(_00206_),
    .Q_N(_13949_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net75),
    .D(_00207_),
    .Q_N(_13948_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in1_sync1$_SDFF_PN0_  (.CLK(clknet_leaf_820_clk),
    .RESET_B(net76),
    .D(_00208_),
    .Q_N(_13947_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in1_sync1 ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in1_sync2$_SDFF_PN0_  (.CLK(clknet_leaf_820_clk),
    .RESET_B(net77),
    .D(_00209_),
    .Q_N(_13946_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in1_sync ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in2_sync1$_SDFF_PN0_  (.CLK(clknet_8_186_0_clk),
    .RESET_B(net78),
    .D(_00210_),
    .Q_N(_13945_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in2_sync1 ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in2_sync2$_SDFF_PN0_  (.CLK(clknet_leaf_728_clk),
    .RESET_B(net79),
    .D(_00211_),
    .Q_N(_13944_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in2_sync ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_io1_oe$_SDFFE_PN0P_  (.CLK(clknet_leaf_424_clk),
    .RESET_B(net80),
    .D(_00212_),
    .Q_N(_13943_),
    .Q(gpio_io1_oe));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_io2_oe$_SDFFE_PN0P_  (.CLK(clknet_leaf_424_clk),
    .RESET_B(net81),
    .D(_00213_),
    .Q_N(_13942_),
    .Q(gpio_io2_oe));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_out1$_SDFFE_PN0P_  (.CLK(clknet_leaf_607_clk),
    .RESET_B(net82),
    .D(_00214_),
    .Q_N(_13941_),
    .Q(gpio_out1));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_out2$_SDFFE_PN0P_  (.CLK(clknet_8_178_0_clk),
    .RESET_B(net83),
    .D(_00215_),
    .Q_N(_13940_),
    .Q(gpio_out2));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_417_clk),
    .RESET_B(net84),
    .D(_00216_),
    .Q_N(_13939_),
    .Q(\u_ac_controller_soc_inst.io_rdata[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net85),
    .D(_00217_),
    .Q_N(_13938_),
    .Q(\u_ac_controller_soc_inst.io_rdata[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_329_clk),
    .RESET_B(net86),
    .D(_00218_),
    .Q_N(_13937_),
    .Q(\u_ac_controller_soc_inst.io_rdata[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net87),
    .D(_00219_),
    .Q_N(_13936_),
    .Q(\u_ac_controller_soc_inst.io_rdata[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_329_clk),
    .RESET_B(net88),
    .D(_00220_),
    .Q_N(_13935_),
    .Q(\u_ac_controller_soc_inst.io_rdata[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_401_clk),
    .RESET_B(net89),
    .D(_00221_),
    .Q_N(_13934_),
    .Q(\u_ac_controller_soc_inst.io_rdata[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net90),
    .D(_00222_),
    .Q_N(_13933_),
    .Q(\u_ac_controller_soc_inst.io_rdata[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_330_clk),
    .RESET_B(net91),
    .D(_00223_),
    .Q_N(_13932_),
    .Q(\u_ac_controller_soc_inst.io_rdata[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[17]$_SDFFE_PN0P_  (.CLK(clknet_8_115_0_clk),
    .RESET_B(net92),
    .D(_00224_),
    .Q_N(_13931_),
    .Q(\u_ac_controller_soc_inst.io_rdata[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_367_clk),
    .RESET_B(net93),
    .D(_00225_),
    .Q_N(_13930_),
    .Q(\u_ac_controller_soc_inst.io_rdata[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_367_clk),
    .RESET_B(net94),
    .D(_00226_),
    .Q_N(_13929_),
    .Q(\u_ac_controller_soc_inst.io_rdata[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net95),
    .D(_00227_),
    .Q_N(_13928_),
    .Q(\u_ac_controller_soc_inst.io_rdata[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_331_clk),
    .RESET_B(net96),
    .D(_00228_),
    .Q_N(_13927_),
    .Q(\u_ac_controller_soc_inst.io_rdata[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_331_clk),
    .RESET_B(net97),
    .D(_00229_),
    .Q_N(_13926_),
    .Q(\u_ac_controller_soc_inst.io_rdata[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_401_clk),
    .RESET_B(net98),
    .D(_00230_),
    .Q_N(_13925_),
    .Q(\u_ac_controller_soc_inst.io_rdata[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_372_clk),
    .RESET_B(net99),
    .D(_00231_),
    .Q_N(_13924_),
    .Q(\u_ac_controller_soc_inst.io_rdata[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_374_clk),
    .RESET_B(net100),
    .D(_00232_),
    .Q_N(_13923_),
    .Q(\u_ac_controller_soc_inst.io_rdata[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_372_clk),
    .RESET_B(net101),
    .D(_00233_),
    .Q_N(_13922_),
    .Q(\u_ac_controller_soc_inst.io_rdata[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_368_clk),
    .RESET_B(net102),
    .D(_00234_),
    .Q_N(_13921_),
    .Q(\u_ac_controller_soc_inst.io_rdata[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_367_clk),
    .RESET_B(net103),
    .D(_00235_),
    .Q_N(_13920_),
    .Q(\u_ac_controller_soc_inst.io_rdata[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_371_clk),
    .RESET_B(net104),
    .D(_00236_),
    .Q_N(_13919_),
    .Q(\u_ac_controller_soc_inst.io_rdata[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_371_clk),
    .RESET_B(net105),
    .D(_00237_),
    .Q_N(_13918_),
    .Q(\u_ac_controller_soc_inst.io_rdata[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net106),
    .D(_00238_),
    .Q_N(_13917_),
    .Q(\u_ac_controller_soc_inst.io_rdata[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_368_clk),
    .RESET_B(net107),
    .D(_00239_),
    .Q_N(_13916_),
    .Q(\u_ac_controller_soc_inst.io_rdata[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_369_clk),
    .RESET_B(net108),
    .D(_00240_),
    .Q_N(_13915_),
    .Q(\u_ac_controller_soc_inst.io_rdata[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net109),
    .D(_00241_),
    .Q_N(_13914_),
    .Q(\u_ac_controller_soc_inst.io_rdata[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net110),
    .D(_00242_),
    .Q_N(_13913_),
    .Q(\u_ac_controller_soc_inst.io_rdata[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net111),
    .D(_00243_),
    .Q_N(_13912_),
    .Q(\u_ac_controller_soc_inst.io_rdata[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net112),
    .D(_00244_),
    .Q_N(_13911_),
    .Q(\u_ac_controller_soc_inst.io_rdata[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net113),
    .D(_00245_),
    .Q_N(_13910_),
    .Q(\u_ac_controller_soc_inst.io_rdata[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net114),
    .D(_00246_),
    .Q_N(_13909_),
    .Q(\u_ac_controller_soc_inst.io_rdata[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net115),
    .D(_00247_),
    .Q_N(_13908_),
    .Q(\u_ac_controller_soc_inst.io_rdata[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_ready$_SDFF_PN0_  (.CLK(clknet_leaf_419_clk),
    .RESET_B(net116),
    .D(_00248_),
    .Q_N(_13907_),
    .Q(\u_ac_controller_soc_inst.io_ready ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net117),
    .D(_00249_),
    .Q_N(_13906_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net118),
    .D(_00250_),
    .Q_N(_13905_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net119),
    .D(_00251_),
    .Q_N(_13904_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[12]$_SDFFE_PN0P_  (.CLK(clknet_8_86_0_clk),
    .RESET_B(net120),
    .D(_00252_),
    .Q_N(_13903_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net121),
    .D(_00253_),
    .Q_N(_13902_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_338_clk),
    .RESET_B(net122),
    .D(_00254_),
    .Q_N(_13901_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net123),
    .D(_00255_),
    .Q_N(_13900_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_335_clk),
    .RESET_B(net124),
    .D(_00256_),
    .Q_N(_13899_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_342_clk),
    .RESET_B(net125),
    .D(_00257_),
    .Q_N(_13898_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_341_clk),
    .RESET_B(net126),
    .D(_00258_),
    .Q_N(_13897_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_341_clk),
    .RESET_B(net127),
    .D(_00259_),
    .Q_N(_13896_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net128),
    .D(_00260_),
    .Q_N(_13895_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_334_clk),
    .RESET_B(net129),
    .D(_00261_),
    .Q_N(_13894_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_334_clk),
    .RESET_B(net130),
    .D(_00262_),
    .Q_N(_13893_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_350_clk),
    .RESET_B(net131),
    .D(_00263_),
    .Q_N(_13892_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_350_clk),
    .RESET_B(net132),
    .D(_00264_),
    .Q_N(_13891_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_355_clk),
    .RESET_B(net133),
    .D(_00265_),
    .Q_N(_13890_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_349_clk),
    .RESET_B(net134),
    .D(_00266_),
    .Q_N(_13889_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_358_clk),
    .RESET_B(net135),
    .D(_00267_),
    .Q_N(_13888_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_355_clk),
    .RESET_B(net136),
    .D(_00268_),
    .Q_N(_13887_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_357_clk),
    .RESET_B(net137),
    .D(_00269_),
    .Q_N(_13886_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_356_clk),
    .RESET_B(net138),
    .D(_00270_),
    .Q_N(_13885_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[2]$_SDFFE_PN0P_  (.CLK(clknet_8_82_0_clk),
    .RESET_B(net139),
    .D(_00271_),
    .Q_N(_13884_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_365_clk),
    .RESET_B(net140),
    .D(_00272_),
    .Q_N(_13883_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[31]$_SDFFE_PN0P_  (.CLK(clknet_8_124_0_clk),
    .RESET_B(net141),
    .D(_00273_),
    .Q_N(_13882_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net142),
    .D(_00274_),
    .Q_N(_13881_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net143),
    .D(_00275_),
    .Q_N(_13880_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net144),
    .D(_00276_),
    .Q_N(_13879_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[6]$_SDFFE_PN0P_  (.CLK(clknet_8_84_0_clk),
    .RESET_B(net145),
    .D(_00277_),
    .Q_N(_13878_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net146),
    .D(_00278_),
    .Q_N(_13877_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net147),
    .D(_00279_),
    .Q_N(_13876_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[9]$_SDFFE_PN0P_  (.CLK(clknet_8_85_0_clk),
    .RESET_B(net148),
    .D(_00280_),
    .Q_N(_13875_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_enable$_SDFFE_PN1P_  (.CLK(clknet_8_91_0_clk),
    .RESET_B(net149),
    .D(_00281_),
    .Q_N(_13874_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_enable ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_out$_SDFF_PN0_  (.CLK(clknet_leaf_360_clk),
    .RESET_B(net150),
    .D(_00282_),
    .Q_N(_13873_),
    .Q(pwm_out));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net151),
    .D(_00283_),
    .Q_N(_13872_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net152),
    .D(_00284_),
    .Q_N(_13871_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[11]$_SDFFE_PN0P_  (.CLK(clknet_8_87_0_clk),
    .RESET_B(net153),
    .D(_00285_),
    .Q_N(_13870_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net154),
    .D(_00286_),
    .Q_N(_13869_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_337_clk),
    .RESET_B(net155),
    .D(_00287_),
    .Q_N(_13868_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_338_clk),
    .RESET_B(net156),
    .D(_00288_),
    .Q_N(_13867_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[15]$_SDFFE_PN0P_  (.CLK(clknet_8_95_0_clk),
    .RESET_B(net157),
    .D(_00289_),
    .Q_N(_13866_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_335_clk),
    .RESET_B(net158),
    .D(_00290_),
    .Q_N(_13865_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_340_clk),
    .RESET_B(net159),
    .D(_00291_),
    .Q_N(_13864_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_342_clk),
    .RESET_B(net160),
    .D(_00292_),
    .Q_N(_13863_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_340_clk),
    .RESET_B(net161),
    .D(_00293_),
    .Q_N(_13862_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[1]$_SDFFE_PN0P_  (.CLK(clknet_8_83_0_clk),
    .RESET_B(net162),
    .D(_00294_),
    .Q_N(_13861_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_333_clk),
    .RESET_B(net163),
    .D(_00295_),
    .Q_N(_13860_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_350_clk),
    .RESET_B(net164),
    .D(_00296_),
    .Q_N(_13859_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_332_clk),
    .RESET_B(net165),
    .D(_00297_),
    .Q_N(_13858_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[23]$_SDFFE_PN0P_  (.CLK(clknet_8_118_0_clk),
    .RESET_B(net166),
    .D(_00298_),
    .Q_N(_13857_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_352_clk),
    .RESET_B(net167),
    .D(_00299_),
    .Q_N(_13856_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_349_clk),
    .RESET_B(net168),
    .D(_00300_),
    .Q_N(_13855_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_358_clk),
    .RESET_B(net169),
    .D(_00301_),
    .Q_N(_13854_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_355_clk),
    .RESET_B(net170),
    .D(_00302_),
    .Q_N(_13853_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_356_clk),
    .RESET_B(net171),
    .D(_00303_),
    .Q_N(_13852_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_357_clk),
    .RESET_B(net172),
    .D(_00304_),
    .Q_N(_13851_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net173),
    .D(_00305_),
    .Q_N(_13850_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_365_clk),
    .RESET_B(net174),
    .D(_00306_),
    .Q_N(_13849_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_365_clk),
    .RESET_B(net175),
    .D(_00307_),
    .Q_N(_13848_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net176),
    .D(_00308_),
    .Q_N(_13847_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[4]$_SDFFE_PN0P_  (.CLK(clknet_8_81_0_clk),
    .RESET_B(net177),
    .D(_00309_),
    .Q_N(_13846_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net178),
    .D(_00310_),
    .Q_N(_13845_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net179),
    .D(_00311_),
    .Q_N(_13844_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[7]$_SDFFE_PN0P_  (.CLK(clknet_8_84_0_clk),
    .RESET_B(net180),
    .D(_00312_),
    .Q_N(_13843_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net181),
    .D(_00313_),
    .Q_N(_13842_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net182),
    .D(_00314_),
    .Q_N(_13841_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_433_clk),
    .RESET_B(net183),
    .D(_00315_),
    .Q_N(_13840_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_432_clk),
    .RESET_B(net184),
    .D(_00316_),
    .Q_N(_13839_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_432_clk),
    .RESET_B(net185),
    .D(_00317_),
    .Q_N(_13838_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3]$_SDFFE_PN0P_  (.CLK(clknet_8_103_0_clk),
    .RESET_B(net186),
    .D(_00318_),
    .Q_N(_13837_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_430_clk),
    .RESET_B(net187),
    .D(_00319_),
    .Q_N(_13836_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_430_clk),
    .RESET_B(net188),
    .D(_00320_),
    .Q_N(_13835_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_410_clk),
    .RESET_B(net189),
    .D(_00321_),
    .Q_N(_13834_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_396_clk),
    .RESET_B(net190),
    .D(_00322_),
    .Q_N(_13833_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_395_clk),
    .RESET_B(net191),
    .D(_00323_),
    .Q_N(_13832_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_397_clk),
    .RESET_B(net192),
    .D(_00324_),
    .Q_N(_13831_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_397_clk),
    .RESET_B(net193),
    .D(_00325_),
    .Q_N(_13830_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[14]$_SDFFE_PN0P_  (.CLK(clknet_8_109_0_clk),
    .RESET_B(net194),
    .D(_00326_),
    .Q_N(_13829_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_384_clk),
    .RESET_B(net195),
    .D(_00327_),
    .Q_N(_13828_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[16]$_SDFFE_PN0P_  (.CLK(clknet_8_122_0_clk),
    .RESET_B(net196),
    .D(_00328_),
    .Q_N(_13827_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_530_clk),
    .RESET_B(net197),
    .D(_00329_),
    .Q_N(_13826_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_530_clk),
    .RESET_B(net198),
    .D(_00330_),
    .Q_N(_13825_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_529_clk),
    .RESET_B(net199),
    .D(_00331_),
    .Q_N(_13824_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_410_clk),
    .RESET_B(net200),
    .D(_00332_),
    .Q_N(_13823_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_384_clk),
    .RESET_B(net201),
    .D(_00333_),
    .Q_N(_13822_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_385_clk),
    .RESET_B(net202),
    .D(_00334_),
    .Q_N(_13821_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_386_clk),
    .RESET_B(net203),
    .D(_00335_),
    .Q_N(_13820_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[23]$_SDFFE_PN0P_  (.CLK(clknet_8_111_0_clk),
    .RESET_B(net204),
    .D(_00336_),
    .Q_N(_13819_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_393_clk),
    .RESET_B(net205),
    .D(_00337_),
    .Q_N(_13818_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_393_clk),
    .RESET_B(net206),
    .D(_00338_),
    .Q_N(_13817_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_391_clk),
    .RESET_B(net207),
    .D(_00339_),
    .Q_N(_13816_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_389_clk),
    .RESET_B(net208),
    .D(_00340_),
    .Q_N(_13815_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_386_clk),
    .RESET_B(net209),
    .D(_00341_),
    .Q_N(_13814_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_391_clk),
    .RESET_B(net210),
    .D(_00342_),
    .Q_N(_13813_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_412_clk),
    .RESET_B(net211),
    .D(_00343_),
    .Q_N(_13812_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_389_clk),
    .RESET_B(net212),
    .D(_00344_),
    .Q_N(_13811_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_385_clk),
    .RESET_B(net213),
    .D(_00345_),
    .Q_N(_00128_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_419_clk),
    .RESET_B(net214),
    .D(_00346_),
    .Q_N(_13810_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_411_clk),
    .RESET_B(net215),
    .D(_00347_),
    .Q_N(_13809_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[5]$_SDFFE_PN0P_  (.CLK(clknet_8_101_0_clk),
    .RESET_B(net216),
    .D(_00348_),
    .Q_N(_13808_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_411_clk),
    .RESET_B(net217),
    .D(_00349_),
    .Q_N(_13807_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_409_clk),
    .RESET_B(net218),
    .D(_00350_),
    .Q_N(_13806_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_409_clk),
    .RESET_B(net219),
    .D(_00351_),
    .Q_N(_13805_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_408_clk),
    .RESET_B(net220),
    .D(_00352_),
    .Q_N(_13804_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_rdata[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net221),
    .D(_00353_),
    .Q_N(_13803_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[10]$_SDFFE_PN0P_  (.CLK(clknet_8_21_0_clk),
    .RESET_B(net222),
    .D(_00354_),
    .Q_N(_13802_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net223),
    .D(_00355_),
    .Q_N(_13801_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net224),
    .D(_00356_),
    .Q_N(_13800_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[13]$_SDFFE_PN0P_  (.CLK(clknet_8_66_0_clk),
    .RESET_B(net225),
    .D(_00357_),
    .Q_N(_13799_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net226),
    .D(_00358_),
    .Q_N(_13798_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net227),
    .D(_00359_),
    .Q_N(_13797_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[16]$_SDFFE_PN0P_  (.CLK(clknet_8_20_0_clk),
    .RESET_B(net228),
    .D(_00360_),
    .Q_N(_13796_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net229),
    .D(_00361_),
    .Q_N(_13795_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[18]$_SDFFE_PN0P_  (.CLK(clknet_8_64_0_clk),
    .RESET_B(net230),
    .D(_00362_),
    .Q_N(_13794_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net231),
    .D(_00363_),
    .Q_N(_13793_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net232),
    .D(_00364_),
    .Q_N(_13792_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[20]$_SDFFE_PN0P_  (.CLK(clknet_8_21_0_clk),
    .RESET_B(net233),
    .D(_00365_),
    .Q_N(_13791_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net234),
    .D(_00366_),
    .Q_N(_13790_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net235),
    .D(_00367_),
    .Q_N(_13789_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net236),
    .D(_00368_),
    .Q_N(_13788_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[24]$_SDFFE_PN0P_  (.CLK(clknet_8_72_0_clk),
    .RESET_B(net237),
    .D(_00369_),
    .Q_N(_13787_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net238),
    .D(_00370_),
    .Q_N(_13786_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net239),
    .D(_00371_),
    .Q_N(_13785_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net240),
    .D(_00372_),
    .Q_N(_13784_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net241),
    .D(_00373_),
    .Q_N(_13783_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net242),
    .D(_00374_),
    .Q_N(_13782_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[2]$_SDFFE_PN0P_  (.CLK(clknet_8_75_0_clk),
    .RESET_B(net243),
    .D(_00375_),
    .Q_N(_13781_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net244),
    .D(_00376_),
    .Q_N(_13780_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net245),
    .D(_00377_),
    .Q_N(_13779_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[32]$_SDFFE_PN0P_  (.CLK(clknet_8_79_0_clk),
    .RESET_B(net246),
    .D(_00378_),
    .Q_N(_13778_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[32] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net247),
    .D(_00379_),
    .Q_N(_13777_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[33] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[34]$_SDFFE_PP0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net248),
    .D(_00380_),
    .Q_N(_13776_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[34] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[35]$_SDFFE_PP0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net249),
    .D(_00381_),
    .Q_N(_13775_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[35] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net250),
    .D(_00382_),
    .Q_N(_13774_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[36] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net251),
    .D(_00383_),
    .Q_N(_13773_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[37] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net252),
    .D(_00384_),
    .Q_N(_13772_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[38] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net253),
    .D(_00385_),
    .Q_N(_13771_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[39] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[3]$_SDFFE_PN0P_  (.CLK(clknet_8_73_0_clk),
    .RESET_B(net254),
    .D(_00386_),
    .Q_N(_13770_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net255),
    .D(_00387_),
    .Q_N(_13769_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net256),
    .D(_00388_),
    .Q_N(_13768_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net257),
    .D(_00389_),
    .Q_N(_13767_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net258),
    .D(_00390_),
    .Q_N(_13766_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[8]$_SDFFE_PN0P_  (.CLK(clknet_8_66_0_clk),
    .RESET_B(net259),
    .D(_00391_),
    .Q_N(_13765_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net260),
    .D(_00392_),
    .Q_N(_13764_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.spi_clk_reg$_SDFF_PN0_  (.CLK(clknet_leaf_429_clk),
    .RESET_B(net261),
    .D(_00393_),
    .Q_N(_00043_),
    .Q(spi_sensor_clk));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.spi_cs_n_reg$_SDFFE_PP1P_  (.CLK(clknet_leaf_428_clk),
    .RESET_B(net262),
    .D(_00394_),
    .Q_N(_00103_),
    .Q(spi_sensor_cs_n));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.spi_sensor_ready_reg$_SDFF_PN0_  (.CLK(clknet_leaf_429_clk),
    .RESET_B(net263),
    .D(_00395_),
    .Q_N(_13763_),
    .Q(\u_ac_controller_soc_inst.spi_sensor_ready ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[3]$_SDFF_PN0_  (.CLK(clknet_leaf_421_clk),
    .RESET_B(net264),
    .D(_00396_),
    .Q_N(_13762_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[4]$_SDFF_PN1_  (.CLK(clknet_leaf_422_clk),
    .RESET_B(net265),
    .D(_00397_),
    .Q_N(_13761_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[5]$_SDFF_PN0_  (.CLK(clknet_leaf_421_clk),
    .RESET_B(net266),
    .D(_00398_),
    .Q_N(_13760_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_420_clk),
    .RESET_B(net267),
    .D(_00399_),
    .Q_N(_13759_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_420_clk),
    .RESET_B(net268),
    .D(_00400_),
    .Q_N(_13758_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[0]$_SDFFE_PP0P_  (.CLK(clknet_8_23_0_clk),
    .RESET_B(net269),
    .D(_00401_),
    .Q_N(_00137_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[1]$_SDFFE_PP0P_  (.CLK(clknet_8_23_0_clk),
    .RESET_B(net270),
    .D(_00402_),
    .Q_N(_13757_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2]$_SDFFE_PP0P_  (.CLK(clknet_8_22_0_clk),
    .RESET_B(net271),
    .D(_00403_),
    .Q_N(_00136_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net272),
    .D(_00404_),
    .Q_N(_00135_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[10]$_SDFFE_PP0P_  (.CLK(clknet_8_16_0_clk),
    .RESET_B(net273),
    .D(_00405_),
    .Q_N(_13756_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net274),
    .D(_00406_),
    .Q_N(_13755_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net275),
    .D(_00407_),
    .Q_N(_13754_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net276),
    .D(_00408_),
    .Q_N(_13753_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net277),
    .D(_00409_),
    .Q_N(_13752_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net278),
    .D(_00410_),
    .Q_N(_13751_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net279),
    .D(_00411_),
    .Q_N(_13750_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net280),
    .D(_00412_),
    .Q_N(_13749_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net281),
    .D(_00413_),
    .Q_N(_13748_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net282),
    .D(_00414_),
    .Q_N(_13747_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net283),
    .D(_00415_),
    .Q_N(_13746_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[20]$_SDFFE_PP0P_  (.CLK(clknet_8_5_0_clk),
    .RESET_B(net284),
    .D(_00416_),
    .Q_N(_13745_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[21]$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net285),
    .D(_00417_),
    .Q_N(_13744_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22]$_SDFFE_PP0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net286),
    .D(_00418_),
    .Q_N(_13743_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[23]$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net287),
    .D(_00419_),
    .Q_N(_13742_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[24]$_SDFFE_PP0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net288),
    .D(_00420_),
    .Q_N(_13741_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[25]$_SDFFE_PP0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net289),
    .D(_00421_),
    .Q_N(_13740_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[26]$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net290),
    .D(_00422_),
    .Q_N(_13739_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[27]$_SDFFE_PP0P_  (.CLK(clknet_8_7_0_clk),
    .RESET_B(net291),
    .D(_00423_),
    .Q_N(_13738_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[28]$_SDFFE_PP0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net292),
    .D(_00424_),
    .Q_N(_13737_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[29]$_SDFFE_PP0P_  (.CLK(clknet_8_6_0_clk),
    .RESET_B(net293),
    .D(_00425_),
    .Q_N(_13736_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net294),
    .D(_00426_),
    .Q_N(_13735_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[30]$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net295),
    .D(_00427_),
    .Q_N(_13734_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[31]$_SDFFE_PP0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net296),
    .D(_00428_),
    .Q_N(_13733_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net297),
    .D(_00429_),
    .Q_N(_13732_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net298),
    .D(_00430_),
    .Q_N(_13731_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net299),
    .D(_00431_),
    .Q_N(_13730_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net300),
    .D(_00432_),
    .Q_N(_13729_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[7]$_SDFFE_PP0P_  (.CLK(clknet_8_17_0_clk),
    .RESET_B(net301),
    .D(_00433_),
    .Q_N(_13728_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[8]$_SDFFE_PP0P_  (.CLK(clknet_8_17_0_clk),
    .RESET_B(net302),
    .D(_00434_),
    .Q_N(_13727_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net303),
    .D(_00435_),
    .Q_N(_13726_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net304),
    .D(_00436_),
    .Q_N(_13725_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net305),
    .D(_00437_),
    .Q_N(_13724_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net306),
    .D(_00438_),
    .Q_N(_13723_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net307),
    .D(_00439_),
    .Q_N(_13722_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net308),
    .D(_00440_),
    .Q_N(_13721_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net309),
    .D(_00441_),
    .Q_N(_13720_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[6]$_SDFFE_PN0P_  (.CLK(clknet_8_88_0_clk),
    .RESET_B(net310),
    .D(_00442_),
    .Q_N(_13719_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net311),
    .D(_00443_),
    .Q_N(_13718_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_416_clk),
    .RESET_B(net312),
    .D(_00444_),
    .Q_N(_13717_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync1$_SDFF_PN1_  (.CLK(clknet_8_237_0_clk),
    .RESET_B(net313),
    .D(_00445_),
    .Q_N(_13716_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync1 ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync2$_SDFF_PN1_  (.CLK(clknet_leaf_613_clk),
    .RESET_B(net314),
    .D(_00446_),
    .Q_N(_13715_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_tx$_SDFFE_PP1P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net315),
    .D(_00447_),
    .Q_N(_13714_),
    .Q(ser_tx));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.start_bit$_SDFFE_PP0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net316),
    .D(_00448_),
    .Q_N(_13713_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.start_bit ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.stop_bit$_SDFFE_PP0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net317),
    .D(_00449_),
    .Q_N(_00096_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.stop_bit ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_417_clk),
    .RESET_B(net318),
    .D(_00450_),
    .Q_N(_13712_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net319),
    .D(_00451_),
    .Q_N(_13711_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_416_clk),
    .RESET_B(net320),
    .D(_00452_),
    .Q_N(_13710_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net321),
    .D(_00453_),
    .Q_N(_13709_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[4]$_SDFFE_PN0P_  (.CLK(clknet_8_89_0_clk),
    .RESET_B(net322),
    .D(_00454_),
    .Q_N(_13708_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net323),
    .D(_00455_),
    .Q_N(_13707_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net324),
    .D(_00456_),
    .Q_N(_13706_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net325),
    .D(_00457_),
    .Q_N(_13705_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[8]$_SDFFE_PN0P_  (.CLK(clknet_8_90_0_clk),
    .RESET_B(net326),
    .D(_00458_),
    .Q_N(_13704_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_ready$_SDFF_PN0_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net327),
    .D(_00459_),
    .Q_N(_13703_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_ready ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net328),
    .D(_00460_),
    .Q_N(_13702_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net329),
    .D(_00461_),
    .Q_N(_13701_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net330),
    .D(_00462_),
    .Q_N(_13700_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net331),
    .D(_00463_),
    .Q_N(_13699_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net332),
    .D(_00464_),
    .Q_N(_13698_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net333),
    .D(_00465_),
    .Q_N(_13697_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[12]$_SDFFE_PN0P_  (.CLK(clknet_8_16_0_clk),
    .RESET_B(net334),
    .D(_00466_),
    .Q_N(_13696_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[13]$_SDFFE_PN0P_  (.CLK(clknet_8_16_0_clk),
    .RESET_B(net335),
    .D(_00467_),
    .Q_N(_13695_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net336),
    .D(_00468_),
    .Q_N(_13694_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net337),
    .D(_00469_),
    .Q_N(_13693_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net338),
    .D(_00470_),
    .Q_N(_13692_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[17]$_SDFFE_PN0P_  (.CLK(clknet_8_4_0_clk),
    .RESET_B(net339),
    .D(_00471_),
    .Q_N(_13691_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net340),
    .D(_00472_),
    .Q_N(_13690_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net341),
    .D(_00473_),
    .Q_N(_13689_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net342),
    .D(_00474_),
    .Q_N(_13688_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net343),
    .D(_00475_),
    .Q_N(_13687_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net344),
    .D(_00476_),
    .Q_N(_13686_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net345),
    .D(_00477_),
    .Q_N(_13685_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net346),
    .D(_00478_),
    .Q_N(_13684_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net347),
    .D(_00479_),
    .Q_N(_13683_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net348),
    .D(_00480_),
    .Q_N(_13682_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net349),
    .D(_00481_),
    .Q_N(_13681_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net350),
    .D(_00482_),
    .Q_N(_13680_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net351),
    .D(_00483_),
    .Q_N(_13679_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[29]$_SDFFE_PN0P_  (.CLK(clknet_8_13_0_clk),
    .RESET_B(net352),
    .D(_00484_),
    .Q_N(_13678_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net353),
    .D(_00485_),
    .Q_N(_13677_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net354),
    .D(_00486_),
    .Q_N(_13676_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net355),
    .D(_00487_),
    .Q_N(_13675_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net356),
    .D(_00488_),
    .Q_N(_13674_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net357),
    .D(_00489_),
    .Q_N(_13673_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[5]$_SDFFE_PN0P_  (.CLK(clknet_8_16_0_clk),
    .RESET_B(net358),
    .D(_00490_),
    .Q_N(_13672_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net359),
    .D(_00491_),
    .Q_N(_13671_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net360),
    .D(_00492_),
    .Q_N(_13670_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net361),
    .D(_00493_),
    .Q_N(_13669_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[9]$_SDFFE_PN0P_  (.CLK(clknet_8_20_0_clk),
    .RESET_B(net362),
    .D(_00494_),
    .Q_N(_13668_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_done$_SDFF_PN0_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net363),
    .D(_00495_),
    .Q_N(_13667_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_done ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout$_SDFF_PP0_  (.CLK(clknet_8_123_0_clk),
    .RESET_B(net364),
    .D(_00496_),
    .Q_N(_00111_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_532_clk),
    .RESET_B(net365),
    .D(_00497_),
    .Q_N(_13666_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[10]$_SDFFE_PN0P_  (.CLK(clknet_8_127_0_clk),
    .RESET_B(net366),
    .D(_00498_),
    .Q_N(_13665_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[11]$_SDFFE_PN0P_  (.CLK(clknet_8_127_0_clk),
    .RESET_B(net367),
    .D(_00499_),
    .Q_N(_13664_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_547_clk),
    .RESET_B(net368),
    .D(_00500_),
    .Q_N(_13663_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_546_clk),
    .RESET_B(net369),
    .D(_00501_),
    .Q_N(_13662_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_547_clk),
    .RESET_B(net370),
    .D(_00502_),
    .Q_N(_13661_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[15]$_SDFFE_PN0P_  (.CLK(clknet_8_127_0_clk),
    .RESET_B(net371),
    .D(_00503_),
    .Q_N(_13660_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_550_clk),
    .RESET_B(net372),
    .D(_00504_),
    .Q_N(_13659_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_550_clk),
    .RESET_B(net373),
    .D(_00505_),
    .Q_N(_13658_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_552_clk),
    .RESET_B(net374),
    .D(_00506_),
    .Q_N(_13657_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_552_clk),
    .RESET_B(net375),
    .D(_00507_),
    .Q_N(_13656_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_541_clk),
    .RESET_B(net376),
    .D(_00508_),
    .Q_N(_13655_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_553_clk),
    .RESET_B(net377),
    .D(_00509_),
    .Q_N(_13654_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[21]$_SDFFE_PN0P_  (.CLK(clknet_8_213_0_clk),
    .RESET_B(net378),
    .D(_00510_),
    .Q_N(_13653_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_546_clk),
    .RESET_B(net379),
    .D(_00511_),
    .Q_N(_13652_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_553_clk),
    .RESET_B(net380),
    .D(_00512_),
    .Q_N(_13651_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_553_clk),
    .RESET_B(net381),
    .D(_00513_),
    .Q_N(_13650_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_554_clk),
    .RESET_B(net382),
    .D(_00514_),
    .Q_N(_13649_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_554_clk),
    .RESET_B(net383),
    .D(_00515_),
    .Q_N(_13648_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_539_clk),
    .RESET_B(net384),
    .D(_00516_),
    .Q_N(_13647_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[28]$_SDFFE_PN0P_  (.CLK(clknet_8_123_0_clk),
    .RESET_B(net385),
    .D(_00517_),
    .Q_N(_13646_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_539_clk),
    .RESET_B(net386),
    .D(_00518_),
    .Q_N(_13645_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_541_clk),
    .RESET_B(net387),
    .D(_00519_),
    .Q_N(_13644_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_539_clk),
    .RESET_B(net388),
    .D(_00520_),
    .Q_N(_13643_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_540_clk),
    .RESET_B(net389),
    .D(_00521_),
    .Q_N(_13642_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_540_clk),
    .RESET_B(net390),
    .D(_00522_),
    .Q_N(_13641_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_543_clk),
    .RESET_B(net391),
    .D(_00523_),
    .Q_N(_13640_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_543_clk),
    .RESET_B(net392),
    .D(_00524_),
    .Q_N(_13639_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_8_126_0_clk),
    .RESET_B(net393),
    .D(_00525_),
    .Q_N(_13638_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_366_clk),
    .RESET_B(net394),
    .D(_00526_),
    .Q_N(_13637_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_366_clk),
    .RESET_B(net395),
    .D(_00527_),
    .Q_N(_13636_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[9]$_SDFFE_PN0P_  (.CLK(clknet_8_126_0_clk),
    .RESET_B(net396),
    .D(_00528_),
    .Q_N(_13635_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfering$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net397),
    .D(_00529_),
    .Q_N(_00097_),
    .Q(\u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfering ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[0]$_DFF_P_  (.CLK(clknet_leaf_470_clk),
    .RESET_B(net398),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[0] ),
    .Q_N(_14022_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[10]$_DFF_P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net399),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[10] ),
    .Q_N(_14023_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[11]$_DFF_P_  (.CLK(clknet_leaf_660_clk),
    .RESET_B(net400),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[11] ),
    .Q_N(_14024_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[12]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net401),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[12] ),
    .Q_N(_14025_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[13]$_DFF_P_  (.CLK(clknet_leaf_660_clk),
    .RESET_B(net402),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[13] ),
    .Q_N(_14026_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[14]$_DFF_P_  (.CLK(clknet_leaf_658_clk),
    .RESET_B(net403),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[14] ),
    .Q_N(_14027_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[15]$_DFF_P_  (.CLK(clknet_8_246_0_clk),
    .RESET_B(net404),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[15] ),
    .Q_N(_14028_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[16]$_DFF_P_  (.CLK(clknet_leaf_654_clk),
    .RESET_B(net405),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[16] ),
    .Q_N(_14029_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[17]$_DFF_P_  (.CLK(clknet_leaf_654_clk),
    .RESET_B(net406),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[17] ),
    .Q_N(_14030_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[18]$_DFF_P_  (.CLK(clknet_leaf_653_clk),
    .RESET_B(net407),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[18] ),
    .Q_N(_14031_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[19]$_DFF_P_  (.CLK(clknet_8_253_0_clk),
    .RESET_B(net408),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[19] ),
    .Q_N(_14032_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[1]$_DFF_P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net409),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[1] ),
    .Q_N(_14033_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[20]$_DFF_P_  (.CLK(clknet_leaf_608_clk),
    .RESET_B(net410),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[20] ),
    .Q_N(_14034_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[21]$_DFF_P_  (.CLK(clknet_leaf_641_clk),
    .RESET_B(net411),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[21] ),
    .Q_N(_14035_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[22]$_DFF_P_  (.CLK(clknet_leaf_606_clk),
    .RESET_B(net412),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[22] ),
    .Q_N(_14036_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[23]$_DFF_P_  (.CLK(clknet_leaf_606_clk),
    .RESET_B(net413),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[23] ),
    .Q_N(_14037_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[24]$_DFF_P_  (.CLK(clknet_leaf_606_clk),
    .RESET_B(net414),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[24] ),
    .Q_N(_14038_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[25]$_DFF_P_  (.CLK(clknet_leaf_604_clk),
    .RESET_B(net415),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[25] ),
    .Q_N(_14039_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[26]$_DFF_P_  (.CLK(clknet_leaf_605_clk),
    .RESET_B(net416),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[26] ),
    .Q_N(_14040_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[27]$_DFF_P_  (.CLK(clknet_leaf_605_clk),
    .RESET_B(net417),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[27] ),
    .Q_N(_14041_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[28]$_DFF_P_  (.CLK(clknet_leaf_607_clk),
    .RESET_B(net418),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[28] ),
    .Q_N(_14042_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[29]$_DFF_P_  (.CLK(clknet_leaf_608_clk),
    .RESET_B(net419),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[29] ),
    .Q_N(_14043_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[2]$_DFF_P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net420),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[2] ),
    .Q_N(_14044_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[30]$_DFF_P_  (.CLK(clknet_leaf_607_clk),
    .RESET_B(net421),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[30] ),
    .Q_N(_14045_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[31]$_DFF_P_  (.CLK(clknet_leaf_641_clk),
    .RESET_B(net422),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[31] ),
    .Q_N(_14046_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[3]$_DFF_P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net423),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[3] ),
    .Q_N(_14047_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[4]$_DFF_P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net424),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[4] ),
    .Q_N(_14048_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[5]$_DFF_P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net425),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[5] ),
    .Q_N(_14049_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[6]$_DFF_P_  (.CLK(clknet_8_28_0_clk),
    .RESET_B(net426),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[6] ),
    .Q_N(_14050_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[7]$_DFF_P_  (.CLK(clknet_8_30_0_clk),
    .RESET_B(net427),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[7] ),
    .Q_N(_14051_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[8]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net428),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[8] ),
    .Q_N(_14052_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.alu_out_q[9]$_DFF_P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net429),
    .D(\u_ac_controller_soc_inst.u_picorv32.alu_out[9] ),
    .Q_N(_13634_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.alu_out_q[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[0]$_SDFF_PN0_  (.CLK(clknet_leaf_529_clk),
    .RESET_B(net430),
    .D(_00530_),
    .Q_N(_00140_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[10]$_SDFF_PN0_  (.CLK(clknet_leaf_509_clk),
    .RESET_B(net431),
    .D(_00531_),
    .Q_N(_13633_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[11]$_SDFF_PN0_  (.CLK(clknet_8_211_0_clk),
    .RESET_B(net432),
    .D(_00532_),
    .Q_N(_13632_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[12]$_SDFF_PN0_  (.CLK(clknet_leaf_513_clk),
    .RESET_B(net433),
    .D(_00533_),
    .Q_N(_13631_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[13]$_SDFF_PN0_  (.CLK(clknet_leaf_505_clk),
    .RESET_B(net434),
    .D(_00534_),
    .Q_N(_13630_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[14]$_SDFF_PN0_  (.CLK(clknet_leaf_566_clk),
    .RESET_B(net435),
    .D(_00535_),
    .Q_N(_13629_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[15]$_SDFF_PN0_  (.CLK(clknet_leaf_506_clk),
    .RESET_B(net436),
    .D(_00536_),
    .Q_N(_13628_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[16]$_SDFF_PN0_  (.CLK(clknet_leaf_506_clk),
    .RESET_B(net437),
    .D(_00537_),
    .Q_N(_13627_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[17]$_SDFF_PN0_  (.CLK(clknet_leaf_493_clk),
    .RESET_B(net438),
    .D(_00538_),
    .Q_N(_13626_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[18]$_SDFF_PN0_  (.CLK(clknet_leaf_625_clk),
    .RESET_B(net439),
    .D(_00539_),
    .Q_N(_13625_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[19]$_SDFF_PN0_  (.CLK(clknet_leaf_624_clk),
    .RESET_B(net440),
    .D(_00540_),
    .Q_N(_13624_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[1]$_SDFF_PN0_  (.CLK(clknet_leaf_525_clk),
    .RESET_B(net441),
    .D(_00541_),
    .Q_N(_13623_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[20]$_SDFF_PN0_  (.CLK(clknet_leaf_624_clk),
    .RESET_B(net442),
    .D(_00542_),
    .Q_N(_13622_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[21]$_SDFF_PN0_  (.CLK(clknet_8_206_0_clk),
    .RESET_B(net443),
    .D(_00543_),
    .Q_N(_13621_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[22]$_SDFF_PN0_  (.CLK(clknet_leaf_621_clk),
    .RESET_B(net444),
    .D(_00544_),
    .Q_N(_13620_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[23]$_SDFF_PN0_  (.CLK(clknet_leaf_592_clk),
    .RESET_B(net445),
    .D(_00545_),
    .Q_N(_13619_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[24]$_SDFF_PN0_  (.CLK(clknet_leaf_591_clk),
    .RESET_B(net446),
    .D(_00546_),
    .Q_N(_13618_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[25]$_SDFF_PN0_  (.CLK(clknet_leaf_621_clk),
    .RESET_B(net447),
    .D(_00547_),
    .Q_N(_13617_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[26]$_SDFF_PN0_  (.CLK(clknet_leaf_593_clk),
    .RESET_B(net448),
    .D(_00548_),
    .Q_N(_13616_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[27]$_SDFF_PN0_  (.CLK(clknet_leaf_593_clk),
    .RESET_B(net449),
    .D(_00549_),
    .Q_N(_13615_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[28]$_SDFF_PN0_  (.CLK(clknet_leaf_624_clk),
    .RESET_B(net450),
    .D(_00550_),
    .Q_N(_13614_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[29]$_SDFF_PN0_  (.CLK(clknet_8_206_0_clk),
    .RESET_B(net451),
    .D(_00551_),
    .Q_N(_13613_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[2]$_SDFF_PN0_  (.CLK(clknet_leaf_528_clk),
    .RESET_B(net452),
    .D(_00552_),
    .Q_N(_13612_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[30]$_SDFF_PN0_  (.CLK(clknet_leaf_495_clk),
    .RESET_B(net453),
    .D(_00553_),
    .Q_N(_13611_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[31]$_SDFF_PN0_  (.CLK(clknet_leaf_572_clk),
    .RESET_B(net454),
    .D(_00554_),
    .Q_N(_13610_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[32]$_SDFF_PN0_  (.CLK(clknet_leaf_507_clk),
    .RESET_B(net455),
    .D(_00555_),
    .Q_N(_13609_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[32] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[33]$_SDFF_PN0_  (.CLK(clknet_leaf_507_clk),
    .RESET_B(net456),
    .D(_00556_),
    .Q_N(_13608_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[33] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[34]$_SDFF_PN0_  (.CLK(clknet_leaf_533_clk),
    .RESET_B(net457),
    .D(_00557_),
    .Q_N(_13607_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[34] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[35]$_SDFF_PN0_  (.CLK(clknet_leaf_532_clk),
    .RESET_B(net458),
    .D(_00558_),
    .Q_N(_13606_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[35] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[36]$_SDFF_PN0_  (.CLK(clknet_leaf_532_clk),
    .RESET_B(net459),
    .D(_00559_),
    .Q_N(_13605_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[36] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[37]$_SDFF_PN0_  (.CLK(clknet_leaf_538_clk),
    .RESET_B(net460),
    .D(_00560_),
    .Q_N(_13604_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[37] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[38]$_SDFF_PN0_  (.CLK(clknet_leaf_535_clk),
    .RESET_B(net461),
    .D(_00561_),
    .Q_N(_13603_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[38] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[39]$_SDFF_PN0_  (.CLK(clknet_leaf_534_clk),
    .RESET_B(net462),
    .D(_00562_),
    .Q_N(_13602_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[39] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[3]$_SDFF_PN0_  (.CLK(clknet_leaf_528_clk),
    .RESET_B(net463),
    .D(_00563_),
    .Q_N(_13601_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[40]$_SDFF_PN0_  (.CLK(clknet_leaf_534_clk),
    .RESET_B(net464),
    .D(_00564_),
    .Q_N(_13600_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[40] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[41]$_SDFF_PN0_  (.CLK(clknet_8_214_0_clk),
    .RESET_B(net465),
    .D(_00565_),
    .Q_N(_13599_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[41] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[42]$_SDFF_PN0_  (.CLK(clknet_leaf_509_clk),
    .RESET_B(net466),
    .D(_00566_),
    .Q_N(_13598_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[42] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[43]$_SDFF_PN0_  (.CLK(clknet_leaf_508_clk),
    .RESET_B(net467),
    .D(_00567_),
    .Q_N(_13597_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[43] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[44]$_SDFF_PN0_  (.CLK(clknet_leaf_564_clk),
    .RESET_B(net468),
    .D(_00568_),
    .Q_N(_13596_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[44] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[45]$_SDFF_PN0_  (.CLK(clknet_leaf_565_clk),
    .RESET_B(net469),
    .D(_00569_),
    .Q_N(_13595_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[45] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[46]$_SDFF_PN0_  (.CLK(clknet_leaf_498_clk),
    .RESET_B(net470),
    .D(_00570_),
    .Q_N(_13594_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[46] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[47]$_SDFF_PN0_  (.CLK(clknet_leaf_571_clk),
    .RESET_B(net471),
    .D(_00571_),
    .Q_N(_13593_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[47] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[48]$_SDFF_PN0_  (.CLK(clknet_leaf_572_clk),
    .RESET_B(net472),
    .D(_00572_),
    .Q_N(_13592_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[48] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[49]$_SDFF_PN0_  (.CLK(clknet_leaf_495_clk),
    .RESET_B(net473),
    .D(_00573_),
    .Q_N(_13591_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[49] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[4]$_SDFF_PN0_  (.CLK(clknet_leaf_526_clk),
    .RESET_B(net474),
    .D(_00574_),
    .Q_N(_13590_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[50]$_SDFF_PN0_  (.CLK(clknet_leaf_574_clk),
    .RESET_B(net475),
    .D(_00575_),
    .Q_N(_13589_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[50] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[51]$_SDFF_PN0_  (.CLK(clknet_leaf_574_clk),
    .RESET_B(net476),
    .D(_00576_),
    .Q_N(_13588_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[51] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[52]$_SDFF_PN0_  (.CLK(clknet_8_206_0_clk),
    .RESET_B(net477),
    .D(_00577_),
    .Q_N(_13587_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[52] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[53]$_SDFF_PN0_  (.CLK(clknet_leaf_574_clk),
    .RESET_B(net478),
    .D(_00578_),
    .Q_N(_13586_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[53] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[54]$_SDFF_PN0_  (.CLK(clknet_leaf_586_clk),
    .RESET_B(net479),
    .D(_00579_),
    .Q_N(_13585_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[54] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[55]$_SDFF_PN0_  (.CLK(clknet_leaf_586_clk),
    .RESET_B(net480),
    .D(_00580_),
    .Q_N(_13584_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[55] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[56]$_SDFF_PN0_  (.CLK(clknet_leaf_592_clk),
    .RESET_B(net481),
    .D(_00581_),
    .Q_N(_13583_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[56] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[57]$_SDFF_PN0_  (.CLK(clknet_8_203_0_clk),
    .RESET_B(net482),
    .D(_00582_),
    .Q_N(_13582_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[57] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[58]$_SDFF_PN0_  (.CLK(clknet_leaf_586_clk),
    .RESET_B(net483),
    .D(_00583_),
    .Q_N(_13581_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[58] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[59]$_SDFF_PN0_  (.CLK(clknet_8_218_0_clk),
    .RESET_B(net484),
    .D(_00584_),
    .Q_N(_13580_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[59] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[5]$_SDFF_PN0_  (.CLK(clknet_8_209_0_clk),
    .RESET_B(net485),
    .D(_00585_),
    .Q_N(_13579_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[60]$_SDFF_PN0_  (.CLK(clknet_leaf_587_clk),
    .RESET_B(net486),
    .D(_00586_),
    .Q_N(_13578_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[60] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[61]$_SDFF_PN0_  (.CLK(clknet_leaf_578_clk),
    .RESET_B(net487),
    .D(_00587_),
    .Q_N(_13577_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[61] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[62]$_SDFF_PN0_  (.CLK(clknet_leaf_570_clk),
    .RESET_B(net488),
    .D(_00588_),
    .Q_N(_13576_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[62] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[63]$_SDFF_PN0_  (.CLK(clknet_leaf_572_clk),
    .RESET_B(net489),
    .D(_00589_),
    .Q_N(_13575_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[63] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[6]$_SDFF_PN0_  (.CLK(clknet_leaf_533_clk),
    .RESET_B(net490),
    .D(_00590_),
    .Q_N(_13574_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[7]$_SDFF_PN0_  (.CLK(clknet_leaf_533_clk),
    .RESET_B(net491),
    .D(_00591_),
    .Q_N(_13573_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[8]$_SDFF_PN0_  (.CLK(clknet_leaf_511_clk),
    .RESET_B(net492),
    .D(_00592_),
    .Q_N(_13572_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_cycle[9]$_SDFF_PN0_  (.CLK(clknet_leaf_511_clk),
    .RESET_B(net493),
    .D(_00593_),
    .Q_N(_13571_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_cycle[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_627_clk),
    .RESET_B(net494),
    .D(_00594_),
    .Q_N(_00141_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_556_clk),
    .RESET_B(net495),
    .D(_00595_),
    .Q_N(_13570_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[11]$_SDFFE_PN0P_  (.CLK(clknet_8_220_0_clk),
    .RESET_B(net496),
    .D(_00596_),
    .Q_N(_13569_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[12]$_SDFFE_PN0P_  (.CLK(clknet_8_221_0_clk),
    .RESET_B(net497),
    .D(_00597_),
    .Q_N(_13568_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_556_clk),
    .RESET_B(net498),
    .D(_00598_),
    .Q_N(_13567_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_558_clk),
    .RESET_B(net499),
    .D(_00599_),
    .Q_N(_13566_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_558_clk),
    .RESET_B(net500),
    .D(_00600_),
    .Q_N(_13565_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_557_clk),
    .RESET_B(net501),
    .D(_00601_),
    .Q_N(_13564_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_569_clk),
    .RESET_B(net502),
    .D(_00602_),
    .Q_N(_13563_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_557_clk),
    .RESET_B(net503),
    .D(_00603_),
    .Q_N(_13562_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_584_clk),
    .RESET_B(net504),
    .D(_00604_),
    .Q_N(_13561_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_625_clk),
    .RESET_B(net505),
    .D(_00605_),
    .Q_N(_13560_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_584_clk),
    .RESET_B(net506),
    .D(_00606_),
    .Q_N(_13559_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_583_clk),
    .RESET_B(net507),
    .D(_00607_),
    .Q_N(_13558_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_583_clk),
    .RESET_B(net508),
    .D(_00608_),
    .Q_N(_13557_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_582_clk),
    .RESET_B(net509),
    .D(_00609_),
    .Q_N(_13556_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_582_clk),
    .RESET_B(net510),
    .D(_00610_),
    .Q_N(_13555_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[25]$_SDFFE_PN0P_  (.CLK(clknet_8_219_0_clk),
    .RESET_B(net511),
    .D(_00611_),
    .Q_N(_13554_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[26]$_SDFFE_PN0P_  (.CLK(clknet_8_219_0_clk),
    .RESET_B(net512),
    .D(_00612_),
    .Q_N(_13553_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_578_clk),
    .RESET_B(net513),
    .D(_00613_),
    .Q_N(_13552_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_578_clk),
    .RESET_B(net514),
    .D(_00614_),
    .Q_N(_13551_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_579_clk),
    .RESET_B(net515),
    .D(_00615_),
    .Q_N(_13550_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_566_clk),
    .RESET_B(net516),
    .D(_00616_),
    .Q_N(_13549_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_569_clk),
    .RESET_B(net517),
    .D(_00617_),
    .Q_N(_13548_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_570_clk),
    .RESET_B(net518),
    .D(_00618_),
    .Q_N(_13547_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_570_clk),
    .RESET_B(net519),
    .D(_00619_),
    .Q_N(_13546_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[32] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_571_clk),
    .RESET_B(net520),
    .D(_00620_),
    .Q_N(_13545_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[33] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_567_clk),
    .RESET_B(net521),
    .D(_00621_),
    .Q_N(_13544_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[34] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_567_clk),
    .RESET_B(net522),
    .D(_00622_),
    .Q_N(_13543_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[35] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_564_clk),
    .RESET_B(net523),
    .D(_00623_),
    .Q_N(_13542_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[36] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_564_clk),
    .RESET_B(net524),
    .D(_00624_),
    .Q_N(_13541_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[37] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_555_clk),
    .RESET_B(net525),
    .D(_00625_),
    .Q_N(_13540_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[38] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_537_clk),
    .RESET_B(net526),
    .D(_00626_),
    .Q_N(_13539_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[39] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[3]$_SDFFE_PN0P_  (.CLK(clknet_8_222_0_clk),
    .RESET_B(net527),
    .D(_00627_),
    .Q_N(_13538_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_554_clk),
    .RESET_B(net528),
    .D(_00628_),
    .Q_N(_13537_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[40] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_554_clk),
    .RESET_B(net529),
    .D(_00629_),
    .Q_N(_13536_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[41] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_555_clk),
    .RESET_B(net530),
    .D(_00630_),
    .Q_N(_13535_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[42] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[43]$_SDFFE_PN0P_  (.CLK(clknet_8_220_0_clk),
    .RESET_B(net531),
    .D(_00631_),
    .Q_N(_13534_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[43] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[44]$_SDFFE_PN0P_  (.CLK(clknet_8_221_0_clk),
    .RESET_B(net532),
    .D(_00632_),
    .Q_N(_13533_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[44] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_559_clk),
    .RESET_B(net533),
    .D(_00633_),
    .Q_N(_13532_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[45] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_559_clk),
    .RESET_B(net534),
    .D(_00634_),
    .Q_N(_13531_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[46] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_559_clk),
    .RESET_B(net535),
    .D(_00635_),
    .Q_N(_13530_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[47] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_569_clk),
    .RESET_B(net536),
    .D(_00636_),
    .Q_N(_13529_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[48] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_581_clk),
    .RESET_B(net537),
    .D(_00637_),
    .Q_N(_13528_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[49] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_565_clk),
    .RESET_B(net538),
    .D(_00638_),
    .Q_N(_13527_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_581_clk),
    .RESET_B(net539),
    .D(_00639_),
    .Q_N(_13526_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[50] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_580_clk),
    .RESET_B(net540),
    .D(_00640_),
    .Q_N(_13525_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[51] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_580_clk),
    .RESET_B(net541),
    .D(_00641_),
    .Q_N(_13524_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[52] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_579_clk),
    .RESET_B(net542),
    .D(_00642_),
    .Q_N(_13523_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[53] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_582_clk),
    .RESET_B(net543),
    .D(_00643_),
    .Q_N(_13522_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[54] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_582_clk),
    .RESET_B(net544),
    .D(_00644_),
    .Q_N(_13521_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[55] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_585_clk),
    .RESET_B(net545),
    .D(_00645_),
    .Q_N(_13520_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[56] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_585_clk),
    .RESET_B(net546),
    .D(_00646_),
    .Q_N(_13519_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[57] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[58]$_SDFFE_PN0P_  (.CLK(clknet_8_218_0_clk),
    .RESET_B(net547),
    .D(_00647_),
    .Q_N(_13518_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[58] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_587_clk),
    .RESET_B(net548),
    .D(_00648_),
    .Q_N(_13517_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[59] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_555_clk),
    .RESET_B(net549),
    .D(_00649_),
    .Q_N(_13516_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_591_clk),
    .RESET_B(net550),
    .D(_00650_),
    .Q_N(_13515_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[60] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_591_clk),
    .RESET_B(net551),
    .D(_00651_),
    .Q_N(_13514_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[61] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_590_clk),
    .RESET_B(net552),
    .D(_00652_),
    .Q_N(_13513_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[62] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_590_clk),
    .RESET_B(net553),
    .D(_00653_),
    .Q_N(_13512_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[63] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_508_clk),
    .RESET_B(net554),
    .D(_00654_),
    .Q_N(_13511_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_535_clk),
    .RESET_B(net555),
    .D(_00655_),
    .Q_N(_13510_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_538_clk),
    .RESET_B(net556),
    .D(_00656_),
    .Q_N(_13509_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.count_instr[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_537_clk),
    .RESET_B(net557),
    .D(_00657_),
    .Q_N(_14053_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.count_instr[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpu_state[0]$_DFF_P_  (.CLK(clknet_leaf_477_clk),
    .RESET_B(net558),
    .D(_00010_),
    .Q_N(_14054_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpu_state[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpu_state[1]$_DFF_P_  (.CLK(clknet_leaf_486_clk),
    .RESET_B(net559),
    .D(_00011_),
    .Q_N(_14055_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpu_state[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpu_state[2]$_DFF_P_  (.CLK(clknet_leaf_465_clk),
    .RESET_B(net560),
    .D(_00012_),
    .Q_N(_14056_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpu_state[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpu_state[3]$_DFF_P_  (.CLK(clknet_8_196_0_clk),
    .RESET_B(net561),
    .D(_00013_),
    .Q_N(_00110_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpu_state[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpu_state[4]$_DFF_P_  (.CLK(clknet_leaf_466_clk),
    .RESET_B(net562),
    .D(_00014_),
    .Q_N(_00109_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpu_state[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpu_state[5]$_DFF_P_  (.CLK(clknet_leaf_472_clk),
    .RESET_B(net563),
    .D(_00015_),
    .Q_N(_00089_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpu_state[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpu_state[6]$_DFF_P_  (.CLK(clknet_leaf_472_clk),
    .RESET_B(net564),
    .D(_00016_),
    .Q_N(_00088_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpu_state[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][0]$_DFFE_PP_  (.CLK(clknet_8_145_0_clk),
    .RESET_B(net565),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][0] ),
    .Q_N(_13508_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_1077_clk),
    .RESET_B(net566),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][10] ),
    .Q_N(_13507_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_831_clk),
    .RESET_B(net567),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][11] ),
    .Q_N(_13506_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][12]$_DFFE_PP_  (.CLK(clknet_8_10_0_clk),
    .RESET_B(net568),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][12] ),
    .Q_N(_13505_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_1020_clk),
    .RESET_B(net569),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][13] ),
    .Q_N(_13504_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_937_clk),
    .RESET_B(net570),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][14] ),
    .Q_N(_13503_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_1147_clk),
    .RESET_B(net571),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][15] ),
    .Q_N(_13502_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_1114_clk),
    .RESET_B(net572),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][16] ),
    .Q_N(_13501_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][17]$_DFFE_PP_  (.CLK(clknet_8_45_0_clk),
    .RESET_B(net573),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][17] ),
    .Q_N(_13500_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_1052_clk),
    .RESET_B(net574),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][18] ),
    .Q_N(_13499_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_707_clk),
    .RESET_B(net575),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][19] ),
    .Q_N(_13498_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net576),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][1] ),
    .Q_N(_13497_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_1067_clk),
    .RESET_B(net577),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][20] ),
    .Q_N(_13496_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][21]$_DFFE_PP_  (.CLK(clknet_8_135_0_clk),
    .RESET_B(net578),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][21] ),
    .Q_N(_13495_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_821_clk),
    .RESET_B(net579),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][22] ),
    .Q_N(_13494_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_845_clk),
    .RESET_B(net580),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][23] ),
    .Q_N(_13493_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][24]$_DFFE_PP_  (.CLK(clknet_8_171_0_clk),
    .RESET_B(net581),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][24] ),
    .Q_N(_13492_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_816_clk),
    .RESET_B(net582),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][25] ),
    .Q_N(_13491_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_725_clk),
    .RESET_B(net583),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][26] ),
    .Q_N(_13490_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][27]$_DFFE_PP_  (.CLK(clknet_8_187_0_clk),
    .RESET_B(net584),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][27] ),
    .Q_N(_13489_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_712_clk),
    .RESET_B(net585),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][28] ),
    .Q_N(_13488_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_817_clk),
    .RESET_B(net586),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][29] ),
    .Q_N(_13487_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][2]$_DFFE_PP_  (.CLK(clknet_8_37_0_clk),
    .RESET_B(net587),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][2] ),
    .Q_N(_13486_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_688_clk),
    .RESET_B(net588),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][30] ),
    .Q_N(_13485_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_701_clk),
    .RESET_B(net589),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][31] ),
    .Q_N(_13484_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_1086_clk),
    .RESET_B(net590),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][3] ),
    .Q_N(_13483_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_1072_clk),
    .RESET_B(net591),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][4] ),
    .Q_N(_13482_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_1093_clk),
    .RESET_B(net592),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][5] ),
    .Q_N(_13481_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net593),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][6] ),
    .Q_N(_13480_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_1150_clk),
    .RESET_B(net594),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][7] ),
    .Q_N(_13479_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][8]$_DFFE_PP_  (.CLK(clknet_8_165_0_clk),
    .RESET_B(net595),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][8] ),
    .Q_N(_13478_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net596),
    .D(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][9] ),
    .Q_N(_13477_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[0][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_998_clk),
    .RESET_B(net597),
    .D(_00690_),
    .Q_N(_13476_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_1116_clk),
    .RESET_B(net598),
    .D(_00691_),
    .Q_N(_13475_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_781_clk),
    .RESET_B(net599),
    .D(_00692_),
    .Q_N(_13474_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][12]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net600),
    .D(_00693_),
    .Q_N(_13473_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][13]$_DFFE_PP_  (.CLK(clknet_leaf_1007_clk),
    .RESET_B(net601),
    .D(_00694_),
    .Q_N(_13472_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][14]$_DFFE_PP_  (.CLK(clknet_leaf_946_clk),
    .RESET_B(net602),
    .D(_00695_),
    .Q_N(_13471_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][15]$_DFFE_PP_  (.CLK(clknet_leaf_1105_clk),
    .RESET_B(net603),
    .D(_00696_),
    .Q_N(_13470_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][16]$_DFFE_PP_  (.CLK(clknet_leaf_1124_clk),
    .RESET_B(net604),
    .D(_00697_),
    .Q_N(_13469_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][17]$_DFFE_PP_  (.CLK(clknet_leaf_1127_clk),
    .RESET_B(net605),
    .D(_00698_),
    .Q_N(_13468_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][18]$_DFFE_PP_  (.CLK(clknet_leaf_924_clk),
    .RESET_B(net606),
    .D(_00699_),
    .Q_N(_13467_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][19]$_DFFE_PP_  (.CLK(clknet_leaf_743_clk),
    .RESET_B(net607),
    .D(_00700_),
    .Q_N(_13466_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net608),
    .D(_00701_),
    .Q_N(_13465_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][20]$_DFFE_PP_  (.CLK(clknet_leaf_888_clk),
    .RESET_B(net609),
    .D(_00702_),
    .Q_N(_13464_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][21]$_DFFE_PP_  (.CLK(clknet_leaf_890_clk),
    .RESET_B(net610),
    .D(_00703_),
    .Q_N(_13463_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][22]$_DFFE_PP_  (.CLK(clknet_leaf_852_clk),
    .RESET_B(net611),
    .D(_00704_),
    .Q_N(_13462_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][23]$_DFFE_PP_  (.CLK(clknet_leaf_905_clk),
    .RESET_B(net612),
    .D(_00705_),
    .Q_N(_13461_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][24]$_DFFE_PP_  (.CLK(clknet_leaf_851_clk),
    .RESET_B(net613),
    .D(_00706_),
    .Q_N(_13460_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][25]$_DFFE_PP_  (.CLK(clknet_leaf_773_clk),
    .RESET_B(net614),
    .D(_00707_),
    .Q_N(_13459_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][26]$_DFFE_PP_  (.CLK(clknet_8_232_0_clk),
    .RESET_B(net615),
    .D(_00708_),
    .Q_N(_13458_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][27]$_DFFE_PP_  (.CLK(clknet_leaf_754_clk),
    .RESET_B(net616),
    .D(_00709_),
    .Q_N(_13457_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][28]$_DFFE_PP_  (.CLK(clknet_leaf_739_clk),
    .RESET_B(net617),
    .D(_00710_),
    .Q_N(_13456_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][29]$_DFFE_PP_  (.CLK(clknet_leaf_775_clk),
    .RESET_B(net618),
    .D(_00711_),
    .Q_N(_13455_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][2]$_DFFE_PP_  (.CLK(clknet_8_56_0_clk),
    .RESET_B(net619),
    .D(_00712_),
    .Q_N(_13454_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][30]$_DFFE_PP_  (.CLK(clknet_leaf_685_clk),
    .RESET_B(net620),
    .D(_00713_),
    .Q_N(_13453_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][31]$_DFFE_PP_  (.CLK(clknet_8_172_0_clk),
    .RESET_B(net621),
    .D(_00714_),
    .Q_N(_13452_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_1106_clk),
    .RESET_B(net622),
    .D(_00715_),
    .Q_N(_13451_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_1071_clk),
    .RESET_B(net623),
    .D(_00716_),
    .Q_N(_13450_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net624),
    .D(_00717_),
    .Q_N(_13449_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net625),
    .D(_00718_),
    .Q_N(_13448_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net626),
    .D(_00719_),
    .Q_N(_13447_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_961_clk),
    .RESET_B(net627),
    .D(_00720_),
    .Q_N(_13446_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net628),
    .D(_00721_),
    .Q_N(_13445_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[10][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_1000_clk),
    .RESET_B(net629),
    .D(_00722_),
    .Q_N(_13444_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][10]$_DFFE_PP_  (.CLK(clknet_8_38_0_clk),
    .RESET_B(net630),
    .D(_00723_),
    .Q_N(_13443_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_778_clk),
    .RESET_B(net631),
    .D(_00724_),
    .Q_N(_13442_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][12]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net632),
    .D(_00725_),
    .Q_N(_13441_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][13]$_DFFE_PP_  (.CLK(clknet_leaf_1007_clk),
    .RESET_B(net633),
    .D(_00726_),
    .Q_N(_13440_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][14]$_DFFE_PP_  (.CLK(clknet_leaf_946_clk),
    .RESET_B(net634),
    .D(_00727_),
    .Q_N(_13439_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][15]$_DFFE_PP_  (.CLK(clknet_leaf_1104_clk),
    .RESET_B(net635),
    .D(_00728_),
    .Q_N(_13438_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][16]$_DFFE_PP_  (.CLK(clknet_leaf_1114_clk),
    .RESET_B(net636),
    .D(_00729_),
    .Q_N(_13437_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][17]$_DFFE_PP_  (.CLK(clknet_leaf_1128_clk),
    .RESET_B(net637),
    .D(_00730_),
    .Q_N(_13436_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][18]$_DFFE_PP_  (.CLK(clknet_8_154_0_clk),
    .RESET_B(net638),
    .D(_00731_),
    .Q_N(_13435_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][19]$_DFFE_PP_  (.CLK(clknet_leaf_744_clk),
    .RESET_B(net639),
    .D(_00732_),
    .Q_N(_13434_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net640),
    .D(_00733_),
    .Q_N(_13433_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][20]$_DFFE_PP_  (.CLK(clknet_8_136_0_clk),
    .RESET_B(net641),
    .D(_00734_),
    .Q_N(_13432_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][21]$_DFFE_PP_  (.CLK(clknet_leaf_888_clk),
    .RESET_B(net642),
    .D(_00735_),
    .Q_N(_13431_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][22]$_DFFE_PP_  (.CLK(clknet_leaf_852_clk),
    .RESET_B(net643),
    .D(_00736_),
    .Q_N(_13430_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][23]$_DFFE_PP_  (.CLK(clknet_leaf_877_clk),
    .RESET_B(net644),
    .D(_00737_),
    .Q_N(_13429_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][24]$_DFFE_PP_  (.CLK(clknet_leaf_853_clk),
    .RESET_B(net645),
    .D(_00738_),
    .Q_N(_13428_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][25]$_DFFE_PP_  (.CLK(clknet_8_182_0_clk),
    .RESET_B(net646),
    .D(_00739_),
    .Q_N(_13427_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][26]$_DFFE_PP_  (.CLK(clknet_leaf_738_clk),
    .RESET_B(net647),
    .D(_00740_),
    .Q_N(_13426_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][27]$_DFFE_PP_  (.CLK(clknet_leaf_757_clk),
    .RESET_B(net648),
    .D(_00741_),
    .Q_N(_13425_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][28]$_DFFE_PP_  (.CLK(clknet_8_238_0_clk),
    .RESET_B(net649),
    .D(_00742_),
    .Q_N(_13424_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][29]$_DFFE_PP_  (.CLK(clknet_leaf_774_clk),
    .RESET_B(net650),
    .D(_00743_),
    .Q_N(_13423_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_1131_clk),
    .RESET_B(net651),
    .D(_00744_),
    .Q_N(_13422_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][30]$_DFFE_PP_  (.CLK(clknet_8_180_0_clk),
    .RESET_B(net652),
    .D(_00745_),
    .Q_N(_13421_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][31]$_DFFE_PP_  (.CLK(clknet_leaf_838_clk),
    .RESET_B(net653),
    .D(_00746_),
    .Q_N(_13420_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_1101_clk),
    .RESET_B(net654),
    .D(_00747_),
    .Q_N(_13419_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_892_clk),
    .RESET_B(net655),
    .D(_00748_),
    .Q_N(_13418_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net656),
    .D(_00749_),
    .Q_N(_13417_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net657),
    .D(_00750_),
    .Q_N(_13416_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net658),
    .D(_00751_),
    .Q_N(_13415_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_961_clk),
    .RESET_B(net659),
    .D(_00752_),
    .Q_N(_13414_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net660),
    .D(_00753_),
    .Q_N(_13413_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[11][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_1005_clk),
    .RESET_B(net661),
    .D(_00754_),
    .Q_N(_13412_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_1113_clk),
    .RESET_B(net662),
    .D(_00755_),
    .Q_N(_13411_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_776_clk),
    .RESET_B(net663),
    .D(_00756_),
    .Q_N(_13410_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][12]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net664),
    .D(_00757_),
    .Q_N(_13409_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][13]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net665),
    .D(_00758_),
    .Q_N(_13408_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][14]$_DFFE_PP_  (.CLK(clknet_leaf_952_clk),
    .RESET_B(net666),
    .D(_00759_),
    .Q_N(_13407_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][15]$_DFFE_PP_  (.CLK(clknet_leaf_1105_clk),
    .RESET_B(net667),
    .D(_00760_),
    .Q_N(_13406_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][16]$_DFFE_PP_  (.CLK(clknet_leaf_1031_clk),
    .RESET_B(net668),
    .D(_00761_),
    .Q_N(_13405_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][17]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net669),
    .D(_00762_),
    .Q_N(_13404_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][18]$_DFFE_PP_  (.CLK(clknet_8_153_0_clk),
    .RESET_B(net670),
    .D(_00763_),
    .Q_N(_13403_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][19]$_DFFE_PP_  (.CLK(clknet_leaf_742_clk),
    .RESET_B(net671),
    .D(_00764_),
    .Q_N(_13402_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net672),
    .D(_00765_),
    .Q_N(_13401_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][20]$_DFFE_PP_  (.CLK(clknet_8_136_0_clk),
    .RESET_B(net673),
    .D(_00766_),
    .Q_N(_13400_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][21]$_DFFE_PP_  (.CLK(clknet_leaf_898_clk),
    .RESET_B(net674),
    .D(_00767_),
    .Q_N(_13399_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][22]$_DFFE_PP_  (.CLK(clknet_leaf_870_clk),
    .RESET_B(net675),
    .D(_00768_),
    .Q_N(_13398_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][23]$_DFFE_PP_  (.CLK(clknet_leaf_884_clk),
    .RESET_B(net676),
    .D(_00769_),
    .Q_N(_13397_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][24]$_DFFE_PP_  (.CLK(clknet_leaf_868_clk),
    .RESET_B(net677),
    .D(_00770_),
    .Q_N(_13396_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][25]$_DFFE_PP_  (.CLK(clknet_leaf_759_clk),
    .RESET_B(net678),
    .D(_00771_),
    .Q_N(_13395_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][26]$_DFFE_PP_  (.CLK(clknet_leaf_721_clk),
    .RESET_B(net679),
    .D(_00772_),
    .Q_N(_13394_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][27]$_DFFE_PP_  (.CLK(clknet_8_189_0_clk),
    .RESET_B(net680),
    .D(_00773_),
    .Q_N(_13393_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][28]$_DFFE_PP_  (.CLK(clknet_leaf_721_clk),
    .RESET_B(net681),
    .D(_00774_),
    .Q_N(_13392_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][29]$_DFFE_PP_  (.CLK(clknet_leaf_774_clk),
    .RESET_B(net682),
    .D(_00775_),
    .Q_N(_13391_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][2]$_DFFE_PP_  (.CLK(clknet_8_51_0_clk),
    .RESET_B(net683),
    .D(_00776_),
    .Q_N(_13390_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][30]$_DFFE_PP_  (.CLK(clknet_leaf_777_clk),
    .RESET_B(net684),
    .D(_00777_),
    .Q_N(_13389_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][31]$_DFFE_PP_  (.CLK(clknet_leaf_681_clk),
    .RESET_B(net685),
    .D(_00778_),
    .Q_N(_13388_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_1110_clk),
    .RESET_B(net686),
    .D(_00779_),
    .Q_N(_13387_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_891_clk),
    .RESET_B(net687),
    .D(_00780_),
    .Q_N(_13386_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net688),
    .D(_00781_),
    .Q_N(_13385_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net689),
    .D(_00782_),
    .Q_N(_13384_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net690),
    .D(_00783_),
    .Q_N(_13383_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_957_clk),
    .RESET_B(net691),
    .D(_00784_),
    .Q_N(_13382_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net692),
    .D(_00785_),
    .Q_N(_13381_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[12][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_1009_clk),
    .RESET_B(net693),
    .D(_00786_),
    .Q_N(_13380_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_1113_clk),
    .RESET_B(net694),
    .D(_00787_),
    .Q_N(_13379_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_781_clk),
    .RESET_B(net695),
    .D(_00788_),
    .Q_N(_13378_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][12]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net696),
    .D(_00789_),
    .Q_N(_13377_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][13]$_DFFE_PP_  (.CLK(clknet_leaf_1015_clk),
    .RESET_B(net697),
    .D(_00790_),
    .Q_N(_13376_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][14]$_DFFE_PP_  (.CLK(clknet_leaf_951_clk),
    .RESET_B(net698),
    .D(_00791_),
    .Q_N(_13375_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][15]$_DFFE_PP_  (.CLK(clknet_8_37_0_clk),
    .RESET_B(net699),
    .D(_00792_),
    .Q_N(_13374_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][16]$_DFFE_PP_  (.CLK(clknet_8_47_0_clk),
    .RESET_B(net700),
    .D(_00793_),
    .Q_N(_13373_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][17]$_DFFE_PP_  (.CLK(clknet_leaf_1127_clk),
    .RESET_B(net701),
    .D(_00794_),
    .Q_N(_13372_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][18]$_DFFE_PP_  (.CLK(clknet_leaf_963_clk),
    .RESET_B(net702),
    .D(_00795_),
    .Q_N(_13371_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][19]$_DFFE_PP_  (.CLK(clknet_leaf_742_clk),
    .RESET_B(net703),
    .D(_00796_),
    .Q_N(_13370_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net704),
    .D(_00797_),
    .Q_N(_13369_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][20]$_DFFE_PP_  (.CLK(clknet_leaf_888_clk),
    .RESET_B(net705),
    .D(_00798_),
    .Q_N(_13368_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][21]$_DFFE_PP_  (.CLK(clknet_8_140_0_clk),
    .RESET_B(net706),
    .D(_00799_),
    .Q_N(_13367_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][22]$_DFFE_PP_  (.CLK(clknet_leaf_869_clk),
    .RESET_B(net707),
    .D(_00800_),
    .Q_N(_13366_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][23]$_DFFE_PP_  (.CLK(clknet_leaf_883_clk),
    .RESET_B(net708),
    .D(_00801_),
    .Q_N(_13365_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][24]$_DFFE_PP_  (.CLK(clknet_leaf_868_clk),
    .RESET_B(net709),
    .D(_00802_),
    .Q_N(_13364_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][25]$_DFFE_PP_  (.CLK(clknet_leaf_797_clk),
    .RESET_B(net710),
    .D(_00803_),
    .Q_N(_13363_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][26]$_DFFE_PP_  (.CLK(clknet_leaf_727_clk),
    .RESET_B(net711),
    .D(_00804_),
    .Q_N(_13362_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][27]$_DFFE_PP_  (.CLK(clknet_8_189_0_clk),
    .RESET_B(net712),
    .D(_00805_),
    .Q_N(_13361_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][28]$_DFFE_PP_  (.CLK(clknet_leaf_726_clk),
    .RESET_B(net713),
    .D(_00806_),
    .Q_N(_13360_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][29]$_DFFE_PP_  (.CLK(clknet_leaf_786_clk),
    .RESET_B(net714),
    .D(_00807_),
    .Q_N(_13359_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net715),
    .D(_00808_),
    .Q_N(_13358_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][30]$_DFFE_PP_  (.CLK(clknet_leaf_685_clk),
    .RESET_B(net716),
    .D(_00809_),
    .Q_N(_13357_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][31]$_DFFE_PP_  (.CLK(clknet_leaf_682_clk),
    .RESET_B(net717),
    .D(_00810_),
    .Q_N(_13356_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_1109_clk),
    .RESET_B(net718),
    .D(_00811_),
    .Q_N(_13355_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_891_clk),
    .RESET_B(net719),
    .D(_00812_),
    .Q_N(_13354_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net720),
    .D(_00813_),
    .Q_N(_13353_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net721),
    .D(_00814_),
    .Q_N(_13352_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net722),
    .D(_00815_),
    .Q_N(_13351_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_962_clk),
    .RESET_B(net723),
    .D(_00816_),
    .Q_N(_13350_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net724),
    .D(_00817_),
    .Q_N(_13349_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[13][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_1005_clk),
    .RESET_B(net725),
    .D(_00818_),
    .Q_N(_13348_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_1110_clk),
    .RESET_B(net726),
    .D(_00819_),
    .Q_N(_13347_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][11]$_DFFE_PP_  (.CLK(clknet_8_176_0_clk),
    .RESET_B(net727),
    .D(_00820_),
    .Q_N(_13346_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][12]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net728),
    .D(_00821_),
    .Q_N(_13345_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][13]$_DFFE_PP_  (.CLK(clknet_leaf_1015_clk),
    .RESET_B(net729),
    .D(_00822_),
    .Q_N(_13344_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][14]$_DFFE_PP_  (.CLK(clknet_leaf_951_clk),
    .RESET_B(net730),
    .D(_00823_),
    .Q_N(_13343_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][15]$_DFFE_PP_  (.CLK(clknet_8_39_0_clk),
    .RESET_B(net731),
    .D(_00824_),
    .Q_N(_13342_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][16]$_DFFE_PP_  (.CLK(clknet_leaf_1033_clk),
    .RESET_B(net732),
    .D(_00825_),
    .Q_N(_13341_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][17]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net733),
    .D(_00826_),
    .Q_N(_13340_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][18]$_DFFE_PP_  (.CLK(clknet_leaf_917_clk),
    .RESET_B(net734),
    .D(_00827_),
    .Q_N(_13339_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][19]$_DFFE_PP_  (.CLK(clknet_leaf_742_clk),
    .RESET_B(net735),
    .D(_00828_),
    .Q_N(_13338_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][1]$_DFFE_PP_  (.CLK(clknet_8_11_0_clk),
    .RESET_B(net736),
    .D(_00829_),
    .Q_N(_13337_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][20]$_DFFE_PP_  (.CLK(clknet_leaf_886_clk),
    .RESET_B(net737),
    .D(_00830_),
    .Q_N(_13336_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][21]$_DFFE_PP_  (.CLK(clknet_leaf_896_clk),
    .RESET_B(net738),
    .D(_00831_),
    .Q_N(_13335_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][22]$_DFFE_PP_  (.CLK(clknet_leaf_869_clk),
    .RESET_B(net739),
    .D(_00832_),
    .Q_N(_13334_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][23]$_DFFE_PP_  (.CLK(clknet_leaf_870_clk),
    .RESET_B(net740),
    .D(_00833_),
    .Q_N(_13333_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][24]$_DFFE_PP_  (.CLK(clknet_leaf_865_clk),
    .RESET_B(net741),
    .D(_00834_),
    .Q_N(_13332_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][25]$_DFFE_PP_  (.CLK(clknet_8_182_0_clk),
    .RESET_B(net742),
    .D(_00835_),
    .Q_N(_13331_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][26]$_DFFE_PP_  (.CLK(clknet_leaf_727_clk),
    .RESET_B(net743),
    .D(_00836_),
    .Q_N(_13330_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][27]$_DFFE_PP_  (.CLK(clknet_8_188_0_clk),
    .RESET_B(net744),
    .D(_00837_),
    .Q_N(_13329_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][28]$_DFFE_PP_  (.CLK(clknet_leaf_722_clk),
    .RESET_B(net745),
    .D(_00838_),
    .Q_N(_13328_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][29]$_DFFE_PP_  (.CLK(clknet_leaf_786_clk),
    .RESET_B(net746),
    .D(_00839_),
    .Q_N(_13327_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][2]$_DFFE_PP_  (.CLK(clknet_8_55_0_clk),
    .RESET_B(net747),
    .D(_00840_),
    .Q_N(_13326_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][30]$_DFFE_PP_  (.CLK(clknet_leaf_775_clk),
    .RESET_B(net748),
    .D(_00841_),
    .Q_N(_13325_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][31]$_DFFE_PP_  (.CLK(clknet_leaf_941_clk),
    .RESET_B(net749),
    .D(_00842_),
    .Q_N(_13324_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_1109_clk),
    .RESET_B(net750),
    .D(_00843_),
    .Q_N(_13323_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_1071_clk),
    .RESET_B(net751),
    .D(_00844_),
    .Q_N(_13322_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net752),
    .D(_00845_),
    .Q_N(_13321_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net753),
    .D(_00846_),
    .Q_N(_13320_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net754),
    .D(_00847_),
    .Q_N(_13319_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][8]$_DFFE_PP_  (.CLK(clknet_8_158_0_clk),
    .RESET_B(net755),
    .D(_00848_),
    .Q_N(_13318_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net756),
    .D(_00849_),
    .Q_N(_13317_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[14][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_1004_clk),
    .RESET_B(net757),
    .D(_00850_),
    .Q_N(_13316_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_1112_clk),
    .RESET_B(net758),
    .D(_00851_),
    .Q_N(_13315_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][11]$_DFFE_PP_  (.CLK(clknet_8_176_0_clk),
    .RESET_B(net759),
    .D(_00852_),
    .Q_N(_13314_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][12]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net760),
    .D(_00853_),
    .Q_N(_13313_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][13]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net761),
    .D(_00854_),
    .Q_N(_13312_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][14]$_DFFE_PP_  (.CLK(clknet_leaf_672_clk),
    .RESET_B(net762),
    .D(_00855_),
    .Q_N(_13311_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][15]$_DFFE_PP_  (.CLK(clknet_leaf_1120_clk),
    .RESET_B(net763),
    .D(_00856_),
    .Q_N(_13310_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][16]$_DFFE_PP_  (.CLK(clknet_leaf_1031_clk),
    .RESET_B(net764),
    .D(_00857_),
    .Q_N(_13309_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][17]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net765),
    .D(_00858_),
    .Q_N(_13308_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][18]$_DFFE_PP_  (.CLK(clknet_leaf_921_clk),
    .RESET_B(net766),
    .D(_00859_),
    .Q_N(_13307_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][19]$_DFFE_PP_  (.CLK(clknet_8_234_0_clk),
    .RESET_B(net767),
    .D(_00860_),
    .Q_N(_13306_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net768),
    .D(_00861_),
    .Q_N(_13305_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][20]$_DFFE_PP_  (.CLK(clknet_leaf_886_clk),
    .RESET_B(net769),
    .D(_00862_),
    .Q_N(_13304_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][21]$_DFFE_PP_  (.CLK(clknet_leaf_896_clk),
    .RESET_B(net770),
    .D(_00863_),
    .Q_N(_13303_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][22]$_DFFE_PP_  (.CLK(clknet_leaf_868_clk),
    .RESET_B(net771),
    .D(_00864_),
    .Q_N(_13302_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][23]$_DFFE_PP_  (.CLK(clknet_8_138_0_clk),
    .RESET_B(net772),
    .D(_00865_),
    .Q_N(_13301_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][24]$_DFFE_PP_  (.CLK(clknet_leaf_865_clk),
    .RESET_B(net773),
    .D(_00866_),
    .Q_N(_13300_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][25]$_DFFE_PP_  (.CLK(clknet_leaf_798_clk),
    .RESET_B(net774),
    .D(_00867_),
    .Q_N(_13299_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][26]$_DFFE_PP_  (.CLK(clknet_leaf_738_clk),
    .RESET_B(net775),
    .D(_00868_),
    .Q_N(_13298_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][27]$_DFFE_PP_  (.CLK(clknet_leaf_744_clk),
    .RESET_B(net776),
    .D(_00869_),
    .Q_N(_13297_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][28]$_DFFE_PP_  (.CLK(clknet_leaf_726_clk),
    .RESET_B(net777),
    .D(_00870_),
    .Q_N(_13296_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][29]$_DFFE_PP_  (.CLK(clknet_leaf_797_clk),
    .RESET_B(net778),
    .D(_00871_),
    .Q_N(_13295_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net779),
    .D(_00872_),
    .Q_N(_13294_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][30]$_DFFE_PP_  (.CLK(clknet_leaf_776_clk),
    .RESET_B(net780),
    .D(_00873_),
    .Q_N(_13293_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][31]$_DFFE_PP_  (.CLK(clknet_8_173_0_clk),
    .RESET_B(net781),
    .D(_00874_),
    .Q_N(_13292_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][3]$_DFFE_PP_  (.CLK(clknet_8_43_0_clk),
    .RESET_B(net782),
    .D(_00875_),
    .Q_N(_13291_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_890_clk),
    .RESET_B(net783),
    .D(_00876_),
    .Q_N(_13290_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net784),
    .D(_00877_),
    .Q_N(_13289_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net785),
    .D(_00878_),
    .Q_N(_13288_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net786),
    .D(_00879_),
    .Q_N(_13287_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_957_clk),
    .RESET_B(net787),
    .D(_00880_),
    .Q_N(_13286_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net788),
    .D(_00881_),
    .Q_N(_13285_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[15][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_1041_clk),
    .RESET_B(net789),
    .D(_00882_),
    .Q_N(_13284_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_1079_clk),
    .RESET_B(net790),
    .D(_00883_),
    .Q_N(_13283_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_840_clk),
    .RESET_B(net791),
    .D(_00884_),
    .Q_N(_13282_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net792),
    .D(_00885_),
    .Q_N(_13281_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][13]$_DFFE_PP_  (.CLK(clknet_leaf_1028_clk),
    .RESET_B(net793),
    .D(_00886_),
    .Q_N(_13280_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][14]$_DFFE_PP_  (.CLK(clknet_leaf_942_clk),
    .RESET_B(net794),
    .D(_00887_),
    .Q_N(_13279_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][15]$_DFFE_PP_  (.CLK(clknet_leaf_1097_clk),
    .RESET_B(net795),
    .D(_00888_),
    .Q_N(_13278_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][16]$_DFFE_PP_  (.CLK(clknet_leaf_1040_clk),
    .RESET_B(net796),
    .D(_00889_),
    .Q_N(_13277_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][17]$_DFFE_PP_  (.CLK(clknet_leaf_1023_clk),
    .RESET_B(net797),
    .D(_00890_),
    .Q_N(_13276_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][18]$_DFFE_PP_  (.CLK(clknet_leaf_926_clk),
    .RESET_B(net798),
    .D(_00891_),
    .Q_N(_13275_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][19]$_DFFE_PP_  (.CLK(clknet_leaf_695_clk),
    .RESET_B(net799),
    .D(_00892_),
    .Q_N(_13274_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net800),
    .D(_00893_),
    .Q_N(_13273_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][20]$_DFFE_PP_  (.CLK(clknet_leaf_903_clk),
    .RESET_B(net801),
    .D(_00894_),
    .Q_N(_13272_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][21]$_DFFE_PP_  (.CLK(clknet_leaf_907_clk),
    .RESET_B(net802),
    .D(_00895_),
    .Q_N(_13271_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][22]$_DFFE_PP_  (.CLK(clknet_leaf_861_clk),
    .RESET_B(net803),
    .D(_00896_),
    .Q_N(_13270_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][23]$_DFFE_PP_  (.CLK(clknet_leaf_842_clk),
    .RESET_B(net804),
    .D(_00897_),
    .Q_N(_13269_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][24]$_DFFE_PP_  (.CLK(clknet_leaf_860_clk),
    .RESET_B(net805),
    .D(_00898_),
    .Q_N(_13268_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][25]$_DFFE_PP_  (.CLK(clknet_leaf_798_clk),
    .RESET_B(net806),
    .D(_00899_),
    .Q_N(_13267_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][26]$_DFFE_PP_  (.CLK(clknet_leaf_769_clk),
    .RESET_B(net807),
    .D(_00900_),
    .Q_N(_13266_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][27]$_DFFE_PP_  (.CLK(clknet_leaf_755_clk),
    .RESET_B(net808),
    .D(_00901_),
    .Q_N(_13265_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][28]$_DFFE_PP_  (.CLK(clknet_leaf_718_clk),
    .RESET_B(net809),
    .D(_00902_),
    .Q_N(_13264_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][29]$_DFFE_PP_  (.CLK(clknet_leaf_800_clk),
    .RESET_B(net810),
    .D(_00903_),
    .Q_N(_13263_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_1142_clk),
    .RESET_B(net811),
    .D(_00904_),
    .Q_N(_13262_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][30]$_DFFE_PP_  (.CLK(clknet_leaf_692_clk),
    .RESET_B(net812),
    .D(_00905_),
    .Q_N(_13261_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][31]$_DFFE_PP_  (.CLK(clknet_leaf_696_clk),
    .RESET_B(net813),
    .D(_00906_),
    .Q_N(_13260_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_1085_clk),
    .RESET_B(net814),
    .D(_00907_),
    .Q_N(_13259_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_1075_clk),
    .RESET_B(net815),
    .D(_00908_),
    .Q_N(_13258_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_1097_clk),
    .RESET_B(net816),
    .D(_00909_),
    .Q_N(_13257_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][6]$_DFFE_PP_  (.CLK(clknet_8_2_0_clk),
    .RESET_B(net817),
    .D(_00910_),
    .Q_N(_13256_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net818),
    .D(_00911_),
    .Q_N(_13255_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_923_clk),
    .RESET_B(net819),
    .D(_00912_),
    .Q_N(_13254_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net820),
    .D(_00913_),
    .Q_N(_13253_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[16][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_1043_clk),
    .RESET_B(net821),
    .D(_00914_),
    .Q_N(_13252_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_1090_clk),
    .RESET_B(net822),
    .D(_00915_),
    .Q_N(_13251_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_838_clk),
    .RESET_B(net823),
    .D(_00916_),
    .Q_N(_13250_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net824),
    .D(_00917_),
    .Q_N(_13249_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][13]$_DFFE_PP_  (.CLK(clknet_leaf_1018_clk),
    .RESET_B(net825),
    .D(_00918_),
    .Q_N(_13248_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][14]$_DFFE_PP_  (.CLK(clknet_8_167_0_clk),
    .RESET_B(net826),
    .D(_00919_),
    .Q_N(_13247_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][15]$_DFFE_PP_  (.CLK(clknet_leaf_1098_clk),
    .RESET_B(net827),
    .D(_00920_),
    .Q_N(_13246_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][16]$_DFFE_PP_  (.CLK(clknet_leaf_1037_clk),
    .RESET_B(net828),
    .D(_00921_),
    .Q_N(_13245_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][17]$_DFFE_PP_  (.CLK(clknet_leaf_1022_clk),
    .RESET_B(net829),
    .D(_00922_),
    .Q_N(_13244_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][18]$_DFFE_PP_  (.CLK(clknet_leaf_926_clk),
    .RESET_B(net830),
    .D(_00923_),
    .Q_N(_13243_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][19]$_DFFE_PP_  (.CLK(clknet_leaf_717_clk),
    .RESET_B(net831),
    .D(_00924_),
    .Q_N(_13242_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net832),
    .D(_00925_),
    .Q_N(_13241_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][20]$_DFFE_PP_  (.CLK(clknet_leaf_903_clk),
    .RESET_B(net833),
    .D(_00926_),
    .Q_N(_13240_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][21]$_DFFE_PP_  (.CLK(clknet_leaf_929_clk),
    .RESET_B(net834),
    .D(_00927_),
    .Q_N(_13239_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][22]$_DFFE_PP_  (.CLK(clknet_leaf_860_clk),
    .RESET_B(net835),
    .D(_00928_),
    .Q_N(_13238_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][23]$_DFFE_PP_  (.CLK(clknet_leaf_841_clk),
    .RESET_B(net836),
    .D(_00929_),
    .Q_N(_13237_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][24]$_DFFE_PP_  (.CLK(clknet_leaf_859_clk),
    .RESET_B(net837),
    .D(_00930_),
    .Q_N(_13236_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][25]$_DFFE_PP_  (.CLK(clknet_8_177_0_clk),
    .RESET_B(net838),
    .D(_00931_),
    .Q_N(_13235_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][26]$_DFFE_PP_  (.CLK(clknet_leaf_770_clk),
    .RESET_B(net839),
    .D(_00932_),
    .Q_N(_13234_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][27]$_DFFE_PP_  (.CLK(clknet_leaf_799_clk),
    .RESET_B(net840),
    .D(_00933_),
    .Q_N(_13233_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][28]$_DFFE_PP_  (.CLK(clknet_leaf_717_clk),
    .RESET_B(net841),
    .D(_00934_),
    .Q_N(_13232_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][29]$_DFFE_PP_  (.CLK(clknet_leaf_800_clk),
    .RESET_B(net842),
    .D(_00935_),
    .Q_N(_13231_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_1142_clk),
    .RESET_B(net843),
    .D(_00936_),
    .Q_N(_13230_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][30]$_DFFE_PP_  (.CLK(clknet_leaf_693_clk),
    .RESET_B(net844),
    .D(_00937_),
    .Q_N(_13229_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][31]$_DFFE_PP_  (.CLK(clknet_leaf_695_clk),
    .RESET_B(net845),
    .D(_00938_),
    .Q_N(_13228_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_1084_clk),
    .RESET_B(net846),
    .D(_00939_),
    .Q_N(_13227_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][4]$_DFFE_PP_  (.CLK(clknet_8_129_0_clk),
    .RESET_B(net847),
    .D(_00940_),
    .Q_N(_13226_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_1148_clk),
    .RESET_B(net848),
    .D(_00941_),
    .Q_N(_13225_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net849),
    .D(_00942_),
    .Q_N(_13224_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net850),
    .D(_00943_),
    .Q_N(_13223_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][8]$_DFFE_PP_  (.CLK(clknet_8_154_0_clk),
    .RESET_B(net851),
    .D(_00944_),
    .Q_N(_13222_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net852),
    .D(_00945_),
    .Q_N(_13221_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[17][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_1004_clk),
    .RESET_B(net853),
    .D(_00946_),
    .Q_N(_13220_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_1078_clk),
    .RESET_B(net854),
    .D(_00947_),
    .Q_N(_13219_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_837_clk),
    .RESET_B(net855),
    .D(_00948_),
    .Q_N(_13218_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][12]$_DFFE_PP_  (.CLK(clknet_8_8_0_clk),
    .RESET_B(net856),
    .D(_00949_),
    .Q_N(_13217_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][13]$_DFFE_PP_  (.CLK(clknet_leaf_1005_clk),
    .RESET_B(net857),
    .D(_00950_),
    .Q_N(_13216_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][14]$_DFFE_PP_  (.CLK(clknet_leaf_941_clk),
    .RESET_B(net858),
    .D(_00951_),
    .Q_N(_13215_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][15]$_DFFE_PP_  (.CLK(clknet_leaf_1148_clk),
    .RESET_B(net859),
    .D(_00952_),
    .Q_N(_13214_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][16]$_DFFE_PP_  (.CLK(clknet_leaf_1034_clk),
    .RESET_B(net860),
    .D(_00953_),
    .Q_N(_13213_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][17]$_DFFE_PP_  (.CLK(clknet_leaf_1023_clk),
    .RESET_B(net861),
    .D(_00954_),
    .Q_N(_13212_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][18]$_DFFE_PP_  (.CLK(clknet_leaf_907_clk),
    .RESET_B(net862),
    .D(_00955_),
    .Q_N(_13211_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][19]$_DFFE_PP_  (.CLK(clknet_8_226_0_clk),
    .RESET_B(net863),
    .D(_00956_),
    .Q_N(_13210_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net864),
    .D(_00957_),
    .Q_N(_13209_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][20]$_DFFE_PP_  (.CLK(clknet_8_141_0_clk),
    .RESET_B(net865),
    .D(_00958_),
    .Q_N(_13208_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][21]$_DFFE_PP_  (.CLK(clknet_leaf_909_clk),
    .RESET_B(net866),
    .D(_00959_),
    .Q_N(_13207_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][22]$_DFFE_PP_  (.CLK(clknet_leaf_863_clk),
    .RESET_B(net867),
    .D(_00960_),
    .Q_N(_13206_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][23]$_DFFE_PP_  (.CLK(clknet_leaf_842_clk),
    .RESET_B(net868),
    .D(_00961_),
    .Q_N(_13205_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][24]$_DFFE_PP_  (.CLK(clknet_leaf_821_clk),
    .RESET_B(net869),
    .D(_00962_),
    .Q_N(_13204_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][25]$_DFFE_PP_  (.CLK(clknet_leaf_798_clk),
    .RESET_B(net870),
    .D(_00963_),
    .Q_N(_13203_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][26]$_DFFE_PP_  (.CLK(clknet_leaf_767_clk),
    .RESET_B(net871),
    .D(_00964_),
    .Q_N(_13202_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][27]$_DFFE_PP_  (.CLK(clknet_leaf_803_clk),
    .RESET_B(net872),
    .D(_00965_),
    .Q_N(_13201_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][28]$_DFFE_PP_  (.CLK(clknet_8_227_0_clk),
    .RESET_B(net873),
    .D(_00966_),
    .Q_N(_13200_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][29]$_DFFE_PP_  (.CLK(clknet_leaf_803_clk),
    .RESET_B(net874),
    .D(_00967_),
    .Q_N(_13199_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_1144_clk),
    .RESET_B(net875),
    .D(_00968_),
    .Q_N(_13198_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][30]$_DFFE_PP_  (.CLK(clknet_leaf_693_clk),
    .RESET_B(net876),
    .D(_00969_),
    .Q_N(_13197_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][31]$_DFFE_PP_  (.CLK(clknet_leaf_696_clk),
    .RESET_B(net877),
    .D(_00970_),
    .Q_N(_13196_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_1085_clk),
    .RESET_B(net878),
    .D(_00971_),
    .Q_N(_13195_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_1073_clk),
    .RESET_B(net879),
    .D(_00972_),
    .Q_N(_13194_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_1097_clk),
    .RESET_B(net880),
    .D(_00973_),
    .Q_N(_13193_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net881),
    .D(_00974_),
    .Q_N(_13192_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net882),
    .D(_00975_),
    .Q_N(_13191_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_920_clk),
    .RESET_B(net883),
    .D(_00976_),
    .Q_N(_13190_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net884),
    .D(_00977_),
    .Q_N(_13189_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[18][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_1046_clk),
    .RESET_B(net885),
    .D(_00978_),
    .Q_N(_13188_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_1078_clk),
    .RESET_B(net886),
    .D(_00979_),
    .Q_N(_13187_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_838_clk),
    .RESET_B(net887),
    .D(_00980_),
    .Q_N(_13186_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][12]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net888),
    .D(_00981_),
    .Q_N(_13185_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][13]$_DFFE_PP_  (.CLK(clknet_leaf_1041_clk),
    .RESET_B(net889),
    .D(_00982_),
    .Q_N(_13184_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][14]$_DFFE_PP_  (.CLK(clknet_leaf_840_clk),
    .RESET_B(net890),
    .D(_00983_),
    .Q_N(_13183_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][15]$_DFFE_PP_  (.CLK(clknet_leaf_1098_clk),
    .RESET_B(net891),
    .D(_00984_),
    .Q_N(_13182_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][16]$_DFFE_PP_  (.CLK(clknet_8_46_0_clk),
    .RESET_B(net892),
    .D(_00985_),
    .Q_N(_13181_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][17]$_DFFE_PP_  (.CLK(clknet_leaf_1022_clk),
    .RESET_B(net893),
    .D(_00986_),
    .Q_N(_13180_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][18]$_DFFE_PP_  (.CLK(clknet_leaf_934_clk),
    .RESET_B(net894),
    .D(_00987_),
    .Q_N(_13179_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][19]$_DFFE_PP_  (.CLK(clknet_leaf_694_clk),
    .RESET_B(net895),
    .D(_00988_),
    .Q_N(_13178_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][1]$_DFFE_PP_  (.CLK(clknet_8_58_0_clk),
    .RESET_B(net896),
    .D(_00989_),
    .Q_N(_13177_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][20]$_DFFE_PP_  (.CLK(clknet_leaf_905_clk),
    .RESET_B(net897),
    .D(_00990_),
    .Q_N(_13176_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][21]$_DFFE_PP_  (.CLK(clknet_leaf_927_clk),
    .RESET_B(net898),
    .D(_00991_),
    .Q_N(_13175_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][22]$_DFFE_PP_  (.CLK(clknet_8_168_0_clk),
    .RESET_B(net899),
    .D(_00992_),
    .Q_N(_13174_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][23]$_DFFE_PP_  (.CLK(clknet_leaf_841_clk),
    .RESET_B(net900),
    .D(_00993_),
    .Q_N(_13173_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][24]$_DFFE_PP_  (.CLK(clknet_8_170_0_clk),
    .RESET_B(net901),
    .D(_00994_),
    .Q_N(_13172_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][25]$_DFFE_PP_  (.CLK(clknet_leaf_800_clk),
    .RESET_B(net902),
    .D(_00995_),
    .Q_N(_13171_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][26]$_DFFE_PP_  (.CLK(clknet_leaf_767_clk),
    .RESET_B(net903),
    .D(_00996_),
    .Q_N(_13170_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][27]$_DFFE_PP_  (.CLK(clknet_leaf_755_clk),
    .RESET_B(net904),
    .D(_00997_),
    .Q_N(_13169_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][28]$_DFFE_PP_  (.CLK(clknet_leaf_718_clk),
    .RESET_B(net905),
    .D(_00998_),
    .Q_N(_13168_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][29]$_DFFE_PP_  (.CLK(clknet_leaf_801_clk),
    .RESET_B(net906),
    .D(_00999_),
    .Q_N(_13167_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_1142_clk),
    .RESET_B(net907),
    .D(_01000_),
    .Q_N(_13166_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][30]$_DFFE_PP_  (.CLK(clknet_leaf_769_clk),
    .RESET_B(net908),
    .D(_01001_),
    .Q_N(_13165_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][31]$_DFFE_PP_  (.CLK(clknet_leaf_695_clk),
    .RESET_B(net909),
    .D(_01002_),
    .Q_N(_13164_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_1084_clk),
    .RESET_B(net910),
    .D(_01003_),
    .Q_N(_13163_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_1075_clk),
    .RESET_B(net911),
    .D(_01004_),
    .Q_N(_13162_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_1148_clk),
    .RESET_B(net912),
    .D(_01005_),
    .Q_N(_13161_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net913),
    .D(_01006_),
    .Q_N(_13160_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net914),
    .D(_01007_),
    .Q_N(_13159_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_923_clk),
    .RESET_B(net915),
    .D(_01008_),
    .Q_N(_13158_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][9]$_DFFE_PP_  (.CLK(clknet_8_54_0_clk),
    .RESET_B(net916),
    .D(_01009_),
    .Q_N(_13157_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[19][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_1003_clk),
    .RESET_B(net917),
    .D(_01010_),
    .Q_N(_13156_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_1076_clk),
    .RESET_B(net918),
    .D(_01011_),
    .Q_N(_13155_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_835_clk),
    .RESET_B(net919),
    .D(_01012_),
    .Q_N(_13154_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net920),
    .D(_01013_),
    .Q_N(_13153_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_1020_clk),
    .RESET_B(net921),
    .D(_01014_),
    .Q_N(_13152_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_937_clk),
    .RESET_B(net922),
    .D(_01015_),
    .Q_N(_13151_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_1144_clk),
    .RESET_B(net923),
    .D(_01016_),
    .Q_N(_13150_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_1032_clk),
    .RESET_B(net924),
    .D(_01017_),
    .Q_N(_13149_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_1026_clk),
    .RESET_B(net925),
    .D(_01018_),
    .Q_N(_13148_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_1051_clk),
    .RESET_B(net926),
    .D(_01019_),
    .Q_N(_13147_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_707_clk),
    .RESET_B(net927),
    .D(_01020_),
    .Q_N(_13146_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net928),
    .D(_01021_),
    .Q_N(_13145_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_1053_clk),
    .RESET_B(net929),
    .D(_01022_),
    .Q_N(_13144_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_1054_clk),
    .RESET_B(net930),
    .D(_01023_),
    .Q_N(_13143_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_823_clk),
    .RESET_B(net931),
    .D(_01024_),
    .Q_N(_13142_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][23]$_DFFE_PP_  (.CLK(clknet_8_163_0_clk),
    .RESET_B(net932),
    .D(_01025_),
    .Q_N(_13141_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_834_clk),
    .RESET_B(net933),
    .D(_01026_),
    .Q_N(_13140_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_792_clk),
    .RESET_B(net934),
    .D(_01027_),
    .Q_N(_13139_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_723_clk),
    .RESET_B(net935),
    .D(_01028_),
    .Q_N(_13138_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_808_clk),
    .RESET_B(net936),
    .D(_01029_),
    .Q_N(_13137_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_711_clk),
    .RESET_B(net937),
    .D(_01030_),
    .Q_N(_13136_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_813_clk),
    .RESET_B(net938),
    .D(_01031_),
    .Q_N(_13135_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_1131_clk),
    .RESET_B(net939),
    .D(_01032_),
    .Q_N(_13134_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_688_clk),
    .RESET_B(net940),
    .D(_01033_),
    .Q_N(_13133_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_706_clk),
    .RESET_B(net941),
    .D(_01034_),
    .Q_N(_13132_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][3]$_DFFE_PP_  (.CLK(clknet_8_35_0_clk),
    .RESET_B(net942),
    .D(_01035_),
    .Q_N(_13131_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_1073_clk),
    .RESET_B(net943),
    .D(_01036_),
    .Q_N(_13130_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_1092_clk),
    .RESET_B(net944),
    .D(_01037_),
    .Q_N(_13129_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net945),
    .D(_01038_),
    .Q_N(_13128_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_1149_clk),
    .RESET_B(net946),
    .D(_01039_),
    .Q_N(_13127_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_960_clk),
    .RESET_B(net947),
    .D(_01040_),
    .Q_N(_13126_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_1149_clk),
    .RESET_B(net948),
    .D(_01041_),
    .Q_N(_13125_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[1][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_1045_clk),
    .RESET_B(net949),
    .D(_01042_),
    .Q_N(_13124_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_1081_clk),
    .RESET_B(net950),
    .D(_01043_),
    .Q_N(_13123_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_832_clk),
    .RESET_B(net951),
    .D(_01044_),
    .Q_N(_13122_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][12]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net952),
    .D(_01045_),
    .Q_N(_13121_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][13]$_DFFE_PP_  (.CLK(clknet_leaf_1018_clk),
    .RESET_B(net953),
    .D(_01046_),
    .Q_N(_13120_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][14]$_DFFE_PP_  (.CLK(clknet_leaf_942_clk),
    .RESET_B(net954),
    .D(_01047_),
    .Q_N(_13119_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][15]$_DFFE_PP_  (.CLK(clknet_8_35_0_clk),
    .RESET_B(net955),
    .D(_01048_),
    .Q_N(_13118_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][16]$_DFFE_PP_  (.CLK(clknet_leaf_1038_clk),
    .RESET_B(net956),
    .D(_01049_),
    .Q_N(_13117_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][17]$_DFFE_PP_  (.CLK(clknet_leaf_1021_clk),
    .RESET_B(net957),
    .D(_01050_),
    .Q_N(_13116_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][18]$_DFFE_PP_  (.CLK(clknet_leaf_927_clk),
    .RESET_B(net958),
    .D(_01051_),
    .Q_N(_13115_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][19]$_DFFE_PP_  (.CLK(clknet_leaf_704_clk),
    .RESET_B(net959),
    .D(_01052_),
    .Q_N(_13114_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net960),
    .D(_01053_),
    .Q_N(_13113_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][20]$_DFFE_PP_  (.CLK(clknet_leaf_905_clk),
    .RESET_B(net961),
    .D(_01054_),
    .Q_N(_13112_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][21]$_DFFE_PP_  (.CLK(clknet_8_143_0_clk),
    .RESET_B(net962),
    .D(_01055_),
    .Q_N(_13111_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][22]$_DFFE_PP_  (.CLK(clknet_leaf_849_clk),
    .RESET_B(net963),
    .D(_01056_),
    .Q_N(_13110_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][23]$_DFFE_PP_  (.CLK(clknet_leaf_849_clk),
    .RESET_B(net964),
    .D(_01057_),
    .Q_N(_13109_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][24]$_DFFE_PP_  (.CLK(clknet_leaf_834_clk),
    .RESET_B(net965),
    .D(_01058_),
    .Q_N(_13108_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][25]$_DFFE_PP_  (.CLK(clknet_leaf_815_clk),
    .RESET_B(net966),
    .D(_01059_),
    .Q_N(_13107_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][26]$_DFFE_PP_  (.CLK(clknet_leaf_724_clk),
    .RESET_B(net967),
    .D(_01060_),
    .Q_N(_13106_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][27]$_DFFE_PP_  (.CLK(clknet_leaf_807_clk),
    .RESET_B(net968),
    .D(_01061_),
    .Q_N(_13105_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][28]$_DFFE_PP_  (.CLK(clknet_8_231_0_clk),
    .RESET_B(net969),
    .D(_01062_),
    .Q_N(_13104_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][29]$_DFFE_PP_  (.CLK(clknet_leaf_813_clk),
    .RESET_B(net970),
    .D(_01063_),
    .Q_N(_13103_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_1140_clk),
    .RESET_B(net971),
    .D(_01064_),
    .Q_N(_13102_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][30]$_DFFE_PP_  (.CLK(clknet_leaf_687_clk),
    .RESET_B(net972),
    .D(_01065_),
    .Q_N(_13101_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][31]$_DFFE_PP_  (.CLK(clknet_leaf_705_clk),
    .RESET_B(net973),
    .D(_01066_),
    .Q_N(_13100_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_1084_clk),
    .RESET_B(net974),
    .D(_01067_),
    .Q_N(_13099_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_1062_clk),
    .RESET_B(net975),
    .D(_01068_),
    .Q_N(_13098_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_1145_clk),
    .RESET_B(net976),
    .D(_01069_),
    .Q_N(_13097_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net977),
    .D(_01070_),
    .Q_N(_13096_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][7]$_DFFE_PP_  (.CLK(clknet_8_55_0_clk),
    .RESET_B(net978),
    .D(_01071_),
    .Q_N(_13095_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_936_clk),
    .RESET_B(net979),
    .D(_01072_),
    .Q_N(_13094_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net980),
    .D(_01073_),
    .Q_N(_13093_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[20][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_1045_clk),
    .RESET_B(net981),
    .D(_01074_),
    .Q_N(_13092_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_1080_clk),
    .RESET_B(net982),
    .D(_01075_),
    .Q_N(_13091_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_833_clk),
    .RESET_B(net983),
    .D(_01076_),
    .Q_N(_13090_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][12]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net984),
    .D(_01077_),
    .Q_N(_13089_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][13]$_DFFE_PP_  (.CLK(clknet_leaf_1019_clk),
    .RESET_B(net985),
    .D(_01078_),
    .Q_N(_13088_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][14]$_DFFE_PP_  (.CLK(clknet_leaf_943_clk),
    .RESET_B(net986),
    .D(_01079_),
    .Q_N(_13087_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][15]$_DFFE_PP_  (.CLK(clknet_leaf_1099_clk),
    .RESET_B(net987),
    .D(_01080_),
    .Q_N(_13086_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][16]$_DFFE_PP_  (.CLK(clknet_leaf_1038_clk),
    .RESET_B(net988),
    .D(_01081_),
    .Q_N(_13085_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][17]$_DFFE_PP_  (.CLK(clknet_8_58_0_clk),
    .RESET_B(net989),
    .D(_01082_),
    .Q_N(_13084_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][18]$_DFFE_PP_  (.CLK(clknet_leaf_924_clk),
    .RESET_B(net990),
    .D(_01083_),
    .Q_N(_13083_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][19]$_DFFE_PP_  (.CLK(clknet_leaf_708_clk),
    .RESET_B(net991),
    .D(_01084_),
    .Q_N(_13082_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net992),
    .D(_01085_),
    .Q_N(_13081_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][20]$_DFFE_PP_  (.CLK(clknet_leaf_930_clk),
    .RESET_B(net993),
    .D(_01086_),
    .Q_N(_13080_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][21]$_DFFE_PP_  (.CLK(clknet_leaf_932_clk),
    .RESET_B(net994),
    .D(_01087_),
    .Q_N(_13079_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][22]$_DFFE_PP_  (.CLK(clknet_leaf_848_clk),
    .RESET_B(net995),
    .D(_01088_),
    .Q_N(_13078_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][23]$_DFFE_PP_  (.CLK(clknet_leaf_851_clk),
    .RESET_B(net996),
    .D(_01089_),
    .Q_N(_13077_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][24]$_DFFE_PP_  (.CLK(clknet_leaf_847_clk),
    .RESET_B(net997),
    .D(_01090_),
    .Q_N(_13076_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][25]$_DFFE_PP_  (.CLK(clknet_leaf_815_clk),
    .RESET_B(net998),
    .D(_01091_),
    .Q_N(_13075_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][26]$_DFFE_PP_  (.CLK(clknet_8_236_0_clk),
    .RESET_B(net999),
    .D(_01092_),
    .Q_N(_13074_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][27]$_DFFE_PP_  (.CLK(clknet_leaf_810_clk),
    .RESET_B(net1000),
    .D(_01093_),
    .Q_N(_13073_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][28]$_DFFE_PP_  (.CLK(clknet_leaf_602_clk),
    .RESET_B(net1001),
    .D(_01094_),
    .Q_N(_13072_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][29]$_DFFE_PP_  (.CLK(clknet_8_184_0_clk),
    .RESET_B(net1002),
    .D(_01095_),
    .Q_N(_13071_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_1140_clk),
    .RESET_B(net1003),
    .D(_01096_),
    .Q_N(_13070_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][30]$_DFFE_PP_  (.CLK(clknet_leaf_688_clk),
    .RESET_B(net1004),
    .D(_01097_),
    .Q_N(_13069_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][31]$_DFFE_PP_  (.CLK(clknet_leaf_705_clk),
    .RESET_B(net1005),
    .D(_01098_),
    .Q_N(_13068_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_1083_clk),
    .RESET_B(net1006),
    .D(_01099_),
    .Q_N(_13067_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_1062_clk),
    .RESET_B(net1007),
    .D(_01100_),
    .Q_N(_13066_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_1146_clk),
    .RESET_B(net1008),
    .D(_01101_),
    .Q_N(_13065_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1009),
    .D(_01102_),
    .Q_N(_13064_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][7]$_DFFE_PP_  (.CLK(clknet_8_49_0_clk),
    .RESET_B(net1010),
    .D(_01103_),
    .Q_N(_13063_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_936_clk),
    .RESET_B(net1011),
    .D(_01104_),
    .Q_N(_13062_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][9]$_DFFE_PP_  (.CLK(clknet_8_49_0_clk),
    .RESET_B(net1012),
    .D(_01105_),
    .Q_N(_13061_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[21][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_1044_clk),
    .RESET_B(net1013),
    .D(_01106_),
    .Q_N(_13060_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_1080_clk),
    .RESET_B(net1014),
    .D(_01107_),
    .Q_N(_13059_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_829_clk),
    .RESET_B(net1015),
    .D(_01108_),
    .Q_N(_13058_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][12]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1016),
    .D(_01109_),
    .Q_N(_13057_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][13]$_DFFE_PP_  (.CLK(clknet_leaf_1027_clk),
    .RESET_B(net1017),
    .D(_01110_),
    .Q_N(_13056_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][14]$_DFFE_PP_  (.CLK(clknet_leaf_681_clk),
    .RESET_B(net1018),
    .D(_01111_),
    .Q_N(_13055_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][15]$_DFFE_PP_  (.CLK(clknet_8_33_0_clk),
    .RESET_B(net1019),
    .D(_01112_),
    .Q_N(_13054_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][16]$_DFFE_PP_  (.CLK(clknet_8_144_0_clk),
    .RESET_B(net1020),
    .D(_01113_),
    .Q_N(_13053_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][17]$_DFFE_PP_  (.CLK(clknet_leaf_1019_clk),
    .RESET_B(net1021),
    .D(_01114_),
    .Q_N(_13052_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][18]$_DFFE_PP_  (.CLK(clknet_leaf_931_clk),
    .RESET_B(net1022),
    .D(_01115_),
    .Q_N(_13051_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][19]$_DFFE_PP_  (.CLK(clknet_leaf_603_clk),
    .RESET_B(net1023),
    .D(_01116_),
    .Q_N(_13050_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1024),
    .D(_01117_),
    .Q_N(_13049_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][20]$_DFFE_PP_  (.CLK(clknet_leaf_930_clk),
    .RESET_B(net1025),
    .D(_01118_),
    .Q_N(_13048_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][21]$_DFFE_PP_  (.CLK(clknet_leaf_931_clk),
    .RESET_B(net1026),
    .D(_01119_),
    .Q_N(_13047_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][22]$_DFFE_PP_  (.CLK(clknet_leaf_848_clk),
    .RESET_B(net1027),
    .D(_01120_),
    .Q_N(_13046_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][23]$_DFFE_PP_  (.CLK(clknet_leaf_851_clk),
    .RESET_B(net1028),
    .D(_01121_),
    .Q_N(_13045_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][24]$_DFFE_PP_  (.CLK(clknet_leaf_845_clk),
    .RESET_B(net1029),
    .D(_01122_),
    .Q_N(_13044_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][25]$_DFFE_PP_  (.CLK(clknet_leaf_816_clk),
    .RESET_B(net1030),
    .D(_01123_),
    .Q_N(_13043_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][26]$_DFFE_PP_  (.CLK(clknet_leaf_596_clk),
    .RESET_B(net1031),
    .D(_01124_),
    .Q_N(_13042_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][27]$_DFFE_PP_  (.CLK(clknet_leaf_810_clk),
    .RESET_B(net1032),
    .D(_01125_),
    .Q_N(_13041_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][28]$_DFFE_PP_  (.CLK(clknet_leaf_602_clk),
    .RESET_B(net1033),
    .D(_01126_),
    .Q_N(_13040_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][29]$_DFFE_PP_  (.CLK(clknet_leaf_817_clk),
    .RESET_B(net1034),
    .D(_01127_),
    .Q_N(_13039_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_1140_clk),
    .RESET_B(net1035),
    .D(_01128_),
    .Q_N(_13038_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][30]$_DFFE_PP_  (.CLK(clknet_leaf_687_clk),
    .RESET_B(net1036),
    .D(_01129_),
    .Q_N(_13037_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][31]$_DFFE_PP_  (.CLK(clknet_leaf_704_clk),
    .RESET_B(net1037),
    .D(_01130_),
    .Q_N(_13036_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_1083_clk),
    .RESET_B(net1038),
    .D(_01131_),
    .Q_N(_13035_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_1063_clk),
    .RESET_B(net1039),
    .D(_01132_),
    .Q_N(_13034_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_1147_clk),
    .RESET_B(net1040),
    .D(_01133_),
    .Q_N(_13033_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1041),
    .D(_01134_),
    .Q_N(_13032_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1042),
    .D(_01135_),
    .Q_N(_13031_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_921_clk),
    .RESET_B(net1043),
    .D(_01136_),
    .Q_N(_13030_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1044),
    .D(_01137_),
    .Q_N(_13029_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[22][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_1049_clk),
    .RESET_B(net1045),
    .D(_01138_),
    .Q_N(_13028_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_1081_clk),
    .RESET_B(net1046),
    .D(_01139_),
    .Q_N(_13027_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_829_clk),
    .RESET_B(net1047),
    .D(_01140_),
    .Q_N(_13026_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][12]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1048),
    .D(_01141_),
    .Q_N(_13025_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][13]$_DFFE_PP_  (.CLK(clknet_leaf_1028_clk),
    .RESET_B(net1049),
    .D(_01142_),
    .Q_N(_13024_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][14]$_DFFE_PP_  (.CLK(clknet_leaf_943_clk),
    .RESET_B(net1050),
    .D(_01143_),
    .Q_N(_13023_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][15]$_DFFE_PP_  (.CLK(clknet_leaf_1099_clk),
    .RESET_B(net1051),
    .D(_01144_),
    .Q_N(_13022_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][16]$_DFFE_PP_  (.CLK(clknet_leaf_1044_clk),
    .RESET_B(net1052),
    .D(_01145_),
    .Q_N(_13021_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][17]$_DFFE_PP_  (.CLK(clknet_leaf_1021_clk),
    .RESET_B(net1053),
    .D(_01146_),
    .Q_N(_13020_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][18]$_DFFE_PP_  (.CLK(clknet_leaf_934_clk),
    .RESET_B(net1054),
    .D(_01147_),
    .Q_N(_13019_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][19]$_DFFE_PP_  (.CLK(clknet_leaf_603_clk),
    .RESET_B(net1055),
    .D(_01148_),
    .Q_N(_13018_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1056),
    .D(_01149_),
    .Q_N(_13017_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][20]$_DFFE_PP_  (.CLK(clknet_leaf_929_clk),
    .RESET_B(net1057),
    .D(_01150_),
    .Q_N(_13016_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][21]$_DFFE_PP_  (.CLK(clknet_leaf_932_clk),
    .RESET_B(net1058),
    .D(_01151_),
    .Q_N(_13015_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][22]$_DFFE_PP_  (.CLK(clknet_leaf_847_clk),
    .RESET_B(net1059),
    .D(_01152_),
    .Q_N(_13014_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][23]$_DFFE_PP_  (.CLK(clknet_leaf_850_clk),
    .RESET_B(net1060),
    .D(_01153_),
    .Q_N(_13013_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][24]$_DFFE_PP_  (.CLK(clknet_leaf_835_clk),
    .RESET_B(net1061),
    .D(_01154_),
    .Q_N(_13012_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][25]$_DFFE_PP_  (.CLK(clknet_leaf_814_clk),
    .RESET_B(net1062),
    .D(_01155_),
    .Q_N(_13011_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][26]$_DFFE_PP_  (.CLK(clknet_leaf_596_clk),
    .RESET_B(net1063),
    .D(_01156_),
    .Q_N(_13010_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][27]$_DFFE_PP_  (.CLK(clknet_8_186_0_clk),
    .RESET_B(net1064),
    .D(_01157_),
    .Q_N(_13009_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][28]$_DFFE_PP_  (.CLK(clknet_leaf_602_clk),
    .RESET_B(net1065),
    .D(_01158_),
    .Q_N(_13008_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][29]$_DFFE_PP_  (.CLK(clknet_leaf_811_clk),
    .RESET_B(net1066),
    .D(_01159_),
    .Q_N(_13007_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_1145_clk),
    .RESET_B(net1067),
    .D(_01160_),
    .Q_N(_13006_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][30]$_DFFE_PP_  (.CLK(clknet_8_224_0_clk),
    .RESET_B(net1068),
    .D(_01161_),
    .Q_N(_13005_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][31]$_DFFE_PP_  (.CLK(clknet_leaf_706_clk),
    .RESET_B(net1069),
    .D(_01162_),
    .Q_N(_13004_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_1061_clk),
    .RESET_B(net1070),
    .D(_01163_),
    .Q_N(_13003_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_1063_clk),
    .RESET_B(net1071),
    .D(_01164_),
    .Q_N(_13002_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_1146_clk),
    .RESET_B(net1072),
    .D(_01165_),
    .Q_N(_13001_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1073),
    .D(_01166_),
    .Q_N(_13000_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1074),
    .D(_01167_),
    .Q_N(_12999_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_936_clk),
    .RESET_B(net1075),
    .D(_01168_),
    .Q_N(_12998_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1076),
    .D(_01169_),
    .Q_N(_12997_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[23][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_1003_clk),
    .RESET_B(net1077),
    .D(_01170_),
    .Q_N(_12996_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_1060_clk),
    .RESET_B(net1078),
    .D(_01171_),
    .Q_N(_12995_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_831_clk),
    .RESET_B(net1079),
    .D(_01172_),
    .Q_N(_12994_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][12]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1080),
    .D(_01173_),
    .Q_N(_12993_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][13]$_DFFE_PP_  (.CLK(clknet_8_63_0_clk),
    .RESET_B(net1081),
    .D(_01174_),
    .Q_N(_12992_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][14]$_DFFE_PP_  (.CLK(clknet_8_158_0_clk),
    .RESET_B(net1082),
    .D(_01175_),
    .Q_N(_12991_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][15]$_DFFE_PP_  (.CLK(clknet_leaf_1138_clk),
    .RESET_B(net1083),
    .D(_01176_),
    .Q_N(_12990_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][16]$_DFFE_PP_  (.CLK(clknet_leaf_1056_clk),
    .RESET_B(net1084),
    .D(_01177_),
    .Q_N(_12989_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][17]$_DFFE_PP_  (.CLK(clknet_8_62_0_clk),
    .RESET_B(net1085),
    .D(_01178_),
    .Q_N(_12988_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][18]$_DFFE_PP_  (.CLK(clknet_8_153_0_clk),
    .RESET_B(net1086),
    .D(_01179_),
    .Q_N(_12987_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][19]$_DFFE_PP_  (.CLK(clknet_8_191_0_clk),
    .RESET_B(net1087),
    .D(_01180_),
    .Q_N(_12986_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1088),
    .D(_01181_),
    .Q_N(_12985_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][20]$_DFFE_PP_  (.CLK(clknet_leaf_884_clk),
    .RESET_B(net1089),
    .D(_01182_),
    .Q_N(_12984_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][21]$_DFFE_PP_  (.CLK(clknet_leaf_893_clk),
    .RESET_B(net1090),
    .D(_01183_),
    .Q_N(_12983_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][22]$_DFFE_PP_  (.CLK(clknet_leaf_870_clk),
    .RESET_B(net1091),
    .D(_01184_),
    .Q_N(_12982_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][23]$_DFFE_PP_  (.CLK(clknet_leaf_884_clk),
    .RESET_B(net1092),
    .D(_01185_),
    .Q_N(_12981_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][24]$_DFFE_PP_  (.CLK(clknet_leaf_867_clk),
    .RESET_B(net1093),
    .D(_01186_),
    .Q_N(_12980_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][25]$_DFFE_PP_  (.CLK(clknet_8_182_0_clk),
    .RESET_B(net1094),
    .D(_01187_),
    .Q_N(_12979_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][26]$_DFFE_PP_  (.CLK(clknet_leaf_731_clk),
    .RESET_B(net1095),
    .D(_01188_),
    .Q_N(_12978_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][27]$_DFFE_PP_  (.CLK(clknet_leaf_754_clk),
    .RESET_B(net1096),
    .D(_01189_),
    .Q_N(_12977_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][28]$_DFFE_PP_  (.CLK(clknet_leaf_730_clk),
    .RESET_B(net1097),
    .D(_01190_),
    .Q_N(_12976_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][29]$_DFFE_PP_  (.CLK(clknet_leaf_789_clk),
    .RESET_B(net1098),
    .D(_01191_),
    .Q_N(_12975_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1099),
    .D(_01192_),
    .Q_N(_12974_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][30]$_DFFE_PP_  (.CLK(clknet_leaf_777_clk),
    .RESET_B(net1100),
    .D(_01193_),
    .Q_N(_12973_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][31]$_DFFE_PP_  (.CLK(clknet_leaf_680_clk),
    .RESET_B(net1101),
    .D(_01194_),
    .Q_N(_12972_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_1061_clk),
    .RESET_B(net1102),
    .D(_01195_),
    .Q_N(_12971_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][4]$_DFFE_PP_  (.CLK(clknet_8_132_0_clk),
    .RESET_B(net1103),
    .D(_01196_),
    .Q_N(_12970_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1104),
    .D(_01197_),
    .Q_N(_12969_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1105),
    .D(_01198_),
    .Q_N(_12968_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1106),
    .D(_01199_),
    .Q_N(_12967_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_963_clk),
    .RESET_B(net1107),
    .D(_01200_),
    .Q_N(_12966_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1108),
    .D(_01201_),
    .Q_N(_12965_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[24][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_1009_clk),
    .RESET_B(net1109),
    .D(_01202_),
    .Q_N(_12964_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][10]$_DFFE_PP_  (.CLK(clknet_8_43_0_clk),
    .RESET_B(net1110),
    .D(_01203_),
    .Q_N(_12963_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][11]$_DFFE_PP_  (.CLK(clknet_8_175_0_clk),
    .RESET_B(net1111),
    .D(_01204_),
    .Q_N(_12962_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][12]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1112),
    .D(_01205_),
    .Q_N(_12961_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][13]$_DFFE_PP_  (.CLK(clknet_leaf_1012_clk),
    .RESET_B(net1113),
    .D(_01206_),
    .Q_N(_12960_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][14]$_DFFE_PP_  (.CLK(clknet_leaf_949_clk),
    .RESET_B(net1114),
    .D(_01207_),
    .Q_N(_12959_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][15]$_DFFE_PP_  (.CLK(clknet_leaf_1138_clk),
    .RESET_B(net1115),
    .D(_01208_),
    .Q_N(_12958_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][16]$_DFFE_PP_  (.CLK(clknet_leaf_1038_clk),
    .RESET_B(net1116),
    .D(_01209_),
    .Q_N(_12957_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][17]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1117),
    .D(_01210_),
    .Q_N(_12956_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][18]$_DFFE_PP_  (.CLK(clknet_leaf_916_clk),
    .RESET_B(net1118),
    .D(_01211_),
    .Q_N(_12955_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][19]$_DFFE_PP_  (.CLK(clknet_leaf_750_clk),
    .RESET_B(net1119),
    .D(_01212_),
    .Q_N(_12954_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1120),
    .D(_01213_),
    .Q_N(_12953_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][20]$_DFFE_PP_  (.CLK(clknet_leaf_887_clk),
    .RESET_B(net1121),
    .D(_01214_),
    .Q_N(_12952_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][21]$_DFFE_PP_  (.CLK(clknet_leaf_893_clk),
    .RESET_B(net1122),
    .D(_01215_),
    .Q_N(_12951_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][22]$_DFFE_PP_  (.CLK(clknet_leaf_873_clk),
    .RESET_B(net1123),
    .D(_01216_),
    .Q_N(_12950_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][23]$_DFFE_PP_  (.CLK(clknet_leaf_882_clk),
    .RESET_B(net1124),
    .D(_01217_),
    .Q_N(_12949_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][24]$_DFFE_PP_  (.CLK(clknet_leaf_867_clk),
    .RESET_B(net1125),
    .D(_01218_),
    .Q_N(_12948_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][25]$_DFFE_PP_  (.CLK(clknet_8_182_0_clk),
    .RESET_B(net1126),
    .D(_01219_),
    .Q_N(_12947_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][26]$_DFFE_PP_  (.CLK(clknet_leaf_736_clk),
    .RESET_B(net1127),
    .D(_01220_),
    .Q_N(_12946_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][27]$_DFFE_PP_  (.CLK(clknet_leaf_752_clk),
    .RESET_B(net1128),
    .D(_01221_),
    .Q_N(_12945_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][28]$_DFFE_PP_  (.CLK(clknet_leaf_730_clk),
    .RESET_B(net1129),
    .D(_01222_),
    .Q_N(_12944_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][29]$_DFFE_PP_  (.CLK(clknet_leaf_788_clk),
    .RESET_B(net1130),
    .D(_01223_),
    .Q_N(_12943_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1131),
    .D(_01224_),
    .Q_N(_12942_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][30]$_DFFE_PP_  (.CLK(clknet_leaf_771_clk),
    .RESET_B(net1132),
    .D(_01225_),
    .Q_N(_12941_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][31]$_DFFE_PP_  (.CLK(clknet_leaf_680_clk),
    .RESET_B(net1133),
    .D(_01226_),
    .Q_N(_12940_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_1060_clk),
    .RESET_B(net1134),
    .D(_01227_),
    .Q_N(_12939_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_1065_clk),
    .RESET_B(net1135),
    .D(_01228_),
    .Q_N(_12938_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1136),
    .D(_01229_),
    .Q_N(_12937_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1137),
    .D(_01230_),
    .Q_N(_12936_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1138),
    .D(_01231_),
    .Q_N(_12935_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_962_clk),
    .RESET_B(net1139),
    .D(_01232_),
    .Q_N(_12934_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][9]$_DFFE_PP_  (.CLK(clknet_8_12_0_clk),
    .RESET_B(net1140),
    .D(_01233_),
    .Q_N(_12933_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[25][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_1010_clk),
    .RESET_B(net1141),
    .D(_01234_),
    .Q_N(_12932_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_1055_clk),
    .RESET_B(net1142),
    .D(_01235_),
    .Q_N(_12931_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_788_clk),
    .RESET_B(net1143),
    .D(_01236_),
    .Q_N(_12930_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][12]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1144),
    .D(_01237_),
    .Q_N(_12929_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][13]$_DFFE_PP_  (.CLK(clknet_leaf_1012_clk),
    .RESET_B(net1145),
    .D(_01238_),
    .Q_N(_12928_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][14]$_DFFE_PP_  (.CLK(clknet_leaf_953_clk),
    .RESET_B(net1146),
    .D(_01239_),
    .Q_N(_12927_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][15]$_DFFE_PP_  (.CLK(clknet_leaf_1139_clk),
    .RESET_B(net1147),
    .D(_01240_),
    .Q_N(_12926_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][16]$_DFFE_PP_  (.CLK(clknet_leaf_1057_clk),
    .RESET_B(net1148),
    .D(_01241_),
    .Q_N(_12925_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][17]$_DFFE_PP_  (.CLK(clknet_leaf_1017_clk),
    .RESET_B(net1149),
    .D(_01242_),
    .Q_N(_12924_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][18]$_DFFE_PP_  (.CLK(clknet_8_152_0_clk),
    .RESET_B(net1150),
    .D(_01243_),
    .Q_N(_12923_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][19]$_DFFE_PP_  (.CLK(clknet_leaf_748_clk),
    .RESET_B(net1151),
    .D(_01244_),
    .Q_N(_12922_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][1]$_DFFE_PP_  (.CLK(clknet_8_14_0_clk),
    .RESET_B(net1152),
    .D(_01245_),
    .Q_N(_12921_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][20]$_DFFE_PP_  (.CLK(clknet_leaf_887_clk),
    .RESET_B(net1153),
    .D(_01246_),
    .Q_N(_12920_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][21]$_DFFE_PP_  (.CLK(clknet_leaf_894_clk),
    .RESET_B(net1154),
    .D(_01247_),
    .Q_N(_12919_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][22]$_DFFE_PP_  (.CLK(clknet_8_138_0_clk),
    .RESET_B(net1155),
    .D(_01248_),
    .Q_N(_12918_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][23]$_DFFE_PP_  (.CLK(clknet_leaf_882_clk),
    .RESET_B(net1156),
    .D(_01249_),
    .Q_N(_12917_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][24]$_DFFE_PP_  (.CLK(clknet_8_168_0_clk),
    .RESET_B(net1157),
    .D(_01250_),
    .Q_N(_12916_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][25]$_DFFE_PP_  (.CLK(clknet_leaf_772_clk),
    .RESET_B(net1158),
    .D(_01251_),
    .Q_N(_12915_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][26]$_DFFE_PP_  (.CLK(clknet_leaf_733_clk),
    .RESET_B(net1159),
    .D(_01252_),
    .Q_N(_12914_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][27]$_DFFE_PP_  (.CLK(clknet_leaf_753_clk),
    .RESET_B(net1160),
    .D(_01253_),
    .Q_N(_12913_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][28]$_DFFE_PP_  (.CLK(clknet_leaf_730_clk),
    .RESET_B(net1161),
    .D(_01254_),
    .Q_N(_12912_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][29]$_DFFE_PP_  (.CLK(clknet_leaf_790_clk),
    .RESET_B(net1162),
    .D(_01255_),
    .Q_N(_12911_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][2]$_DFFE_PP_  (.CLK(clknet_8_48_0_clk),
    .RESET_B(net1163),
    .D(_01256_),
    .Q_N(_12910_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][30]$_DFFE_PP_  (.CLK(clknet_8_181_0_clk),
    .RESET_B(net1164),
    .D(_01257_),
    .Q_N(_12909_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][31]$_DFFE_PP_  (.CLK(clknet_leaf_684_clk),
    .RESET_B(net1165),
    .D(_01258_),
    .Q_N(_12908_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_1058_clk),
    .RESET_B(net1166),
    .D(_01259_),
    .Q_N(_12907_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_1055_clk),
    .RESET_B(net1167),
    .D(_01260_),
    .Q_N(_12906_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][5]$_DFFE_PP_  (.CLK(clknet_8_48_0_clk),
    .RESET_B(net1168),
    .D(_01261_),
    .Q_N(_12905_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1169),
    .D(_01262_),
    .Q_N(_12904_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1170),
    .D(_01263_),
    .Q_N(_12903_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_963_clk),
    .RESET_B(net1171),
    .D(_01264_),
    .Q_N(_12902_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1172),
    .D(_01265_),
    .Q_N(_12901_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[26][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_997_clk),
    .RESET_B(net1173),
    .D(_01266_),
    .Q_N(_12900_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_1058_clk),
    .RESET_B(net1174),
    .D(_01267_),
    .Q_N(_12899_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_788_clk),
    .RESET_B(net1175),
    .D(_01268_),
    .Q_N(_12898_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][12]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1176),
    .D(_01269_),
    .Q_N(_12897_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][13]$_DFFE_PP_  (.CLK(clknet_leaf_1011_clk),
    .RESET_B(net1177),
    .D(_01270_),
    .Q_N(_12896_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][14]$_DFFE_PP_  (.CLK(clknet_leaf_952_clk),
    .RESET_B(net1178),
    .D(_01271_),
    .Q_N(_12895_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][15]$_DFFE_PP_  (.CLK(clknet_leaf_1139_clk),
    .RESET_B(net1179),
    .D(_01272_),
    .Q_N(_12894_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][16]$_DFFE_PP_  (.CLK(clknet_leaf_1056_clk),
    .RESET_B(net1180),
    .D(_01273_),
    .Q_N(_12893_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][17]$_DFFE_PP_  (.CLK(clknet_8_63_0_clk),
    .RESET_B(net1181),
    .D(_01274_),
    .Q_N(_12892_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][18]$_DFFE_PP_  (.CLK(clknet_leaf_917_clk),
    .RESET_B(net1182),
    .D(_01275_),
    .Q_N(_12891_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][19]$_DFFE_PP_  (.CLK(clknet_leaf_749_clk),
    .RESET_B(net1183),
    .D(_01276_),
    .Q_N(_12890_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1184),
    .D(_01277_),
    .Q_N(_12889_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][20]$_DFFE_PP_  (.CLK(clknet_leaf_882_clk),
    .RESET_B(net1185),
    .D(_01278_),
    .Q_N(_12888_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][21]$_DFFE_PP_  (.CLK(clknet_8_137_0_clk),
    .RESET_B(net1186),
    .D(_01279_),
    .Q_N(_12887_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][22]$_DFFE_PP_  (.CLK(clknet_leaf_874_clk),
    .RESET_B(net1187),
    .D(_01280_),
    .Q_N(_12886_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][23]$_DFFE_PP_  (.CLK(clknet_leaf_873_clk),
    .RESET_B(net1188),
    .D(_01281_),
    .Q_N(_12885_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][24]$_DFFE_PP_  (.CLK(clknet_leaf_863_clk),
    .RESET_B(net1189),
    .D(_01282_),
    .Q_N(_12884_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][25]$_DFFE_PP_  (.CLK(clknet_8_188_0_clk),
    .RESET_B(net1190),
    .D(_01283_),
    .Q_N(_12883_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][26]$_DFFE_PP_  (.CLK(clknet_leaf_733_clk),
    .RESET_B(net1191),
    .D(_01284_),
    .Q_N(_12882_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][27]$_DFFE_PP_  (.CLK(clknet_leaf_753_clk),
    .RESET_B(net1192),
    .D(_01285_),
    .Q_N(_12881_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][28]$_DFFE_PP_  (.CLK(clknet_leaf_728_clk),
    .RESET_B(net1193),
    .D(_01286_),
    .Q_N(_12880_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][29]$_DFFE_PP_  (.CLK(clknet_leaf_787_clk),
    .RESET_B(net1194),
    .D(_01287_),
    .Q_N(_12879_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_1136_clk),
    .RESET_B(net1195),
    .D(_01288_),
    .Q_N(_12878_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][30]$_DFFE_PP_  (.CLK(clknet_leaf_771_clk),
    .RESET_B(net1196),
    .D(_01289_),
    .Q_N(_12877_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][31]$_DFFE_PP_  (.CLK(clknet_leaf_680_clk),
    .RESET_B(net1197),
    .D(_01290_),
    .Q_N(_12876_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_1065_clk),
    .RESET_B(net1198),
    .D(_01291_),
    .Q_N(_12875_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_1066_clk),
    .RESET_B(net1199),
    .D(_01292_),
    .Q_N(_12874_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1200),
    .D(_01293_),
    .Q_N(_12873_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1201),
    .D(_01294_),
    .Q_N(_12872_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1202),
    .D(_01295_),
    .Q_N(_12871_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_962_clk),
    .RESET_B(net1203),
    .D(_01296_),
    .Q_N(_12870_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1204),
    .D(_01297_),
    .Q_N(_12869_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[27][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_999_clk),
    .RESET_B(net1205),
    .D(_01298_),
    .Q_N(_12868_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_1034_clk),
    .RESET_B(net1206),
    .D(_01299_),
    .Q_N(_12867_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][11]$_DFFE_PP_  (.CLK(clknet_8_174_0_clk),
    .RESET_B(net1207),
    .D(_01300_),
    .Q_N(_12866_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][12]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1208),
    .D(_01301_),
    .Q_N(_12865_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][13]$_DFFE_PP_  (.CLK(clknet_8_149_0_clk),
    .RESET_B(net1209),
    .D(_01302_),
    .Q_N(_12864_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][14]$_DFFE_PP_  (.CLK(clknet_leaf_672_clk),
    .RESET_B(net1210),
    .D(_01303_),
    .Q_N(_12863_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][15]$_DFFE_PP_  (.CLK(clknet_leaf_1122_clk),
    .RESET_B(net1211),
    .D(_01304_),
    .Q_N(_12862_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][16]$_DFFE_PP_  (.CLK(clknet_8_146_0_clk),
    .RESET_B(net1212),
    .D(_01305_),
    .Q_N(_12861_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][17]$_DFFE_PP_  (.CLK(clknet_8_62_0_clk),
    .RESET_B(net1213),
    .D(_01306_),
    .Q_N(_12860_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][18]$_DFFE_PP_  (.CLK(clknet_leaf_1048_clk),
    .RESET_B(net1214),
    .D(_01307_),
    .Q_N(_12859_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][19]$_DFFE_PP_  (.CLK(clknet_leaf_747_clk),
    .RESET_B(net1215),
    .D(_01308_),
    .Q_N(_12858_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1216),
    .D(_01309_),
    .Q_N(_12857_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][20]$_DFFE_PP_  (.CLK(clknet_leaf_902_clk),
    .RESET_B(net1217),
    .D(_01310_),
    .Q_N(_12856_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][21]$_DFFE_PP_  (.CLK(clknet_leaf_898_clk),
    .RESET_B(net1218),
    .D(_01311_),
    .Q_N(_12855_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][22]$_DFFE_PP_  (.CLK(clknet_leaf_875_clk),
    .RESET_B(net1219),
    .D(_01312_),
    .Q_N(_12854_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][23]$_DFFE_PP_  (.CLK(clknet_leaf_879_clk),
    .RESET_B(net1220),
    .D(_01313_),
    .Q_N(_12853_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][24]$_DFFE_PP_  (.CLK(clknet_8_161_0_clk),
    .RESET_B(net1221),
    .D(_01314_),
    .Q_N(_12852_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][25]$_DFFE_PP_  (.CLK(clknet_leaf_765_clk),
    .RESET_B(net1222),
    .D(_01315_),
    .Q_N(_12851_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][26]$_DFFE_PP_  (.CLK(clknet_leaf_736_clk),
    .RESET_B(net1223),
    .D(_01316_),
    .Q_N(_12850_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][27]$_DFFE_PP_  (.CLK(clknet_leaf_750_clk),
    .RESET_B(net1224),
    .D(_01317_),
    .Q_N(_12849_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][28]$_DFFE_PP_  (.CLK(clknet_leaf_731_clk),
    .RESET_B(net1225),
    .D(_01318_),
    .Q_N(_12848_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][29]$_DFFE_PP_  (.CLK(clknet_leaf_791_clk),
    .RESET_B(net1226),
    .D(_01319_),
    .Q_N(_12847_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_1136_clk),
    .RESET_B(net1227),
    .D(_01320_),
    .Q_N(_12846_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][30]$_DFFE_PP_  (.CLK(clknet_leaf_770_clk),
    .RESET_B(net1228),
    .D(_01321_),
    .Q_N(_12845_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][31]$_DFFE_PP_  (.CLK(clknet_leaf_677_clk),
    .RESET_B(net1229),
    .D(_01322_),
    .Q_N(_12844_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_1037_clk),
    .RESET_B(net1230),
    .D(_01323_),
    .Q_N(_12843_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_1066_clk),
    .RESET_B(net1231),
    .D(_01324_),
    .Q_N(_12842_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1232),
    .D(_01325_),
    .Q_N(_12841_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1233),
    .D(_01326_),
    .Q_N(_12840_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][7]$_DFFE_PP_  (.CLK(clknet_8_13_0_clk),
    .RESET_B(net1234),
    .D(_01327_),
    .Q_N(_12839_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_956_clk),
    .RESET_B(net1235),
    .D(_01328_),
    .Q_N(_12838_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1236),
    .D(_01329_),
    .Q_N(_12837_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[28][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_1000_clk),
    .RESET_B(net1237),
    .D(_01330_),
    .Q_N(_12836_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_1035_clk),
    .RESET_B(net1238),
    .D(_01331_),
    .Q_N(_12835_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_789_clk),
    .RESET_B(net1239),
    .D(_01332_),
    .Q_N(_12834_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][12]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1240),
    .D(_01333_),
    .Q_N(_12833_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][13]$_DFFE_PP_  (.CLK(clknet_leaf_1010_clk),
    .RESET_B(net1241),
    .D(_01334_),
    .Q_N(_12832_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][14]$_DFFE_PP_  (.CLK(clknet_leaf_679_clk),
    .RESET_B(net1242),
    .D(_01335_),
    .Q_N(_12831_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][15]$_DFFE_PP_  (.CLK(clknet_leaf_1113_clk),
    .RESET_B(net1243),
    .D(_01336_),
    .Q_N(_12830_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][16]$_DFFE_PP_  (.CLK(clknet_leaf_1055_clk),
    .RESET_B(net1244),
    .D(_01337_),
    .Q_N(_12829_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][17]$_DFFE_PP_  (.CLK(clknet_8_61_0_clk),
    .RESET_B(net1245),
    .D(_01338_),
    .Q_N(_12828_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][18]$_DFFE_PP_  (.CLK(clknet_leaf_916_clk),
    .RESET_B(net1246),
    .D(_01339_),
    .Q_N(_12827_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][19]$_DFFE_PP_  (.CLK(clknet_leaf_747_clk),
    .RESET_B(net1247),
    .D(_01340_),
    .Q_N(_12826_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1248),
    .D(_01341_),
    .Q_N(_12825_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][20]$_DFFE_PP_  (.CLK(clknet_leaf_902_clk),
    .RESET_B(net1249),
    .D(_01342_),
    .Q_N(_12824_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][21]$_DFFE_PP_  (.CLK(clknet_leaf_899_clk),
    .RESET_B(net1250),
    .D(_01343_),
    .Q_N(_12823_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][22]$_DFFE_PP_  (.CLK(clknet_leaf_875_clk),
    .RESET_B(net1251),
    .D(_01344_),
    .Q_N(_12822_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][23]$_DFFE_PP_  (.CLK(clknet_leaf_878_clk),
    .RESET_B(net1252),
    .D(_01345_),
    .Q_N(_12821_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][24]$_DFFE_PP_  (.CLK(clknet_leaf_854_clk),
    .RESET_B(net1253),
    .D(_01346_),
    .Q_N(_12820_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][25]$_DFFE_PP_  (.CLK(clknet_leaf_759_clk),
    .RESET_B(net1254),
    .D(_01347_),
    .Q_N(_12819_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][26]$_DFFE_PP_  (.CLK(clknet_leaf_734_clk),
    .RESET_B(net1255),
    .D(_01348_),
    .Q_N(_12818_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][27]$_DFFE_PP_  (.CLK(clknet_leaf_749_clk),
    .RESET_B(net1256),
    .D(_01349_),
    .Q_N(_12817_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][28]$_DFFE_PP_  (.CLK(clknet_8_235_0_clk),
    .RESET_B(net1257),
    .D(_01350_),
    .Q_N(_12816_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][29]$_DFFE_PP_  (.CLK(clknet_leaf_790_clk),
    .RESET_B(net1258),
    .D(_01351_),
    .Q_N(_12815_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_1133_clk),
    .RESET_B(net1259),
    .D(_01352_),
    .Q_N(_12814_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][30]$_DFFE_PP_  (.CLK(clknet_leaf_772_clk),
    .RESET_B(net1260),
    .D(_01353_),
    .Q_N(_12813_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][31]$_DFFE_PP_  (.CLK(clknet_leaf_678_clk),
    .RESET_B(net1261),
    .D(_01354_),
    .Q_N(_12812_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][3]$_DFFE_PP_  (.CLK(clknet_8_46_0_clk),
    .RESET_B(net1262),
    .D(_01355_),
    .Q_N(_12811_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][4]$_DFFE_PP_  (.CLK(clknet_8_134_0_clk),
    .RESET_B(net1263),
    .D(_01356_),
    .Q_N(_12810_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_1135_clk),
    .RESET_B(net1264),
    .D(_01357_),
    .Q_N(_12809_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][6]$_DFFE_PP_  (.CLK(clknet_8_9_0_clk),
    .RESET_B(net1265),
    .D(_01358_),
    .Q_N(_12808_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1266),
    .D(_01359_),
    .Q_N(_12807_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_956_clk),
    .RESET_B(net1267),
    .D(_01360_),
    .Q_N(_12806_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1268),
    .D(_01361_),
    .Q_N(_12805_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[29][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_1043_clk),
    .RESET_B(net1269),
    .D(_01362_),
    .Q_N(_12804_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_1077_clk),
    .RESET_B(net1270),
    .D(_01363_),
    .Q_N(_12803_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_833_clk),
    .RESET_B(net1271),
    .D(_01364_),
    .Q_N(_12802_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1272),
    .D(_01365_),
    .Q_N(_12801_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_1027_clk),
    .RESET_B(net1273),
    .D(_01366_),
    .Q_N(_12800_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][14]$_DFFE_PP_  (.CLK(clknet_8_167_0_clk),
    .RESET_B(net1274),
    .D(_01367_),
    .Q_N(_12799_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_1144_clk),
    .RESET_B(net1275),
    .D(_01368_),
    .Q_N(_12798_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_1032_clk),
    .RESET_B(net1276),
    .D(_01369_),
    .Q_N(_12797_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_1026_clk),
    .RESET_B(net1277),
    .D(_01370_),
    .Q_N(_12796_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_1051_clk),
    .RESET_B(net1278),
    .D(_01371_),
    .Q_N(_12795_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_708_clk),
    .RESET_B(net1279),
    .D(_01372_),
    .Q_N(_12794_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1280),
    .D(_01373_),
    .Q_N(_12793_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_1066_clk),
    .RESET_B(net1281),
    .D(_01374_),
    .Q_N(_12792_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_1053_clk),
    .RESET_B(net1282),
    .D(_01375_),
    .Q_N(_12791_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][22]$_DFFE_PP_  (.CLK(clknet_8_170_0_clk),
    .RESET_B(net1283),
    .D(_01376_),
    .Q_N(_12790_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_836_clk),
    .RESET_B(net1284),
    .D(_01377_),
    .Q_N(_12789_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_824_clk),
    .RESET_B(net1285),
    .D(_01378_),
    .Q_N(_12788_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_792_clk),
    .RESET_B(net1286),
    .D(_01379_),
    .Q_N(_12787_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_724_clk),
    .RESET_B(net1287),
    .D(_01380_),
    .Q_N(_12786_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_808_clk),
    .RESET_B(net1288),
    .D(_01381_),
    .Q_N(_12785_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_711_clk),
    .RESET_B(net1289),
    .D(_01382_),
    .Q_N(_12784_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_811_clk),
    .RESET_B(net1290),
    .D(_01383_),
    .Q_N(_12783_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][2]$_DFFE_PP_  (.CLK(clknet_8_37_0_clk),
    .RESET_B(net1291),
    .D(_01384_),
    .Q_N(_12782_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_689_clk),
    .RESET_B(net1292),
    .D(_01385_),
    .Q_N(_12781_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_701_clk),
    .RESET_B(net1293),
    .D(_01386_),
    .Q_N(_12780_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_1086_clk),
    .RESET_B(net1294),
    .D(_01387_),
    .Q_N(_12779_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_1072_clk),
    .RESET_B(net1295),
    .D(_01388_),
    .Q_N(_12778_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_1092_clk),
    .RESET_B(net1296),
    .D(_01389_),
    .Q_N(_12777_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1297),
    .D(_01390_),
    .Q_N(_12776_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_1150_clk),
    .RESET_B(net1298),
    .D(_01391_),
    .Q_N(_12775_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_949_clk),
    .RESET_B(net1299),
    .D(_01392_),
    .Q_N(_12774_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][9]$_DFFE_PP_  (.CLK(clknet_8_52_0_clk),
    .RESET_B(net1300),
    .D(_01393_),
    .Q_N(_12773_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[2][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_998_clk),
    .RESET_B(net1301),
    .D(_01394_),
    .Q_N(_12772_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_1112_clk),
    .RESET_B(net1302),
    .D(_01395_),
    .Q_N(_12771_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_828_clk),
    .RESET_B(net1303),
    .D(_01396_),
    .Q_N(_12770_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][12]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1304),
    .D(_01397_),
    .Q_N(_12769_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][13]$_DFFE_PP_  (.CLK(clknet_leaf_1011_clk),
    .RESET_B(net1305),
    .D(_01398_),
    .Q_N(_12768_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][14]$_DFFE_PP_  (.CLK(clknet_leaf_678_clk),
    .RESET_B(net1306),
    .D(_01399_),
    .Q_N(_12767_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][15]$_DFFE_PP_  (.CLK(clknet_8_39_0_clk),
    .RESET_B(net1307),
    .D(_01400_),
    .Q_N(_12766_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][16]$_DFFE_PP_  (.CLK(clknet_leaf_1052_clk),
    .RESET_B(net1308),
    .D(_01401_),
    .Q_N(_12765_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][17]$_DFFE_PP_  (.CLK(clknet_8_61_0_clk),
    .RESET_B(net1309),
    .D(_01402_),
    .Q_N(_12764_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][18]$_DFFE_PP_  (.CLK(clknet_leaf_1048_clk),
    .RESET_B(net1310),
    .D(_01403_),
    .Q_N(_12763_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][19]$_DFFE_PP_  (.CLK(clknet_leaf_748_clk),
    .RESET_B(net1311),
    .D(_01404_),
    .Q_N(_12762_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1312),
    .D(_01405_),
    .Q_N(_12761_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][20]$_DFFE_PP_  (.CLK(clknet_8_137_0_clk),
    .RESET_B(net1313),
    .D(_01406_),
    .Q_N(_12760_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][21]$_DFFE_PP_  (.CLK(clknet_leaf_900_clk),
    .RESET_B(net1314),
    .D(_01407_),
    .Q_N(_12759_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][22]$_DFFE_PP_  (.CLK(clknet_8_139_0_clk),
    .RESET_B(net1315),
    .D(_01408_),
    .Q_N(_12758_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][23]$_DFFE_PP_  (.CLK(clknet_leaf_879_clk),
    .RESET_B(net1316),
    .D(_01409_),
    .Q_N(_12757_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][24]$_DFFE_PP_  (.CLK(clknet_leaf_861_clk),
    .RESET_B(net1317),
    .D(_01410_),
    .Q_N(_12756_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][25]$_DFFE_PP_  (.CLK(clknet_leaf_799_clk),
    .RESET_B(net1318),
    .D(_01411_),
    .Q_N(_12755_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][26]$_DFFE_PP_  (.CLK(clknet_8_234_0_clk),
    .RESET_B(net1319),
    .D(_01412_),
    .Q_N(_12754_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][27]$_DFFE_PP_  (.CLK(clknet_leaf_749_clk),
    .RESET_B(net1320),
    .D(_01413_),
    .Q_N(_12753_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][28]$_DFFE_PP_  (.CLK(clknet_8_235_0_clk),
    .RESET_B(net1321),
    .D(_01414_),
    .Q_N(_12752_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][29]$_DFFE_PP_  (.CLK(clknet_leaf_791_clk),
    .RESET_B(net1322),
    .D(_01415_),
    .Q_N(_12751_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][2]$_DFFE_PP_  (.CLK(clknet_8_36_0_clk),
    .RESET_B(net1323),
    .D(_01416_),
    .Q_N(_12750_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][30]$_DFFE_PP_  (.CLK(clknet_leaf_770_clk),
    .RESET_B(net1324),
    .D(_01417_),
    .Q_N(_12749_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][31]$_DFFE_PP_  (.CLK(clknet_leaf_678_clk),
    .RESET_B(net1325),
    .D(_01418_),
    .Q_N(_12748_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_1037_clk),
    .RESET_B(net1326),
    .D(_01419_),
    .Q_N(_12747_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_1069_clk),
    .RESET_B(net1327),
    .D(_01420_),
    .Q_N(_12746_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_1135_clk),
    .RESET_B(net1328),
    .D(_01421_),
    .Q_N(_12745_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1329),
    .D(_01422_),
    .Q_N(_12744_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1330),
    .D(_01423_),
    .Q_N(_12743_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_956_clk),
    .RESET_B(net1331),
    .D(_01424_),
    .Q_N(_12742_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1332),
    .D(_01425_),
    .Q_N(_12741_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[30][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_1000_clk),
    .RESET_B(net1333),
    .D(_01426_),
    .Q_N(_12740_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_1035_clk),
    .RESET_B(net1334),
    .D(_01427_),
    .Q_N(_12739_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_828_clk),
    .RESET_B(net1335),
    .D(_01428_),
    .Q_N(_12738_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][12]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1336),
    .D(_01429_),
    .Q_N(_12737_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][13]$_DFFE_PP_  (.CLK(clknet_8_148_0_clk),
    .RESET_B(net1337),
    .D(_01430_),
    .Q_N(_12736_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][14]$_DFFE_PP_  (.CLK(clknet_leaf_679_clk),
    .RESET_B(net1338),
    .D(_01431_),
    .Q_N(_12735_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][15]$_DFFE_PP_  (.CLK(clknet_leaf_1116_clk),
    .RESET_B(net1339),
    .D(_01432_),
    .Q_N(_12734_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][16]$_DFFE_PP_  (.CLK(clknet_leaf_1049_clk),
    .RESET_B(net1340),
    .D(_01433_),
    .Q_N(_12733_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][17]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1341),
    .D(_01434_),
    .Q_N(_12732_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][18]$_DFFE_PP_  (.CLK(clknet_leaf_1048_clk),
    .RESET_B(net1342),
    .D(_01435_),
    .Q_N(_12731_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][19]$_DFFE_PP_  (.CLK(clknet_leaf_748_clk),
    .RESET_B(net1343),
    .D(_01436_),
    .Q_N(_12730_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1344),
    .D(_01437_),
    .Q_N(_12729_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][20]$_DFFE_PP_  (.CLK(clknet_8_137_0_clk),
    .RESET_B(net1345),
    .D(_01438_),
    .Q_N(_12728_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][21]$_DFFE_PP_  (.CLK(clknet_8_140_0_clk),
    .RESET_B(net1346),
    .D(_01439_),
    .Q_N(_12727_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][22]$_DFFE_PP_  (.CLK(clknet_leaf_874_clk),
    .RESET_B(net1347),
    .D(_01440_),
    .Q_N(_12726_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][23]$_DFFE_PP_  (.CLK(clknet_leaf_878_clk),
    .RESET_B(net1348),
    .D(_01441_),
    .Q_N(_12725_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][24]$_DFFE_PP_  (.CLK(clknet_8_160_0_clk),
    .RESET_B(net1349),
    .D(_01442_),
    .Q_N(_12724_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][25]$_DFFE_PP_  (.CLK(clknet_leaf_758_clk),
    .RESET_B(net1350),
    .D(_01443_),
    .Q_N(_12723_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][26]$_DFFE_PP_  (.CLK(clknet_leaf_734_clk),
    .RESET_B(net1351),
    .D(_01444_),
    .Q_N(_12722_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][27]$_DFFE_PP_  (.CLK(clknet_leaf_752_clk),
    .RESET_B(net1352),
    .D(_01445_),
    .Q_N(_12721_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][28]$_DFFE_PP_  (.CLK(clknet_leaf_733_clk),
    .RESET_B(net1353),
    .D(_01446_),
    .Q_N(_12720_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][29]$_DFFE_PP_  (.CLK(clknet_8_171_0_clk),
    .RESET_B(net1354),
    .D(_01447_),
    .Q_N(_12719_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_1133_clk),
    .RESET_B(net1355),
    .D(_01448_),
    .Q_N(_12718_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][30]$_DFFE_PP_  (.CLK(clknet_leaf_692_clk),
    .RESET_B(net1356),
    .D(_01449_),
    .Q_N(_12717_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][31]$_DFFE_PP_  (.CLK(clknet_leaf_677_clk),
    .RESET_B(net1357),
    .D(_01450_),
    .Q_N(_12716_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_1057_clk),
    .RESET_B(net1358),
    .D(_01451_),
    .Q_N(_12715_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_1067_clk),
    .RESET_B(net1359),
    .D(_01452_),
    .Q_N(_12714_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_1135_clk),
    .RESET_B(net1360),
    .D(_01453_),
    .Q_N(_12713_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1361),
    .D(_01454_),
    .Q_N(_12712_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1362),
    .D(_01455_),
    .Q_N(_12711_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][8]$_DFFE_PP_  (.CLK(clknet_8_158_0_clk),
    .RESET_B(net1363),
    .D(_01456_),
    .Q_N(_12710_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1364),
    .D(_01457_),
    .Q_N(_12709_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[31][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][0]$_DFFE_PP_  (.CLK(clknet_8_147_0_clk),
    .RESET_B(net1365),
    .D(_01458_),
    .Q_N(_12708_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_1076_clk),
    .RESET_B(net1366),
    .D(_01459_),
    .Q_N(_12707_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_832_clk),
    .RESET_B(net1367),
    .D(_01460_),
    .Q_N(_12706_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1368),
    .D(_01461_),
    .Q_N(_12705_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_1020_clk),
    .RESET_B(net1369),
    .D(_01462_),
    .Q_N(_12704_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_937_clk),
    .RESET_B(net1370),
    .D(_01463_),
    .Q_N(_12703_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_1104_clk),
    .RESET_B(net1371),
    .D(_01464_),
    .Q_N(_12702_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_1033_clk),
    .RESET_B(net1372),
    .D(_01465_),
    .Q_N(_12701_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_1027_clk),
    .RESET_B(net1373),
    .D(_01466_),
    .Q_N(_12700_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][18]$_DFFE_PP_  (.CLK(clknet_8_152_0_clk),
    .RESET_B(net1374),
    .D(_01467_),
    .Q_N(_12699_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][19]$_DFFE_PP_  (.CLK(clknet_8_230_0_clk),
    .RESET_B(net1375),
    .D(_01468_),
    .Q_N(_12698_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][1]$_DFFE_PP_  (.CLK(clknet_8_59_0_clk),
    .RESET_B(net1376),
    .D(_01469_),
    .Q_N(_12697_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_1054_clk),
    .RESET_B(net1377),
    .D(_01470_),
    .Q_N(_12696_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_1052_clk),
    .RESET_B(net1378),
    .D(_01471_),
    .Q_N(_12695_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_824_clk),
    .RESET_B(net1379),
    .D(_01472_),
    .Q_N(_12694_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_845_clk),
    .RESET_B(net1380),
    .D(_01473_),
    .Q_N(_12693_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_824_clk),
    .RESET_B(net1381),
    .D(_01474_),
    .Q_N(_12692_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_815_clk),
    .RESET_B(net1382),
    .D(_01475_),
    .Q_N(_12691_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_725_clk),
    .RESET_B(net1383),
    .D(_01476_),
    .Q_N(_12690_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][27]$_DFFE_PP_  (.CLK(clknet_8_187_0_clk),
    .RESET_B(net1384),
    .D(_01477_),
    .Q_N(_12689_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_723_clk),
    .RESET_B(net1385),
    .D(_01478_),
    .Q_N(_12688_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_814_clk),
    .RESET_B(net1386),
    .D(_01479_),
    .Q_N(_12687_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_1120_clk),
    .RESET_B(net1387),
    .D(_01480_),
    .Q_N(_12686_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_690_clk),
    .RESET_B(net1388),
    .D(_01481_),
    .Q_N(_12685_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][31]$_DFFE_PP_  (.CLK(clknet_8_254_0_clk),
    .RESET_B(net1389),
    .D(_01482_),
    .Q_N(_12684_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_1086_clk),
    .RESET_B(net1390),
    .D(_01483_),
    .Q_N(_12683_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_1070_clk),
    .RESET_B(net1391),
    .D(_01484_),
    .Q_N(_12682_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][5]$_DFFE_PP_  (.CLK(clknet_8_40_0_clk),
    .RESET_B(net1392),
    .D(_01485_),
    .Q_N(_12681_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1393),
    .D(_01486_),
    .Q_N(_12680_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][7]$_DFFE_PP_  (.CLK(clknet_8_52_0_clk),
    .RESET_B(net1394),
    .D(_01487_),
    .Q_N(_12679_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_948_clk),
    .RESET_B(net1395),
    .D(_01488_),
    .Q_N(_12678_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1396),
    .D(_01489_),
    .Q_N(_12677_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[3][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_1047_clk),
    .RESET_B(net1397),
    .D(_01490_),
    .Q_N(_12676_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_1091_clk),
    .RESET_B(net1398),
    .D(_01491_),
    .Q_N(_12675_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_837_clk),
    .RESET_B(net1399),
    .D(_01492_),
    .Q_N(_12674_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1400),
    .D(_01493_),
    .Q_N(_12673_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_1017_clk),
    .RESET_B(net1401),
    .D(_01494_),
    .Q_N(_12672_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_938_clk),
    .RESET_B(net1402),
    .D(_01495_),
    .Q_N(_12671_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][15]$_DFFE_PP_  (.CLK(clknet_8_34_0_clk),
    .RESET_B(net1403),
    .D(_01496_),
    .Q_N(_12670_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_1028_clk),
    .RESET_B(net1404),
    .D(_01497_),
    .Q_N(_12669_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_1124_clk),
    .RESET_B(net1405),
    .D(_01498_),
    .Q_N(_12668_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_914_clk),
    .RESET_B(net1406),
    .D(_01499_),
    .Q_N(_12667_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_714_clk),
    .RESET_B(net1407),
    .D(_01500_),
    .Q_N(_12666_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1408),
    .D(_01501_),
    .Q_N(_12665_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_899_clk),
    .RESET_B(net1409),
    .D(_01502_),
    .Q_N(_12664_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_910_clk),
    .RESET_B(net1410),
    .D(_01503_),
    .Q_N(_12663_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][22]$_DFFE_PP_  (.CLK(clknet_8_169_0_clk),
    .RESET_B(net1411),
    .D(_01504_),
    .Q_N(_12662_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_933_clk),
    .RESET_B(net1412),
    .D(_01505_),
    .Q_N(_12661_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_859_clk),
    .RESET_B(net1413),
    .D(_01506_),
    .Q_N(_12660_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_795_clk),
    .RESET_B(net1414),
    .D(_01507_),
    .Q_N(_12659_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_768_clk),
    .RESET_B(net1415),
    .D(_01508_),
    .Q_N(_12658_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_801_clk),
    .RESET_B(net1416),
    .D(_01509_),
    .Q_N(_12657_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_712_clk),
    .RESET_B(net1417),
    .D(_01510_),
    .Q_N(_12656_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_794_clk),
    .RESET_B(net1418),
    .D(_01511_),
    .Q_N(_12655_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_1122_clk),
    .RESET_B(net1419),
    .D(_01512_),
    .Q_N(_12654_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_689_clk),
    .RESET_B(net1420),
    .D(_01513_),
    .Q_N(_12653_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_697_clk),
    .RESET_B(net1421),
    .D(_01514_),
    .Q_N(_12652_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_1088_clk),
    .RESET_B(net1422),
    .D(_01515_),
    .Q_N(_12651_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_1074_clk),
    .RESET_B(net1423),
    .D(_01516_),
    .Q_N(_12650_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_1096_clk),
    .RESET_B(net1424),
    .D(_01517_),
    .Q_N(_12649_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][6]$_DFFE_PP_  (.CLK(clknet_8_53_0_clk),
    .RESET_B(net1425),
    .D(_01518_),
    .Q_N(_12648_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1426),
    .D(_01519_),
    .Q_N(_12647_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_924_clk),
    .RESET_B(net1427),
    .D(_01520_),
    .Q_N(_12646_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1428),
    .D(_01521_),
    .Q_N(_12645_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[4][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_1046_clk),
    .RESET_B(net1429),
    .D(_01522_),
    .Q_N(_12644_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_1091_clk),
    .RESET_B(net1430),
    .D(_01523_),
    .Q_N(_12643_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_837_clk),
    .RESET_B(net1431),
    .D(_01524_),
    .Q_N(_12642_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][12]$_DFFE_PP_  (.CLK(clknet_8_8_0_clk),
    .RESET_B(net1432),
    .D(_01525_),
    .Q_N(_12641_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_1007_clk),
    .RESET_B(net1433),
    .D(_01526_),
    .Q_N(_12640_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_933_clk),
    .RESET_B(net1434),
    .D(_01527_),
    .Q_N(_12639_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_1087_clk),
    .RESET_B(net1435),
    .D(_01528_),
    .Q_N(_12638_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_1040_clk),
    .RESET_B(net1436),
    .D(_01529_),
    .Q_N(_12637_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_1125_clk),
    .RESET_B(net1437),
    .D(_01530_),
    .Q_N(_12636_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_914_clk),
    .RESET_B(net1438),
    .D(_01531_),
    .Q_N(_12635_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_714_clk),
    .RESET_B(net1439),
    .D(_01532_),
    .Q_N(_12634_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1440),
    .D(_01533_),
    .Q_N(_12633_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_899_clk),
    .RESET_B(net1441),
    .D(_01534_),
    .Q_N(_12632_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_910_clk),
    .RESET_B(net1442),
    .D(_01535_),
    .Q_N(_12631_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_857_clk),
    .RESET_B(net1443),
    .D(_01536_),
    .Q_N(_12630_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_850_clk),
    .RESET_B(net1444),
    .D(_01537_),
    .Q_N(_12629_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_857_clk),
    .RESET_B(net1445),
    .D(_01538_),
    .Q_N(_12628_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_793_clk),
    .RESET_B(net1446),
    .D(_01539_),
    .Q_N(_12627_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][26]$_DFFE_PP_  (.CLK(clknet_8_232_0_clk),
    .RESET_B(net1447),
    .D(_01540_),
    .Q_N(_12626_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_806_clk),
    .RESET_B(net1448),
    .D(_01541_),
    .Q_N(_12625_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][28]$_DFFE_PP_  (.CLK(clknet_8_227_0_clk),
    .RESET_B(net1449),
    .D(_01542_),
    .Q_N(_12624_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_794_clk),
    .RESET_B(net1450),
    .D(_01543_),
    .Q_N(_12623_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_1129_clk),
    .RESET_B(net1451),
    .D(_01544_),
    .Q_N(_12622_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_698_clk),
    .RESET_B(net1452),
    .D(_01545_),
    .Q_N(_12621_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_697_clk),
    .RESET_B(net1453),
    .D(_01546_),
    .Q_N(_12620_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_1088_clk),
    .RESET_B(net1454),
    .D(_01547_),
    .Q_N(_12619_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_1069_clk),
    .RESET_B(net1455),
    .D(_01548_),
    .Q_N(_12618_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_1096_clk),
    .RESET_B(net1456),
    .D(_01549_),
    .Q_N(_12617_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1457),
    .D(_01550_),
    .Q_N(_12616_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1458),
    .D(_01551_),
    .Q_N(_12615_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_934_clk),
    .RESET_B(net1459),
    .D(_01552_),
    .Q_N(_12614_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][9]$_DFFE_PP_  (.CLK(clknet_8_53_0_clk),
    .RESET_B(net1460),
    .D(_01553_),
    .Q_N(_12613_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[5][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_1047_clk),
    .RESET_B(net1461),
    .D(_01554_),
    .Q_N(_12612_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_1090_clk),
    .RESET_B(net1462),
    .D(_01555_),
    .Q_N(_12611_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_836_clk),
    .RESET_B(net1463),
    .D(_01556_),
    .Q_N(_12610_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1464),
    .D(_01557_),
    .Q_N(_12609_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_1006_clk),
    .RESET_B(net1465),
    .D(_01558_),
    .Q_N(_12608_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_938_clk),
    .RESET_B(net1466),
    .D(_01559_),
    .Q_N(_12607_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_1087_clk),
    .RESET_B(net1467),
    .D(_01560_),
    .Q_N(_12606_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_1041_clk),
    .RESET_B(net1468),
    .D(_01561_),
    .Q_N(_12605_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_1125_clk),
    .RESET_B(net1469),
    .D(_01562_),
    .Q_N(_12604_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_912_clk),
    .RESET_B(net1470),
    .D(_01563_),
    .Q_N(_12603_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_707_clk),
    .RESET_B(net1471),
    .D(_01564_),
    .Q_N(_12602_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1472),
    .D(_01565_),
    .Q_N(_12601_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_900_clk),
    .RESET_B(net1473),
    .D(_01566_),
    .Q_N(_12600_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_912_clk),
    .RESET_B(net1474),
    .D(_01567_),
    .Q_N(_12599_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_858_clk),
    .RESET_B(net1475),
    .D(_01568_),
    .Q_N(_12598_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][23]$_DFFE_PP_  (.CLK(clknet_8_163_0_clk),
    .RESET_B(net1476),
    .D(_01569_),
    .Q_N(_12597_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_858_clk),
    .RESET_B(net1477),
    .D(_01570_),
    .Q_N(_12596_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_795_clk),
    .RESET_B(net1478),
    .D(_01571_),
    .Q_N(_12595_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_768_clk),
    .RESET_B(net1479),
    .D(_01572_),
    .Q_N(_12594_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_806_clk),
    .RESET_B(net1480),
    .D(_01573_),
    .Q_N(_12593_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_712_clk),
    .RESET_B(net1481),
    .D(_01574_),
    .Q_N(_12592_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_806_clk),
    .RESET_B(net1482),
    .D(_01575_),
    .Q_N(_12591_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_1128_clk),
    .RESET_B(net1483),
    .D(_01576_),
    .Q_N(_12590_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_690_clk),
    .RESET_B(net1484),
    .D(_01577_),
    .Q_N(_12589_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_697_clk),
    .RESET_B(net1485),
    .D(_01578_),
    .Q_N(_12588_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_1089_clk),
    .RESET_B(net1486),
    .D(_01579_),
    .Q_N(_12587_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_1074_clk),
    .RESET_B(net1487),
    .D(_01580_),
    .Q_N(_12586_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_1092_clk),
    .RESET_B(net1488),
    .D(_01581_),
    .Q_N(_12585_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1489),
    .D(_01582_),
    .Q_N(_12584_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1490),
    .D(_01583_),
    .Q_N(_12583_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_935_clk),
    .RESET_B(net1491),
    .D(_01584_),
    .Q_N(_12582_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1492),
    .D(_01585_),
    .Q_N(_12581_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[6][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_1046_clk),
    .RESET_B(net1493),
    .D(_01586_),
    .Q_N(_12580_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_1079_clk),
    .RESET_B(net1494),
    .D(_01587_),
    .Q_N(_12579_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][11]$_DFFE_PP_  (.CLK(clknet_8_176_0_clk),
    .RESET_B(net1495),
    .D(_01588_),
    .Q_N(_12578_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1496),
    .D(_01589_),
    .Q_N(_12577_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_1006_clk),
    .RESET_B(net1497),
    .D(_01590_),
    .Q_N(_12576_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][14]$_DFFE_PP_  (.CLK(clknet_8_166_0_clk),
    .RESET_B(net1498),
    .D(_01591_),
    .Q_N(_12575_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][15]$_DFFE_PP_  (.CLK(clknet_8_34_0_clk),
    .RESET_B(net1499),
    .D(_01592_),
    .Q_N(_12574_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][16]$_DFFE_PP_  (.CLK(clknet_8_47_0_clk),
    .RESET_B(net1500),
    .D(_01593_),
    .Q_N(_12573_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_1026_clk),
    .RESET_B(net1501),
    .D(_01594_),
    .Q_N(_12572_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][18]$_DFFE_PP_  (.CLK(clknet_8_152_0_clk),
    .RESET_B(net1502),
    .D(_01595_),
    .Q_N(_12571_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][19]$_DFFE_PP_  (.CLK(clknet_8_230_0_clk),
    .RESET_B(net1503),
    .D(_01596_),
    .Q_N(_12570_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1504),
    .D(_01597_),
    .Q_N(_12569_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_909_clk),
    .RESET_B(net1505),
    .D(_01598_),
    .Q_N(_12568_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][21]$_DFFE_PP_  (.CLK(clknet_8_141_0_clk),
    .RESET_B(net1506),
    .D(_01599_),
    .Q_N(_12567_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_859_clk),
    .RESET_B(net1507),
    .D(_01600_),
    .Q_N(_12566_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][23]$_DFFE_PP_  (.CLK(clknet_8_166_0_clk),
    .RESET_B(net1508),
    .D(_01601_),
    .Q_N(_12565_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_823_clk),
    .RESET_B(net1509),
    .D(_01602_),
    .Q_N(_12564_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_793_clk),
    .RESET_B(net1510),
    .D(_01603_),
    .Q_N(_12563_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_694_clk),
    .RESET_B(net1511),
    .D(_01604_),
    .Q_N(_12562_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][27]$_DFFE_PP_  (.CLK(clknet_8_185_0_clk),
    .RESET_B(net1512),
    .D(_01605_),
    .Q_N(_12561_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_722_clk),
    .RESET_B(net1513),
    .D(_01606_),
    .Q_N(_12560_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_807_clk),
    .RESET_B(net1514),
    .D(_01607_),
    .Q_N(_12559_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_1126_clk),
    .RESET_B(net1515),
    .D(_01608_),
    .Q_N(_12558_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_696_clk),
    .RESET_B(net1516),
    .D(_01609_),
    .Q_N(_12557_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_698_clk),
    .RESET_B(net1517),
    .D(_01610_),
    .Q_N(_12556_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_1089_clk),
    .RESET_B(net1518),
    .D(_01611_),
    .Q_N(_12555_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_1070_clk),
    .RESET_B(net1519),
    .D(_01612_),
    .Q_N(_12554_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_1093_clk),
    .RESET_B(net1520),
    .D(_01613_),
    .Q_N(_12553_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1521),
    .D(_01614_),
    .Q_N(_12552_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][7]$_DFFE_PP_  (.CLK(clknet_8_0_0_clk),
    .RESET_B(net1522),
    .D(_01615_),
    .Q_N(_12551_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_935_clk),
    .RESET_B(net1523),
    .D(_01616_),
    .Q_N(_12550_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1524),
    .D(_01617_),
    .Q_N(_12549_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[7][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_997_clk),
    .RESET_B(net1525),
    .D(_01618_),
    .Q_N(_12548_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_1106_clk),
    .RESET_B(net1526),
    .D(_01619_),
    .Q_N(_12547_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_780_clk),
    .RESET_B(net1527),
    .D(_01620_),
    .Q_N(_12546_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][12]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1528),
    .D(_01621_),
    .Q_N(_12545_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][13]$_DFFE_PP_  (.CLK(clknet_8_63_0_clk),
    .RESET_B(net1529),
    .D(_01622_),
    .Q_N(_12544_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][14]$_DFFE_PP_  (.CLK(clknet_leaf_948_clk),
    .RESET_B(net1530),
    .D(_01623_),
    .Q_N(_12543_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][15]$_DFFE_PP_  (.CLK(clknet_8_36_0_clk),
    .RESET_B(net1531),
    .D(_01624_),
    .Q_N(_12542_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][16]$_DFFE_PP_  (.CLK(clknet_8_44_0_clk),
    .RESET_B(net1532),
    .D(_01625_),
    .Q_N(_12541_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][17]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1533),
    .D(_01626_),
    .Q_N(_12540_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][18]$_DFFE_PP_  (.CLK(clknet_leaf_920_clk),
    .RESET_B(net1534),
    .D(_01627_),
    .Q_N(_12539_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][19]$_DFFE_PP_  (.CLK(clknet_leaf_765_clk),
    .RESET_B(net1535),
    .D(_01628_),
    .Q_N(_12538_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][1]$_DFFE_PP_  (.CLK(clknet_8_10_0_clk),
    .RESET_B(net1536),
    .D(_01629_),
    .Q_N(_12537_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][20]$_DFFE_PP_  (.CLK(clknet_leaf_886_clk),
    .RESET_B(net1537),
    .D(_01630_),
    .Q_N(_12536_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][21]$_DFFE_PP_  (.CLK(clknet_leaf_890_clk),
    .RESET_B(net1538),
    .D(_01631_),
    .Q_N(_12535_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][22]$_DFFE_PP_  (.CLK(clknet_leaf_852_clk),
    .RESET_B(net1539),
    .D(_01632_),
    .Q_N(_12534_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][23]$_DFFE_PP_  (.CLK(clknet_leaf_904_clk),
    .RESET_B(net1540),
    .D(_01633_),
    .Q_N(_12533_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][24]$_DFFE_PP_  (.CLK(clknet_leaf_853_clk),
    .RESET_B(net1541),
    .D(_01634_),
    .Q_N(_12532_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][25]$_DFFE_PP_  (.CLK(clknet_leaf_773_clk),
    .RESET_B(net1542),
    .D(_01635_),
    .Q_N(_12531_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][26]$_DFFE_PP_  (.CLK(clknet_leaf_739_clk),
    .RESET_B(net1543),
    .D(_01636_),
    .Q_N(_12530_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][27]$_DFFE_PP_  (.CLK(clknet_leaf_758_clk),
    .RESET_B(net1544),
    .D(_01637_),
    .Q_N(_12529_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][28]$_DFFE_PP_  (.CLK(clknet_leaf_740_clk),
    .RESET_B(net1545),
    .D(_01638_),
    .Q_N(_12528_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][29]$_DFFE_PP_  (.CLK(clknet_leaf_787_clk),
    .RESET_B(net1546),
    .D(_01639_),
    .Q_N(_12527_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_1134_clk),
    .RESET_B(net1547),
    .D(_01640_),
    .Q_N(_12526_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][30]$_DFFE_PP_  (.CLK(clknet_leaf_778_clk),
    .RESET_B(net1548),
    .D(_01641_),
    .Q_N(_12525_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][31]$_DFFE_PP_  (.CLK(clknet_leaf_780_clk),
    .RESET_B(net1549),
    .D(_01642_),
    .Q_N(_12524_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][3]$_DFFE_PP_  (.CLK(clknet_8_38_0_clk),
    .RESET_B(net1550),
    .D(_01643_),
    .Q_N(_12523_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_1069_clk),
    .RESET_B(net1551),
    .D(_01644_),
    .Q_N(_12522_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1552),
    .D(_01645_),
    .Q_N(_12521_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1553),
    .D(_01646_),
    .Q_N(_12520_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1554),
    .D(_01647_),
    .Q_N(_12519_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_961_clk),
    .RESET_B(net1555),
    .D(_01648_),
    .Q_N(_12518_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1556),
    .D(_01649_),
    .Q_N(_12517_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[8][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_999_clk),
    .RESET_B(net1557),
    .D(_01650_),
    .Q_N(_12516_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_1106_clk),
    .RESET_B(net1558),
    .D(_01651_),
    .Q_N(_12515_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_778_clk),
    .RESET_B(net1559),
    .D(_01652_),
    .Q_N(_12514_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][12]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1560),
    .D(_01653_),
    .Q_N(_12513_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][13]$_DFFE_PP_  (.CLK(clknet_leaf_1017_clk),
    .RESET_B(net1561),
    .D(_01654_),
    .Q_N(_12512_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][14]$_DFFE_PP_  (.CLK(clknet_8_165_0_clk),
    .RESET_B(net1562),
    .D(_01655_),
    .Q_N(_12511_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][15]$_DFFE_PP_  (.CLK(clknet_leaf_1104_clk),
    .RESET_B(net1563),
    .D(_01656_),
    .Q_N(_12510_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][16]$_DFFE_PP_  (.CLK(clknet_leaf_1122_clk),
    .RESET_B(net1564),
    .D(_01657_),
    .Q_N(_12509_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][17]$_DFFE_PP_  (.CLK(clknet_leaf_1126_clk),
    .RESET_B(net1565),
    .D(_01658_),
    .Q_N(_12508_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][18]$_DFFE_PP_  (.CLK(clknet_leaf_920_clk),
    .RESET_B(net1566),
    .D(_01659_),
    .Q_N(_12507_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][19]$_DFFE_PP_  (.CLK(clknet_leaf_743_clk),
    .RESET_B(net1567),
    .D(_01660_),
    .Q_N(_12506_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1568),
    .D(_01661_),
    .Q_N(_12505_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][20]$_DFFE_PP_  (.CLK(clknet_leaf_883_clk),
    .RESET_B(net1569),
    .D(_01662_),
    .Q_N(_12504_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][21]$_DFFE_PP_  (.CLK(clknet_leaf_894_clk),
    .RESET_B(net1570),
    .D(_01663_),
    .Q_N(_12503_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][22]$_DFFE_PP_  (.CLK(clknet_leaf_877_clk),
    .RESET_B(net1571),
    .D(_01664_),
    .Q_N(_12502_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][23]$_DFFE_PP_  (.CLK(clknet_leaf_904_clk),
    .RESET_B(net1572),
    .D(_01665_),
    .Q_N(_12501_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][24]$_DFFE_PP_  (.CLK(clknet_leaf_854_clk),
    .RESET_B(net1573),
    .D(_01666_),
    .Q_N(_12500_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][25]$_DFFE_PP_  (.CLK(clknet_leaf_773_clk),
    .RESET_B(net1574),
    .D(_01667_),
    .Q_N(_12499_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][26]$_DFFE_PP_  (.CLK(clknet_leaf_739_clk),
    .RESET_B(net1575),
    .D(_01668_),
    .Q_N(_12498_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][27]$_DFFE_PP_  (.CLK(clknet_leaf_757_clk),
    .RESET_B(net1576),
    .D(_01669_),
    .Q_N(_12497_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][28]$_DFFE_PP_  (.CLK(clknet_leaf_740_clk),
    .RESET_B(net1577),
    .D(_01670_),
    .Q_N(_12496_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][29]$_DFFE_PP_  (.CLK(clknet_leaf_786_clk),
    .RESET_B(net1578),
    .D(_01671_),
    .Q_N(_12495_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_1129_clk),
    .RESET_B(net1579),
    .D(_01672_),
    .Q_N(_12494_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][30]$_DFFE_PP_  (.CLK(clknet_leaf_684_clk),
    .RESET_B(net1580),
    .D(_01673_),
    .Q_N(_12493_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][31]$_DFFE_PP_  (.CLK(clknet_leaf_682_clk),
    .RESET_B(net1581),
    .D(_01674_),
    .Q_N(_12492_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_1101_clk),
    .RESET_B(net1582),
    .D(_01675_),
    .Q_N(_12491_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_892_clk),
    .RESET_B(net1583),
    .D(_01676_),
    .Q_N(_12490_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_1134_clk),
    .RESET_B(net1584),
    .D(_01677_),
    .Q_N(_12489_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1585),
    .D(_01678_),
    .Q_N(_12488_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1586),
    .D(_01679_),
    .Q_N(_12487_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_960_clk),
    .RESET_B(net1587),
    .D(_01680_),
    .Q_N(_12486_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1588),
    .D(_01681_),
    .Q_N(_12485_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.cpuregs[9][9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_437_clk),
    .RESET_B(net1589),
    .D(_01682_),
    .Q_N(_00054_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[10]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_457_clk),
    .RESET_B(net1590),
    .D(_01683_),
    .Q_N(_12484_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[11]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_455_clk),
    .RESET_B(net1591),
    .D(_01684_),
    .Q_N(_12483_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[12]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_456_clk),
    .RESET_B(net1592),
    .D(_01685_),
    .Q_N(_12482_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[13]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_657_clk),
    .RESET_B(net1593),
    .D(_01686_),
    .Q_N(_12481_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[14]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_656_clk),
    .RESET_B(net1594),
    .D(_01687_),
    .Q_N(_12480_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[15]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_652_clk),
    .RESET_B(net1595),
    .D(_01688_),
    .Q_N(_12479_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[16]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_645_clk),
    .RESET_B(net1596),
    .D(_01689_),
    .Q_N(_12478_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[17]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_644_clk),
    .RESET_B(net1597),
    .D(_01690_),
    .Q_N(_12477_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[18]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_644_clk),
    .RESET_B(net1598),
    .D(_01691_),
    .Q_N(_12476_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[19]$_SDFFCE_PN0P_  (.CLK(clknet_8_198_0_clk),
    .RESET_B(net1599),
    .D(_01692_),
    .Q_N(_12475_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_452_clk),
    .RESET_B(net1600),
    .D(_01693_),
    .Q_N(_12474_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[20]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_646_clk),
    .RESET_B(net1601),
    .D(_01694_),
    .Q_N(_12473_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[21]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_647_clk),
    .RESET_B(net1602),
    .D(_01695_),
    .Q_N(_12472_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[22]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_646_clk),
    .RESET_B(net1603),
    .D(_01696_),
    .Q_N(_12471_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[23]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_645_clk),
    .RESET_B(net1604),
    .D(_01697_),
    .Q_N(_12470_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[24]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_645_clk),
    .RESET_B(net1605),
    .D(_01698_),
    .Q_N(_12469_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[25]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_647_clk),
    .RESET_B(net1606),
    .D(_01699_),
    .Q_N(_12468_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[26]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_647_clk),
    .RESET_B(net1607),
    .D(_01700_),
    .Q_N(_12467_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[27]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_636_clk),
    .RESET_B(net1608),
    .D(_01701_),
    .Q_N(_12466_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[28]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_636_clk),
    .RESET_B(net1609),
    .D(_01702_),
    .Q_N(_12465_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[29]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_640_clk),
    .RESET_B(net1610),
    .D(_01703_),
    .Q_N(_12464_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_450_clk),
    .RESET_B(net1611),
    .D(_01704_),
    .Q_N(_12463_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[30]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_636_clk),
    .RESET_B(net1612),
    .D(_01705_),
    .Q_N(_12462_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[31]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_640_clk),
    .RESET_B(net1613),
    .D(_01706_),
    .Q_N(_12461_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_450_clk),
    .RESET_B(net1614),
    .D(_01707_),
    .Q_N(_12460_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[4]$_SDFFCE_PN0P_  (.CLK(clknet_8_31_0_clk),
    .RESET_B(net1615),
    .D(_01708_),
    .Q_N(_12459_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[5]$_SDFFCE_PN0P_  (.CLK(clknet_8_241_0_clk),
    .RESET_B(net1616),
    .D(_01709_),
    .Q_N(_12458_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1617),
    .D(_01710_),
    .Q_N(_12457_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[7]$_SDFFCE_PN0P_  (.CLK(clknet_8_31_0_clk),
    .RESET_B(net1618),
    .D(_01711_),
    .Q_N(_12456_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[8]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_453_clk),
    .RESET_B(net1619),
    .D(_01712_),
    .Q_N(_12455_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm[9]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_453_clk),
    .RESET_B(net1620),
    .D(_01713_),
    .Q_N(_12454_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[10]$_DFFE_PN_  (.CLK(clknet_8_106_0_clk),
    .RESET_B(net1621),
    .D(_01714_),
    .Q_N(_12453_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11]$_DFFE_PN_  (.CLK(clknet_leaf_969_clk),
    .RESET_B(net1622),
    .D(_00033_),
    .Q_N(_12452_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12]$_DFFE_PN_  (.CLK(clknet_leaf_526_clk),
    .RESET_B(net1623),
    .D(_01715_),
    .Q_N(_12451_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[13]$_DFFE_PN_  (.CLK(clknet_leaf_467_clk),
    .RESET_B(net1624),
    .D(_01716_),
    .Q_N(_12450_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[14]$_DFFE_PN_  (.CLK(clknet_leaf_464_clk),
    .RESET_B(net1625),
    .D(_01717_),
    .Q_N(_12449_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15]$_DFFE_PN_  (.CLK(clknet_leaf_650_clk),
    .RESET_B(net1626),
    .D(_00038_),
    .Q_N(_12448_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[16]$_DFFE_PN_  (.CLK(clknet_8_194_0_clk),
    .RESET_B(net1627),
    .D(_00039_),
    .Q_N(_12447_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17]$_DFFE_PN_  (.CLK(clknet_leaf_634_clk),
    .RESET_B(net1628),
    .D(_00040_),
    .Q_N(_12446_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18]$_DFFE_PN_  (.CLK(clknet_leaf_648_clk),
    .RESET_B(net1629),
    .D(_00041_),
    .Q_N(_12445_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[19]$_DFFE_PN_  (.CLK(clknet_8_198_0_clk),
    .RESET_B(net1630),
    .D(_00042_),
    .Q_N(_00132_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1]$_DFFE_PN_  (.CLK(clknet_leaf_968_clk),
    .RESET_B(net1631),
    .D(_00034_),
    .Q_N(_12444_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20]$_DFFE_PN_  (.CLK(clknet_8_200_0_clk),
    .RESET_B(net1632),
    .D(_01718_),
    .Q_N(_00133_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2]$_DFFE_PN_  (.CLK(clknet_leaf_990_clk),
    .RESET_B(net1633),
    .D(_00035_),
    .Q_N(_12443_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3]$_DFFE_PN_  (.CLK(clknet_8_240_0_clk),
    .RESET_B(net1634),
    .D(_00036_),
    .Q_N(_12442_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[4]$_DFFE_PN_  (.CLK(clknet_leaf_991_clk),
    .RESET_B(net1635),
    .D(_00037_),
    .Q_N(_00131_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[5]$_DFFE_PN_  (.CLK(clknet_leaf_439_clk),
    .RESET_B(net1636),
    .D(_01719_),
    .Q_N(_12441_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[6]$_DFFE_PN_  (.CLK(clknet_leaf_439_clk),
    .RESET_B(net1637),
    .D(_01720_),
    .Q_N(_12440_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[7]$_DFFE_PN_  (.CLK(clknet_leaf_447_clk),
    .RESET_B(net1638),
    .D(_01721_),
    .Q_N(_12439_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[8]$_DFFE_PN_  (.CLK(clknet_leaf_447_clk),
    .RESET_B(net1639),
    .D(_01722_),
    .Q_N(_12438_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[9]$_DFFE_PN_  (.CLK(clknet_8_106_0_clk),
    .RESET_B(net1640),
    .D(_01723_),
    .Q_N(_12437_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_rd[0]$_DFFE_PN_  (.CLK(clknet_8_192_0_clk),
    .RESET_B(net1641),
    .D(_01724_),
    .Q_N(_12436_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_rd[1]$_DFFE_PN_  (.CLK(clknet_leaf_994_clk),
    .RESET_B(net1642),
    .D(_01725_),
    .Q_N(_12435_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_rd[2]$_DFFE_PN_  (.CLK(clknet_8_150_0_clk),
    .RESET_B(net1643),
    .D(_01726_),
    .Q_N(_12434_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_rd[3]$_DFFE_PN_  (.CLK(clknet_leaf_994_clk),
    .RESET_B(net1644),
    .D(_01727_),
    .Q_N(_12433_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoded_rd[4]$_DFFE_PN_  (.CLK(clknet_leaf_995_clk),
    .RESET_B(net1645),
    .D(_01728_),
    .Q_N(_12432_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoded_rd[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoder_pseudo_trigger$_SDFF_PN0_  (.CLK(clknet_8_193_0_clk),
    .RESET_B(net1646),
    .D(_01729_),
    .Q_N(_14057_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoder_pseudo_trigger ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.decoder_trigger$_DFF_P_  (.CLK(clknet_leaf_481_clk),
    .RESET_B(net1647),
    .D(_00044_),
    .Q_N(_00107_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.decoder_trigger ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_add$_SDFFE_PN0P_  (.CLK(clknet_leaf_502_clk),
    .RESET_B(net1648),
    .D(_01730_),
    .Q_N(_12431_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_add ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_addi$_SDFFE_PN0P_  (.CLK(clknet_leaf_505_clk),
    .RESET_B(net1649),
    .D(_01731_),
    .Q_N(_12430_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_addi ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_and$_SDFFE_PN0P_  (.CLK(clknet_leaf_490_clk),
    .RESET_B(net1650),
    .D(_01732_),
    .Q_N(_12429_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_and ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_andi$_SDFFE_PN0P_  (.CLK(clknet_leaf_491_clk),
    .RESET_B(net1651),
    .D(_01733_),
    .Q_N(_12428_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_andi ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_auipc$_DFFE_PN_  (.CLK(clknet_leaf_519_clk),
    .RESET_B(net1652),
    .D(_01734_),
    .Q_N(_12427_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_auipc ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_beq$_SDFFE_PN0P_  (.CLK(clknet_8_216_0_clk),
    .RESET_B(net1653),
    .D(_01735_),
    .Q_N(_12426_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_beq ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_bge$_SDFFE_PN0P_  (.CLK(clknet_8_198_0_clk),
    .RESET_B(net1654),
    .D(_01736_),
    .Q_N(_12425_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_bge ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_bgeu$_SDFFE_PN0P_  (.CLK(clknet_leaf_486_clk),
    .RESET_B(net1655),
    .D(_01737_),
    .Q_N(_12424_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_bgeu ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_blt$_SDFFE_PN0P_  (.CLK(clknet_leaf_501_clk),
    .RESET_B(net1656),
    .D(_01738_),
    .Q_N(_12423_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_blt ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_bltu$_SDFFE_PN0P_  (.CLK(clknet_8_199_0_clk),
    .RESET_B(net1657),
    .D(_01739_),
    .Q_N(_12422_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_bltu ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_bne$_SDFFE_PN0P_  (.CLK(clknet_leaf_491_clk),
    .RESET_B(net1658),
    .D(_01740_),
    .Q_N(_12421_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_bne ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_fence$_SDFFE_PN0P_  (.CLK(clknet_8_210_0_clk),
    .RESET_B(net1659),
    .D(_01741_),
    .Q_N(_12420_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_fence ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_jal$_DFFE_PN_  (.CLK(clknet_leaf_465_clk),
    .RESET_B(net1660),
    .D(_01742_),
    .Q_N(_00108_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_jal ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_jalr$_DFFE_PN_  (.CLK(clknet_leaf_518_clk),
    .RESET_B(net1661),
    .D(_01743_),
    .Q_N(_00051_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_jalr ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_lb$_DFFE_PP_  (.CLK(clknet_leaf_477_clk),
    .RESET_B(net1662),
    .D(_01744_),
    .Q_N(_12419_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_lb ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_lbu$_DFFE_PP_  (.CLK(clknet_8_210_0_clk),
    .RESET_B(net1663),
    .D(_01745_),
    .Q_N(_12418_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_lbu ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_lh$_DFFE_PP_  (.CLK(clknet_8_210_0_clk),
    .RESET_B(net1664),
    .D(_01746_),
    .Q_N(_12417_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_lh ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_lhu$_DFFE_PP_  (.CLK(clknet_leaf_478_clk),
    .RESET_B(net1665),
    .D(_01747_),
    .Q_N(_12416_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_lhu ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_lui$_DFFE_PN_  (.CLK(clknet_leaf_512_clk),
    .RESET_B(net1666),
    .D(_01748_),
    .Q_N(_12415_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_lui ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_lw$_DFFE_PP_  (.CLK(clknet_leaf_478_clk),
    .RESET_B(net1667),
    .D(_01749_),
    .Q_N(_12414_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_lw ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_or$_SDFFE_PN0P_  (.CLK(clknet_8_216_0_clk),
    .RESET_B(net1668),
    .D(_01750_),
    .Q_N(_12413_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_or ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_ori$_SDFFE_PN0P_  (.CLK(clknet_leaf_498_clk),
    .RESET_B(net1669),
    .D(_01751_),
    .Q_N(_12412_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_ori ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_rdcycle$_DFFE_PP_  (.CLK(clknet_leaf_485_clk),
    .RESET_B(net1670),
    .D(_01752_),
    .Q_N(_12411_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycle ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_rdcycleh$_DFFE_PP_  (.CLK(clknet_leaf_497_clk),
    .RESET_B(net1671),
    .D(_01753_),
    .Q_N(_12410_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_rdcycleh ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_rdinstr$_DFFE_PP_  (.CLK(clknet_leaf_497_clk),
    .RESET_B(net1672),
    .D(_01754_),
    .Q_N(_12409_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstr ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh$_DFFE_PP_  (.CLK(clknet_leaf_495_clk),
    .RESET_B(net1673),
    .D(_01755_),
    .Q_N(_12408_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_sb$_DFFE_PP_  (.CLK(clknet_leaf_517_clk),
    .RESET_B(net1674),
    .D(_01756_),
    .Q_N(_12407_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_sb ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_sh$_DFFE_PP_  (.CLK(clknet_leaf_477_clk),
    .RESET_B(net1675),
    .D(_01757_),
    .Q_N(_12406_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_sh ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_sll$_SDFFE_PN0P_  (.CLK(clknet_leaf_490_clk),
    .RESET_B(net1676),
    .D(_01758_),
    .Q_N(_12405_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_sll ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_slli$_DFFE_PP_  (.CLK(clknet_leaf_487_clk),
    .RESET_B(net1677),
    .D(_01759_),
    .Q_N(_12404_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_slli ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_slt$_SDFFE_PN0P_  (.CLK(clknet_leaf_496_clk),
    .RESET_B(net1678),
    .D(_01760_),
    .Q_N(_12403_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_slt ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_slti$_SDFFE_PN0P_  (.CLK(clknet_leaf_496_clk),
    .RESET_B(net1679),
    .D(_01761_),
    .Q_N(_12402_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_slti ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_sltiu$_SDFFE_PN0P_  (.CLK(clknet_leaf_490_clk),
    .RESET_B(net1680),
    .D(_01762_),
    .Q_N(_12401_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_sltiu ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_sltu$_SDFFE_PN0P_  (.CLK(clknet_leaf_493_clk),
    .RESET_B(net1681),
    .D(_01763_),
    .Q_N(_12400_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_sltu ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_sra$_SDFFE_PN0P_  (.CLK(clknet_leaf_489_clk),
    .RESET_B(net1682),
    .D(_01764_),
    .Q_N(_12399_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_sra ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_srai$_DFFE_PP_  (.CLK(clknet_leaf_489_clk),
    .RESET_B(net1683),
    .D(_01765_),
    .Q_N(_12398_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_srai ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_srl$_SDFFE_PN0P_  (.CLK(clknet_leaf_492_clk),
    .RESET_B(net1684),
    .D(_01766_),
    .Q_N(_12397_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_srl ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_srli$_DFFE_PP_  (.CLK(clknet_leaf_492_clk),
    .RESET_B(net1685),
    .D(_01767_),
    .Q_N(_12396_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_srli ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_sub$_SDFFE_PN0P_  (.CLK(clknet_leaf_502_clk),
    .RESET_B(net1686),
    .D(_01768_),
    .Q_N(_12395_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_sub ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_sw$_DFFE_PP_  (.CLK(clknet_leaf_478_clk),
    .RESET_B(net1687),
    .D(_01769_),
    .Q_N(_12394_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_sw ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_xor$_SDFFE_PN0P_  (.CLK(clknet_leaf_487_clk),
    .RESET_B(net1688),
    .D(_01770_),
    .Q_N(_12393_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_xor ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.instr_xori$_SDFFE_PN0P_  (.CLK(clknet_leaf_501_clk),
    .RESET_B(net1689),
    .D(_01771_),
    .Q_N(_12392_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.instr_xori ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_alu_reg_imm$_DFFE_PN_  (.CLK(clknet_8_211_0_clk),
    .RESET_B(net1690),
    .D(_01772_),
    .Q_N(_00122_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_alu_reg_imm ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_alu_reg_reg$_DFFE_PN_  (.CLK(clknet_leaf_513_clk),
    .RESET_B(net1691),
    .D(_01773_),
    .Q_N(_00123_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_alu_reg_reg ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_beq_bne_blt_bge_bltu_bgeu$_SDFFE_PN0N_  (.CLK(clknet_8_208_0_clk),
    .RESET_B(net1692),
    .D(_01774_),
    .Q_N(_00102_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_beq_bne_blt_bge_bltu_bgeu ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_compare$_SDFF_PP0_  (.CLK(clknet_leaf_485_clk),
    .RESET_B(net1693),
    .D(_01775_),
    .Q_N(_00138_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_compare ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_jalr_addi_slti_sltiu_xori_ori_andi$_DFFE_PP_  (.CLK(clknet_leaf_488_clk),
    .RESET_B(net1694),
    .D(_01776_),
    .Q_N(_12391_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_jalr_addi_slti_sltiu_xori_ori_andi ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_lb_lh_lw_lbu_lhu$_DFFE_PN_  (.CLK(clknet_leaf_517_clk),
    .RESET_B(net1695),
    .D(_01777_),
    .Q_N(_00101_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_lb_lh_lw_lbu_lhu ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_lui_auipc_jal$_DFF_P_  (.CLK(clknet_leaf_482_clk),
    .RESET_B(net1696),
    .D(_00045_),
    .Q_N(_12390_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_lui_auipc_jal ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_sb_sh_sw$_DFFE_PN_  (.CLK(clknet_leaf_512_clk),
    .RESET_B(net1697),
    .D(_01778_),
    .Q_N(_12389_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_sb_sh_sw ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_sll_srl_sra$_DFFE_PP_  (.CLK(clknet_leaf_489_clk),
    .RESET_B(net1698),
    .D(_01779_),
    .Q_N(_12388_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_sll_srl_sra ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_slli_srli_srai$_DFFE_PP_  (.CLK(clknet_leaf_488_clk),
    .RESET_B(net1699),
    .D(_01780_),
    .Q_N(_14058_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_slli_srli_srai ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_slti_blt_slt$_DFF_P_  (.CLK(clknet_leaf_492_clk),
    .RESET_B(net1700),
    .D(_00046_),
    .Q_N(_14059_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_slti_blt_slt ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.is_sltiu_bltu_sltu$_DFF_P_  (.CLK(clknet_leaf_627_clk),
    .RESET_B(net1701),
    .D(_00047_),
    .Q_N(_12387_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.is_sltiu_bltu_sltu ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.latched_branch$_SDFFE_PN0P_  (.CLK(clknet_leaf_482_clk),
    .RESET_B(net1702),
    .D(_01781_),
    .Q_N(_12386_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.latched_branch ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.latched_is_lb$_SDFFE_PN0P_  (.CLK(clknet_leaf_475_clk),
    .RESET_B(net1703),
    .D(_01782_),
    .Q_N(_12385_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.latched_is_lb ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.latched_is_lh$_SDFFE_PN0P_  (.CLK(clknet_leaf_474_clk),
    .RESET_B(net1704),
    .D(_01783_),
    .Q_N(_12384_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.latched_is_lh ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.latched_rd[0]$_SDFFCE_PP0P_  (.CLK(clknet_8_157_0_clk),
    .RESET_B(net1705),
    .D(_01784_),
    .Q_N(_12383_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.latched_rd[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.latched_rd[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_968_clk),
    .RESET_B(net1706),
    .D(_01785_),
    .Q_N(_12382_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.latched_rd[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.latched_rd[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_965_clk),
    .RESET_B(net1707),
    .D(_01786_),
    .Q_N(_00084_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.latched_rd[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.latched_rd[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_965_clk),
    .RESET_B(net1708),
    .D(_01787_),
    .Q_N(_12381_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.latched_rd[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.latched_rd[4]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_995_clk),
    .RESET_B(net1709),
    .D(_01788_),
    .Q_N(_12380_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.latched_rd[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.latched_stalu$_SDFFE_PN0P_  (.CLK(clknet_8_247_0_clk),
    .RESET_B(net1710),
    .D(_01789_),
    .Q_N(_12379_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.latched_stalu ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.latched_store$_SDFFE_PN0P_  (.CLK(clknet_leaf_481_clk),
    .RESET_B(net1711),
    .D(_01790_),
    .Q_N(_12378_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.latched_store ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[10]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1712),
    .D(_01791_),
    .Q_N(_12377_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[11]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1713),
    .D(_01792_),
    .Q_N(_12376_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[12]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1714),
    .D(_01793_),
    .Q_N(_12375_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[13]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1715),
    .D(_01794_),
    .Q_N(_12374_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[14]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1716),
    .D(_01795_),
    .Q_N(_12373_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[15]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1717),
    .D(_01796_),
    .Q_N(_12372_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[16]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1718),
    .D(_01797_),
    .Q_N(_12371_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[17]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1719),
    .D(_01798_),
    .Q_N(_12370_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[18]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1720),
    .D(_01799_),
    .Q_N(_12369_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[19]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1721),
    .D(_01800_),
    .Q_N(_12368_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[20]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1722),
    .D(_01801_),
    .Q_N(_12367_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[21]$_DFFE_PP_  (.CLK(clknet_8_97_0_clk),
    .RESET_B(net1723),
    .D(_01802_),
    .Q_N(_12366_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[22]$_DFFE_PP_  (.CLK(clknet_leaf_444_clk),
    .RESET_B(net1724),
    .D(_01803_),
    .Q_N(_12365_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[23]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1725),
    .D(_01804_),
    .Q_N(_12364_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[24]$_DFFE_PP_  (.CLK(clknet_leaf_443_clk),
    .RESET_B(net1726),
    .D(_01805_),
    .Q_N(_12363_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[25]$_DFFE_PP_  (.CLK(clknet_leaf_428_clk),
    .RESET_B(net1727),
    .D(_01806_),
    .Q_N(_12362_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[26]$_DFFE_PP_  (.CLK(clknet_leaf_440_clk),
    .RESET_B(net1728),
    .D(_01807_),
    .Q_N(_12361_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[27]$_DFFE_PP_  (.CLK(clknet_leaf_426_clk),
    .RESET_B(net1729),
    .D(_01808_),
    .Q_N(_12360_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[28]$_DFFE_PP_  (.CLK(clknet_leaf_426_clk),
    .RESET_B(net1730),
    .D(_01809_),
    .Q_N(_00104_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[29]$_DFFE_PP_  (.CLK(clknet_leaf_426_clk),
    .RESET_B(net1731),
    .D(_01810_),
    .Q_N(_00105_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[2]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1732),
    .D(_01811_),
    .Q_N(_12359_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[30]$_DFFE_PP_  (.CLK(clknet_leaf_425_clk),
    .RESET_B(net1733),
    .D(_01812_),
    .Q_N(_12358_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[31]$_DFFE_PP_  (.CLK(clknet_leaf_425_clk),
    .RESET_B(net1734),
    .D(_01813_),
    .Q_N(_12357_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[3]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1735),
    .D(_01814_),
    .Q_N(_12356_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[4]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1736),
    .D(_01815_),
    .Q_N(_12355_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[5]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1737),
    .D(_01816_),
    .Q_N(_12354_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[6]$_DFFE_PP_  (.CLK(clknet_8_78_0_clk),
    .RESET_B(net1738),
    .D(_01817_),
    .Q_N(_12353_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[7]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1739),
    .D(_01818_),
    .Q_N(_12352_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[8]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1740),
    .D(_01819_),
    .Q_N(_12351_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_addr[9]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1741),
    .D(_01820_),
    .Q_N(_12350_),
    .Q(\u_ac_controller_soc_inst.cbus_addr[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_do_prefetch$_SDFFE_PP0P_  (.CLK(clknet_8_208_0_clk),
    .RESET_B(net1742),
    .D(_01821_),
    .Q_N(_00085_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_do_prefetch ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_do_rdata$_SDFFE_PP1P_  (.CLK(clknet_leaf_474_clk),
    .RESET_B(net1743),
    .D(_01822_),
    .Q_N(_12349_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_do_rdata ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_do_rinst$_SDFFE_PP1P_  (.CLK(clknet_8_110_0_clk),
    .RESET_B(net1744),
    .D(_01823_),
    .Q_N(_00087_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_do_rinst ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_do_wdata$_SDFFE_PP1P_  (.CLK(clknet_leaf_434_clk),
    .RESET_B(net1745),
    .D(_01824_),
    .Q_N(_00112_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_do_wdata ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[0]$_DFFE_PP_  (.CLK(clknet_leaf_387_clk),
    .RESET_B(net1746),
    .D(_00113_),
    .Q_N(_12348_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[10]$_DFFE_PP_  (.CLK(clknet_leaf_452_clk),
    .RESET_B(net1747),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[10] ),
    .Q_N(_12347_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[11]$_DFFE_PP_  (.CLK(clknet_8_106_0_clk),
    .RESET_B(net1748),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[11] ),
    .Q_N(_12346_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[12]$_DFFE_PP_  (.CLK(clknet_leaf_519_clk),
    .RESET_B(net1749),
    .D(_08474_),
    .Q_N(_12345_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[13]$_DFFE_PP_  (.CLK(clknet_leaf_518_clk),
    .RESET_B(net1750),
    .D(_08468_),
    .Q_N(_12344_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[14]$_DFFE_PP_  (.CLK(clknet_leaf_517_clk),
    .RESET_B(net1751),
    .D(_08480_),
    .Q_N(_00121_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[15]$_DFFE_PP_  (.CLK(clknet_8_195_0_clk),
    .RESET_B(net1752),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[15] ),
    .Q_N(_12343_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[16]$_DFFE_PP_  (.CLK(clknet_leaf_463_clk),
    .RESET_B(net1753),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[16] ),
    .Q_N(_12342_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[17]$_DFFE_PP_  (.CLK(clknet_leaf_634_clk),
    .RESET_B(net1754),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[17] ),
    .Q_N(_12341_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[18]$_DFFE_PP_  (.CLK(clknet_8_193_0_clk),
    .RESET_B(net1755),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[18] ),
    .Q_N(_12340_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[19]$_DFFE_PP_  (.CLK(clknet_leaf_633_clk),
    .RESET_B(net1756),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[19] ),
    .Q_N(_12339_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[1]$_DFFE_PP_  (.CLK(clknet_leaf_387_clk),
    .RESET_B(net1757),
    .D(_00114_),
    .Q_N(_12338_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[20]$_DFFE_PP_  (.CLK(clknet_8_193_0_clk),
    .RESET_B(net1758),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[20] ),
    .Q_N(_12337_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[21]$_DFFE_PP_  (.CLK(clknet_leaf_469_clk),
    .RESET_B(net1759),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[21] ),
    .Q_N(_12336_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[22]$_DFFE_PP_  (.CLK(clknet_leaf_439_clk),
    .RESET_B(net1760),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[22] ),
    .Q_N(_12335_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[23]$_DFFE_PP_  (.CLK(clknet_leaf_440_clk),
    .RESET_B(net1761),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[23] ),
    .Q_N(_12334_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[24]$_DFFE_PP_  (.CLK(clknet_leaf_440_clk),
    .RESET_B(net1762),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[24] ),
    .Q_N(_12333_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[25]$_DFFE_PP_  (.CLK(clknet_leaf_435_clk),
    .RESET_B(net1763),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[25] ),
    .Q_N(_12332_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[26]$_DFFE_PP_  (.CLK(clknet_leaf_438_clk),
    .RESET_B(net1764),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[26] ),
    .Q_N(_12331_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27]$_DFFE_PP_  (.CLK(clknet_leaf_435_clk),
    .RESET_B(net1765),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[27] ),
    .Q_N(_12330_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[28]$_DFFE_PP_  (.CLK(clknet_leaf_436_clk),
    .RESET_B(net1766),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[28] ),
    .Q_N(_12329_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[29]$_DFFE_PP_  (.CLK(clknet_leaf_436_clk),
    .RESET_B(net1767),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[29] ),
    .Q_N(_12328_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[2]$_DFFE_PP_  (.CLK(clknet_8_209_0_clk),
    .RESET_B(net1768),
    .D(_00115_),
    .Q_N(_12327_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[30]$_DFFE_PP_  (.CLK(clknet_leaf_470_clk),
    .RESET_B(net1769),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[30] ),
    .Q_N(_12326_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[31]$_DFFE_PP_  (.CLK(clknet_leaf_485_clk),
    .RESET_B(net1770),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[31] ),
    .Q_N(_12325_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[3]$_DFFE_PP_  (.CLK(clknet_leaf_523_clk),
    .RESET_B(net1771),
    .D(_08441_),
    .Q_N(_12324_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[4]$_DFFE_PP_  (.CLK(clknet_leaf_525_clk),
    .RESET_B(net1772),
    .D(_08449_),
    .Q_N(_12323_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[5]$_DFFE_PP_  (.CLK(clknet_leaf_523_clk),
    .RESET_B(net1773),
    .D(_08455_),
    .Q_N(_12322_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[6]$_DFFE_PP_  (.CLK(clknet_leaf_525_clk),
    .RESET_B(net1774),
    .D(_08460_),
    .Q_N(_12321_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[7]$_DFFE_PP_  (.CLK(clknet_leaf_467_clk),
    .RESET_B(net1775),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[7] ),
    .Q_N(_12320_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[8]$_DFFE_PP_  (.CLK(clknet_leaf_437_clk),
    .RESET_B(net1776),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[8] ),
    .Q_N(_12319_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[9]$_DFFE_PP_  (.CLK(clknet_leaf_438_clk),
    .RESET_B(net1777),
    .D(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_latched[9] ),
    .Q_N(_12318_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_state[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_388_clk),
    .RESET_B(net1778),
    .D(_01825_),
    .Q_N(_12317_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_state[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_state[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_388_clk),
    .RESET_B(net1779),
    .D(_01826_),
    .Q_N(_12316_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_state[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_valid$_SDFFCE_PN0P_  (.CLK(clknet_8_105_0_clk),
    .RESET_B(net1780),
    .D(_01827_),
    .Q_N(_00086_),
    .Q(\u_ac_controller_soc_inst.cbus_valid ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1781),
    .D(_01828_),
    .Q_N(_12315_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1782),
    .D(_01829_),
    .Q_N(_12314_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1783),
    .D(_01830_),
    .Q_N(_12313_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1784),
    .D(_01831_),
    .Q_N(_12312_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1785),
    .D(_01832_),
    .Q_N(_12311_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1786),
    .D(_01833_),
    .Q_N(_12310_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1787),
    .D(_01834_),
    .Q_N(_12309_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[16]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1788),
    .D(_01835_),
    .Q_N(_12308_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[17]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1789),
    .D(_01836_),
    .Q_N(_12307_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[18]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1790),
    .D(_01837_),
    .Q_N(_12306_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[19]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1791),
    .D(_01838_),
    .Q_N(_12305_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1792),
    .D(_01839_),
    .Q_N(_12304_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[20]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1793),
    .D(_01840_),
    .Q_N(_12303_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[21]$_DFFE_PP_  (.CLK(clknet_8_27_0_clk),
    .RESET_B(net1794),
    .D(_01841_),
    .Q_N(_12302_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[22]$_DFFE_PP_  (.CLK(clknet_8_27_0_clk),
    .RESET_B(net1795),
    .D(_01842_),
    .Q_N(_12301_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[23]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1796),
    .D(_01843_),
    .Q_N(_12300_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[24]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1797),
    .D(_01844_),
    .Q_N(_12299_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[25]$_DFFE_PP_  (.CLK(clknet_8_27_0_clk),
    .RESET_B(net1798),
    .D(_01845_),
    .Q_N(_12298_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[26]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1799),
    .D(_01846_),
    .Q_N(_12297_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[27]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1800),
    .D(_01847_),
    .Q_N(_12296_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[28]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1801),
    .D(_01848_),
    .Q_N(_12295_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[29]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1802),
    .D(_01849_),
    .Q_N(_12294_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1803),
    .D(_01850_),
    .Q_N(_12293_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[30]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1804),
    .D(_01851_),
    .Q_N(_12292_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[31]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1805),
    .D(_01852_),
    .Q_N(_12291_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1806),
    .D(_01853_),
    .Q_N(_12290_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1807),
    .D(_01854_),
    .Q_N(_12289_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1808),
    .D(_01855_),
    .Q_N(_12288_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1809),
    .D(_01856_),
    .Q_N(_12287_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1810),
    .D(_01857_),
    .Q_N(_12286_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1811),
    .D(_01858_),
    .Q_N(_12285_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1812),
    .D(_01859_),
    .Q_N(_14060_),
    .Q(\u_ac_controller_soc_inst.cbus_wdata[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wordsize[0]$_DFF_P_  (.CLK(clknet_leaf_473_clk),
    .RESET_B(net1813),
    .D(_00017_),
    .Q_N(_14061_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wordsize[1]$_DFF_P_  (.CLK(clknet_leaf_434_clk),
    .RESET_B(net1814),
    .D(_00018_),
    .Q_N(_00129_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wordsize[2]$_DFF_P_  (.CLK(clknet_leaf_433_clk),
    .RESET_B(net1815),
    .D(_00019_),
    .Q_N(_00052_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_wordsize[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wstrb[0]$_DFFE_PP_  (.CLK(clknet_8_102_0_clk),
    .RESET_B(net1816),
    .D(_01860_),
    .Q_N(_00106_),
    .Q(\u_ac_controller_soc_inst.cbus_wstrb[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wstrb[1]$_DFFE_PP_  (.CLK(clknet_leaf_427_clk),
    .RESET_B(net1817),
    .D(_01861_),
    .Q_N(_12284_),
    .Q(\u_ac_controller_soc_inst.cbus_wstrb[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wstrb[2]$_DFFE_PP_  (.CLK(clknet_leaf_427_clk),
    .RESET_B(net1818),
    .D(_01862_),
    .Q_N(_12283_),
    .Q(\u_ac_controller_soc_inst.cbus_wstrb[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.mem_wstrb[3]$_DFFE_PP_  (.CLK(clknet_leaf_427_clk),
    .RESET_B(net1819),
    .D(_01863_),
    .Q_N(_12282_),
    .Q(\u_ac_controller_soc_inst.cbus_wstrb[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_457_clk),
    .RESET_B(net1820),
    .D(_01864_),
    .Q_N(_12281_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[11]$_SDFFE_PN0P_  (.CLK(clknet_8_194_0_clk),
    .RESET_B(net1821),
    .D(_01865_),
    .Q_N(_12280_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_445_clk),
    .RESET_B(net1822),
    .D(_01866_),
    .Q_N(_12279_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[13]$_SDFFE_PN0P_  (.CLK(clknet_8_245_0_clk),
    .RESET_B(net1823),
    .D(_01867_),
    .Q_N(_12278_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_461_clk),
    .RESET_B(net1824),
    .D(_01868_),
    .Q_N(_12277_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_461_clk),
    .RESET_B(net1825),
    .D(_01869_),
    .Q_N(_12276_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_650_clk),
    .RESET_B(net1826),
    .D(_01870_),
    .Q_N(_12275_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_648_clk),
    .RESET_B(net1827),
    .D(_01871_),
    .Q_N(_12274_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_633_clk),
    .RESET_B(net1828),
    .D(_01872_),
    .Q_N(_12273_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_631_clk),
    .RESET_B(net1829),
    .D(_01873_),
    .Q_N(_12272_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1830),
    .D(_01874_),
    .Q_N(_12271_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[20]$_SDFFE_PN0P_  (.CLK(clknet_8_201_0_clk),
    .RESET_B(net1831),
    .D(_01875_),
    .Q_N(_12270_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[21]$_SDFFE_PN0P_  (.CLK(clknet_8_255_0_clk),
    .RESET_B(net1832),
    .D(_01876_),
    .Q_N(_12269_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[22]$_SDFFE_PN0P_  (.CLK(clknet_8_228_0_clk),
    .RESET_B(net1833),
    .D(_01877_),
    .Q_N(_12268_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_615_clk),
    .RESET_B(net1834),
    .D(_01878_),
    .Q_N(_12267_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_599_clk),
    .RESET_B(net1835),
    .D(_01879_),
    .Q_N(_12266_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[25]$_SDFFE_PN0P_  (.CLK(clknet_8_202_0_clk),
    .RESET_B(net1836),
    .D(_01880_),
    .Q_N(_12265_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[26]$_SDFFE_PN0P_  (.CLK(clknet_8_202_0_clk),
    .RESET_B(net1837),
    .D(_01881_),
    .Q_N(_12264_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_615_clk),
    .RESET_B(net1838),
    .D(_01882_),
    .Q_N(_12263_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_594_clk),
    .RESET_B(net1839),
    .D(_01883_),
    .Q_N(_12262_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[29]$_SDFFE_PN0P_  (.CLK(clknet_8_201_0_clk),
    .RESET_B(net1840),
    .D(_01884_),
    .Q_N(_12261_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[2]$_SDFFE_PN0P_  (.CLK(clknet_8_98_0_clk),
    .RESET_B(net1841),
    .D(_01885_),
    .Q_N(_12260_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_594_clk),
    .RESET_B(net1842),
    .D(_01886_),
    .Q_N(_12259_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[31]$_SDFFE_PN0P_  (.CLK(clknet_8_200_0_clk),
    .RESET_B(net1843),
    .D(_01887_),
    .Q_N(_12258_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1844),
    .D(_01888_),
    .Q_N(_12257_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1845),
    .D(_01889_),
    .Q_N(_12256_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[5]$_SDFFE_PN0P_  (.CLK(clknet_8_96_0_clk),
    .RESET_B(net1846),
    .D(_01890_),
    .Q_N(_12255_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1847),
    .D(_01891_),
    .Q_N(_12254_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1848),
    .D(_01892_),
    .Q_N(_12253_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_446_clk),
    .RESET_B(net1849),
    .D(_01893_),
    .Q_N(_12252_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_445_clk),
    .RESET_B(net1850),
    .D(_01894_),
    .Q_N(_12251_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_next_pc[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[0]$_DFFE_PP_  (.CLK(clknet_8_240_0_clk),
    .RESET_B(net1851),
    .D(_01895_),
    .Q_N(_00056_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[10]$_DFFE_PP_  (.CLK(clknet_8_151_0_clk),
    .RESET_B(net1852),
    .D(_01896_),
    .Q_N(_00064_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[11]$_DFFE_PP_  (.CLK(clknet_8_242_0_clk),
    .RESET_B(net1853),
    .D(_01897_),
    .Q_N(_00065_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[12]$_DFFE_PP_  (.CLK(clknet_8_157_0_clk),
    .RESET_B(net1854),
    .D(_01898_),
    .Q_N(_00066_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[13]$_DFFE_PP_  (.CLK(clknet_leaf_969_clk),
    .RESET_B(net1855),
    .D(_01899_),
    .Q_N(_00067_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[14]$_DFFE_PP_  (.CLK(clknet_8_242_0_clk),
    .RESET_B(net1856),
    .D(_01900_),
    .Q_N(_00068_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[15]$_DFFE_PP_  (.CLK(clknet_leaf_972_clk),
    .RESET_B(net1857),
    .D(_01901_),
    .Q_N(_00069_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[16]$_DFFE_PP_  (.CLK(clknet_leaf_972_clk),
    .RESET_B(net1858),
    .D(_01902_),
    .Q_N(_00070_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[17]$_DFFE_PP_  (.CLK(clknet_8_159_0_clk),
    .RESET_B(net1859),
    .D(_01903_),
    .Q_N(_00071_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[18]$_DFFE_PP_  (.CLK(clknet_leaf_955_clk),
    .RESET_B(net1860),
    .D(_01904_),
    .Q_N(_00072_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[19]$_DFFE_PP_  (.CLK(clknet_8_248_0_clk),
    .RESET_B(net1861),
    .D(_01905_),
    .Q_N(_00073_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[1]$_DFFE_PP_  (.CLK(clknet_leaf_988_clk),
    .RESET_B(net1862),
    .D(_01906_),
    .Q_N(_00053_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[20]$_DFFE_PP_  (.CLK(clknet_leaf_954_clk),
    .RESET_B(net1863),
    .D(_01907_),
    .Q_N(_00074_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[21]$_DFFE_PP_  (.CLK(clknet_leaf_954_clk),
    .RESET_B(net1864),
    .D(_01908_),
    .Q_N(_00075_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[22]$_DFFE_PP_  (.CLK(clknet_8_249_0_clk),
    .RESET_B(net1865),
    .D(_01909_),
    .Q_N(_00076_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[23]$_DFFE_PP_  (.CLK(clknet_leaf_671_clk),
    .RESET_B(net1866),
    .D(_01910_),
    .Q_N(_00077_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[24]$_DFFE_PP_  (.CLK(clknet_leaf_671_clk),
    .RESET_B(net1867),
    .D(_01911_),
    .Q_N(_00078_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[25]$_DFFE_PP_  (.CLK(clknet_8_249_0_clk),
    .RESET_B(net1868),
    .D(_01912_),
    .Q_N(_00079_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[26]$_DFFE_PP_  (.CLK(clknet_8_250_0_clk),
    .RESET_B(net1869),
    .D(_01913_),
    .Q_N(_00080_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[27]$_DFFE_PP_  (.CLK(clknet_8_249_0_clk),
    .RESET_B(net1870),
    .D(_01914_),
    .Q_N(_00081_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[28]$_DFFE_PP_  (.CLK(clknet_leaf_676_clk),
    .RESET_B(net1871),
    .D(_01915_),
    .Q_N(_00082_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[29]$_DFFE_PP_  (.CLK(clknet_leaf_676_clk),
    .RESET_B(net1872),
    .D(_01916_),
    .Q_N(_00083_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[2]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1873),
    .D(_01917_),
    .Q_N(_00057_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[30]$_DFFE_PP_  (.CLK(clknet_leaf_699_clk),
    .RESET_B(net1874),
    .D(_01918_),
    .Q_N(_12250_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[31]$_DFFE_PP_  (.CLK(clknet_leaf_669_clk),
    .RESET_B(net1875),
    .D(_01919_),
    .Q_N(_12249_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[3]$_DFFE_PP_  (.CLK(clknet_leaf_988_clk),
    .RESET_B(net1876),
    .D(_01920_),
    .Q_N(_00059_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[4]$_DFFE_PP_  (.CLK(clknet_leaf_990_clk),
    .RESET_B(net1877),
    .D(_01921_),
    .Q_N(_00055_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[5]$_DFFE_PP_  (.CLK(clknet_8_149_0_clk),
    .RESET_B(net1878),
    .D(_01922_),
    .Q_N(_00058_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[6]$_DFFE_PP_  (.CLK(clknet_leaf_988_clk),
    .RESET_B(net1879),
    .D(_01923_),
    .Q_N(_00060_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[7]$_DFFE_PP_  (.CLK(clknet_8_151_0_clk),
    .RESET_B(net1880),
    .D(_01924_),
    .Q_N(_00061_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[8]$_DFFE_PP_  (.CLK(clknet_8_240_0_clk),
    .RESET_B(net1881),
    .D(_01925_),
    .Q_N(_00062_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op1[9]$_DFFE_PP_  (.CLK(clknet_8_151_0_clk),
    .RESET_B(net1882),
    .D(_01926_),
    .Q_N(_00063_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs1[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[0]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1883),
    .D(_01927_),
    .Q_N(_12248_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[10]$_DFFE_PP_  (.CLK(clknet_8_241_0_clk),
    .RESET_B(net1884),
    .D(_01928_),
    .Q_N(_12247_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[11]$_DFFE_PP_  (.CLK(clknet_leaf_978_clk),
    .RESET_B(net1885),
    .D(_01929_),
    .Q_N(_12246_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[12]$_DFFE_PP_  (.CLK(clknet_leaf_982_clk),
    .RESET_B(net1886),
    .D(_01930_),
    .Q_N(_12245_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[13]$_DFFE_PP_  (.CLK(clknet_leaf_978_clk),
    .RESET_B(net1887),
    .D(_01931_),
    .Q_N(_12244_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[14]$_DFFE_PP_  (.CLK(clknet_leaf_974_clk),
    .RESET_B(net1888),
    .D(_01932_),
    .Q_N(_12243_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[15]$_DFFE_PP_  (.CLK(clknet_leaf_974_clk),
    .RESET_B(net1889),
    .D(_01933_),
    .Q_N(_12242_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[16]$_DFFE_PP_  (.CLK(clknet_8_243_0_clk),
    .RESET_B(net1890),
    .D(_01934_),
    .Q_N(_12241_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[17]$_DFFE_PP_  (.CLK(clknet_8_243_0_clk),
    .RESET_B(net1891),
    .D(_01935_),
    .Q_N(_12240_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[18]$_DFFE_PP_  (.CLK(clknet_8_243_0_clk),
    .RESET_B(net1892),
    .D(_01936_),
    .Q_N(_12239_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[19]$_DFFE_PP_  (.CLK(clknet_leaf_666_clk),
    .RESET_B(net1893),
    .D(_01937_),
    .Q_N(_12238_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[1]$_DFFE_PP_  (.CLK(clknet_8_26_0_clk),
    .RESET_B(net1894),
    .D(_01938_),
    .Q_N(_12237_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[20]$_DFFE_PP_  (.CLK(clknet_leaf_668_clk),
    .RESET_B(net1895),
    .D(_01939_),
    .Q_N(_12236_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[21]$_DFFE_PP_  (.CLK(clknet_leaf_668_clk),
    .RESET_B(net1896),
    .D(_01940_),
    .Q_N(_12235_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[22]$_DFFE_PP_  (.CLK(clknet_leaf_666_clk),
    .RESET_B(net1897),
    .D(_01941_),
    .Q_N(_12234_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[23]$_DFFE_PP_  (.CLK(clknet_leaf_667_clk),
    .RESET_B(net1898),
    .D(_01942_),
    .Q_N(_12233_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[24]$_DFFE_PP_  (.CLK(clknet_leaf_667_clk),
    .RESET_B(net1899),
    .D(_01943_),
    .Q_N(_12232_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[25]$_DFFE_PP_  (.CLK(clknet_leaf_700_clk),
    .RESET_B(net1900),
    .D(_01944_),
    .Q_N(_12231_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[26]$_DFFE_PP_  (.CLK(clknet_leaf_703_clk),
    .RESET_B(net1901),
    .D(_01945_),
    .Q_N(_12230_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[27]$_DFFE_PP_  (.CLK(clknet_leaf_669_clk),
    .RESET_B(net1902),
    .D(_01946_),
    .Q_N(_12229_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[28]$_DFFE_PP_  (.CLK(clknet_leaf_703_clk),
    .RESET_B(net1903),
    .D(_01947_),
    .Q_N(_12228_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[29]$_DFFE_PP_  (.CLK(clknet_leaf_700_clk),
    .RESET_B(net1904),
    .D(_01948_),
    .Q_N(_12227_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[2]$_DFFE_PP_  (.CLK(clknet_8_15_0_clk),
    .RESET_B(net1905),
    .D(_01949_),
    .Q_N(_12226_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[30]$_DFFE_PP_  (.CLK(clknet_leaf_699_clk),
    .RESET_B(net1906),
    .D(_01950_),
    .Q_N(_12225_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[31]$_DFFE_PP_  (.CLK(clknet_leaf_703_clk),
    .RESET_B(net1907),
    .D(_01951_),
    .Q_N(_12224_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[3]$_DFFE_PP_  (.CLK(clknet_8_26_0_clk),
    .RESET_B(net1908),
    .D(_01952_),
    .Q_N(_12223_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[4]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1909),
    .D(_01953_),
    .Q_N(_12222_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[5]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1910),
    .D(_01954_),
    .Q_N(_12221_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[6]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1911),
    .D(_01955_),
    .Q_N(_12220_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[7]$_DFFE_PP_  (.CLK(clknet_8_240_0_clk),
    .RESET_B(net1912),
    .D(_01956_),
    .Q_N(_12219_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.mem_la_wdata[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[8]$_DFFE_PP_  (.CLK(clknet_leaf_982_clk),
    .RESET_B(net1913),
    .D(_01957_),
    .Q_N(_12218_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_op2[9]$_DFFE_PP_  (.CLK(clknet_8_241_0_clk),
    .RESET_B(net1914),
    .D(_01958_),
    .Q_N(_14062_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.pcpi_rs2[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[0]$_DFF_P_  (.CLK(clknet_leaf_473_clk),
    .RESET_B(net1915),
    .D(_02144_),
    .Q_N(_14063_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[10]$_DFF_P_  (.CLK(clknet_leaf_470_clk),
    .RESET_B(net1916),
    .D(_02145_),
    .Q_N(_14064_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[11]$_DFF_P_  (.CLK(clknet_leaf_469_clk),
    .RESET_B(net1917),
    .D(_02146_),
    .Q_N(_14065_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[12]$_DFF_P_  (.CLK(clknet_leaf_446_clk),
    .RESET_B(net1918),
    .D(_02147_),
    .Q_N(_14066_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[13]$_DFF_P_  (.CLK(clknet_leaf_456_clk),
    .RESET_B(net1919),
    .D(_02148_),
    .Q_N(_14067_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[14]$_DFF_P_  (.CLK(clknet_leaf_466_clk),
    .RESET_B(net1920),
    .D(_02149_),
    .Q_N(_14068_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[15]$_DFF_P_  (.CLK(clknet_leaf_464_clk),
    .RESET_B(net1921),
    .D(_02150_),
    .Q_N(_14069_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[16]$_DFF_P_  (.CLK(clknet_leaf_463_clk),
    .RESET_B(net1922),
    .D(_02151_),
    .Q_N(_14070_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[17]$_DFF_P_  (.CLK(clknet_8_195_0_clk),
    .RESET_B(net1923),
    .D(_02152_),
    .Q_N(_14071_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[18]$_DFF_P_  (.CLK(clknet_leaf_634_clk),
    .RESET_B(net1924),
    .D(_02153_),
    .Q_N(_14072_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[19]$_DFF_P_  (.CLK(clknet_leaf_627_clk),
    .RESET_B(net1925),
    .D(_02154_),
    .Q_N(_14073_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[1]$_DFF_P_  (.CLK(clknet_leaf_446_clk),
    .RESET_B(net1926),
    .D(_02155_),
    .Q_N(_14074_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[20]$_DFF_P_  (.CLK(clknet_leaf_622_clk),
    .RESET_B(net1927),
    .D(_02156_),
    .Q_N(_14075_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[21]$_DFF_P_  (.CLK(clknet_8_207_0_clk),
    .RESET_B(net1928),
    .D(_02157_),
    .Q_N(_14076_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[22]$_DFF_P_  (.CLK(clknet_leaf_622_clk),
    .RESET_B(net1929),
    .D(_02158_),
    .Q_N(_14077_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[23]$_DFF_P_  (.CLK(clknet_leaf_620_clk),
    .RESET_B(net1930),
    .D(_02159_),
    .Q_N(_14078_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[24]$_DFF_P_  (.CLK(clknet_8_201_0_clk),
    .RESET_B(net1931),
    .D(_02160_),
    .Q_N(_14079_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[25]$_DFF_P_  (.CLK(clknet_leaf_620_clk),
    .RESET_B(net1932),
    .D(_02161_),
    .Q_N(_14080_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[26]$_DFF_P_  (.CLK(clknet_leaf_620_clk),
    .RESET_B(net1933),
    .D(_02162_),
    .Q_N(_14081_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[27]$_DFF_P_  (.CLK(clknet_leaf_615_clk),
    .RESET_B(net1934),
    .D(_02163_),
    .Q_N(_14082_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[28]$_DFF_P_  (.CLK(clknet_leaf_618_clk),
    .RESET_B(net1935),
    .D(_02164_),
    .Q_N(_14083_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[29]$_DFF_P_  (.CLK(clknet_leaf_618_clk),
    .RESET_B(net1936),
    .D(_02165_),
    .Q_N(_14084_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[2]$_DFF_P_  (.CLK(clknet_leaf_443_clk),
    .RESET_B(net1937),
    .D(_02166_),
    .Q_N(_14085_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[30]$_DFF_P_  (.CLK(clknet_leaf_618_clk),
    .RESET_B(net1938),
    .D(_02167_),
    .Q_N(_14086_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[31]$_DFF_P_  (.CLK(clknet_8_204_0_clk),
    .RESET_B(net1939),
    .D(_02168_),
    .Q_N(_14087_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[3]$_DFF_P_  (.CLK(clknet_leaf_444_clk),
    .RESET_B(net1940),
    .D(_02169_),
    .Q_N(_14088_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[4]$_DFF_P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1941),
    .D(_02170_),
    .Q_N(_14089_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[5]$_DFF_P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1942),
    .D(_02171_),
    .Q_N(_14090_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[6]$_DFF_P_  (.CLK(clknet_leaf_445_clk),
    .RESET_B(net1943),
    .D(_02172_),
    .Q_N(_14091_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[7]$_DFF_P_  (.CLK(clknet_leaf_442_clk),
    .RESET_B(net1944),
    .D(_02173_),
    .Q_N(_14092_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[8]$_DFF_P_  (.CLK(clknet_8_104_0_clk),
    .RESET_B(net1945),
    .D(_02174_),
    .Q_N(_14093_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_out[9]$_DFF_P_  (.CLK(clknet_leaf_442_clk),
    .RESET_B(net1946),
    .D(_02175_),
    .Q_N(_12217_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_out[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[10]$_SDFFE_PN0P_  (.CLK(clknet_8_244_0_clk),
    .RESET_B(net1947),
    .D(_01959_),
    .Q_N(_12216_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_658_clk),
    .RESET_B(net1948),
    .D(_01960_),
    .Q_N(_12215_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_455_clk),
    .RESET_B(net1949),
    .D(_01961_),
    .Q_N(_12214_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_657_clk),
    .RESET_B(net1950),
    .D(_01962_),
    .Q_N(_12213_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_656_clk),
    .RESET_B(net1951),
    .D(_01963_),
    .Q_N(_12212_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[15]$_SDFFE_PN0P_  (.CLK(clknet_8_243_0_clk),
    .RESET_B(net1952),
    .D(_01964_),
    .Q_N(_12211_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_652_clk),
    .RESET_B(net1953),
    .D(_01965_),
    .Q_N(_12210_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_653_clk),
    .RESET_B(net1954),
    .D(_01966_),
    .Q_N(_12209_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_631_clk),
    .RESET_B(net1955),
    .D(_01967_),
    .Q_N(_12208_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_611_clk),
    .RESET_B(net1956),
    .D(_01968_),
    .Q_N(_12207_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1957),
    .D(_01969_),
    .Q_N(_12206_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_611_clk),
    .RESET_B(net1958),
    .D(_01970_),
    .Q_N(_12205_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_609_clk),
    .RESET_B(net1959),
    .D(_01971_),
    .Q_N(_12204_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_609_clk),
    .RESET_B(net1960),
    .D(_01972_),
    .Q_N(_12203_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[23]$_SDFFE_PN0P_  (.CLK(clknet_8_229_0_clk),
    .RESET_B(net1961),
    .D(_01973_),
    .Q_N(_12202_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_604_clk),
    .RESET_B(net1962),
    .D(_01974_),
    .Q_N(_12201_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_613_clk),
    .RESET_B(net1963),
    .D(_01975_),
    .Q_N(_12200_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[26]$_SDFFE_PN0P_  (.CLK(clknet_8_229_0_clk),
    .RESET_B(net1964),
    .D(_01976_),
    .Q_N(_12199_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_601_clk),
    .RESET_B(net1965),
    .D(_01977_),
    .Q_N(_12198_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_601_clk),
    .RESET_B(net1966),
    .D(_01978_),
    .Q_N(_12197_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_599_clk),
    .RESET_B(net1967),
    .D(_01979_),
    .Q_N(_12196_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1968),
    .D(_01980_),
    .Q_N(_00130_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_599_clk),
    .RESET_B(net1969),
    .D(_01981_),
    .Q_N(_12195_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[31]$_SDFFE_PN0P_  (.CLK(clknet_8_200_0_clk),
    .RESET_B(net1970),
    .D(_01982_),
    .Q_N(_12194_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1971),
    .D(_01983_),
    .Q_N(_12193_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[4]$_SDFFE_PN0P_  (.CLK(clknet_8_28_0_clk),
    .RESET_B(net1972),
    .D(_01984_),
    .Q_N(_12192_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[5]$_SDFFE_PN0P_  (.CLK(clknet_8_30_0_clk),
    .RESET_B(net1973),
    .D(_01985_),
    .Q_N(_12191_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1974),
    .D(_01986_),
    .Q_N(_12190_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1975),
    .D(_01987_),
    .Q_N(_12189_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1976),
    .D(_01988_),
    .Q_N(_12188_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_pc[9]$_SDFFE_PN0P_  (.CLK(clknet_8_28_0_clk),
    .RESET_B(net1977),
    .D(_01989_),
    .Q_N(_12187_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_pc[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_sh[0]$_DFFE_PP_  (.CLK(clknet_8_159_0_clk),
    .RESET_B(net1978),
    .D(_01990_),
    .Q_N(_12186_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_sh[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_sh[1]$_DFFE_PP_  (.CLK(clknet_8_156_0_clk),
    .RESET_B(net1979),
    .D(_01991_),
    .Q_N(_14094_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_sh[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_sh[2]$_DFF_P_  (.CLK(clknet_leaf_969_clk),
    .RESET_B(net1980),
    .D(_00048_),
    .Q_N(_00134_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_sh[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_sh[3]$_DFF_P_  (.CLK(clknet_leaf_966_clk),
    .RESET_B(net1981),
    .D(_00049_),
    .Q_N(_14095_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_sh[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.reg_sh[4]$_DFF_P_  (.CLK(clknet_leaf_966_clk),
    .RESET_B(net1982),
    .D(_00050_),
    .Q_N(_12185_),
    .Q(\u_ac_controller_soc_inst.u_picorv32.reg_sh[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_picorv32.trap$_SDFF_PN0_  (.CLK(clknet_leaf_475_clk),
    .RESET_B(net1983),
    .D(_01992_),
    .Q_N(_12184_),
    .Q(\u_ac_controller_soc_inst.trap ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[0]$_DFFE_PP_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1984),
    .D(_01993_),
    .Q_N(_12183_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[10]$_DFFE_PP_  (.CLK(clknet_8_114_0_clk),
    .RESET_B(net1985),
    .D(_01994_),
    .Q_N(_12182_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[11]$_DFFE_PP_  (.CLK(clknet_leaf_400_clk),
    .RESET_B(net1986),
    .D(_01995_),
    .Q_N(_12181_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[12]$_DFFE_PP_  (.CLK(clknet_leaf_404_clk),
    .RESET_B(net1987),
    .D(_01996_),
    .Q_N(_12180_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[13]$_DFFE_PP_  (.CLK(clknet_leaf_396_clk),
    .RESET_B(net1988),
    .D(_01997_),
    .Q_N(_12179_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[14]$_DFFE_PP_  (.CLK(clknet_leaf_374_clk),
    .RESET_B(net1989),
    .D(_01998_),
    .Q_N(_12178_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[15]$_DFFE_PP_  (.CLK(clknet_leaf_376_clk),
    .RESET_B(net1990),
    .D(_01999_),
    .Q_N(_12177_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[16]$_DFFE_PP_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1991),
    .D(_02000_),
    .Q_N(_12176_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[17]$_DFFE_PP_  (.CLK(clknet_8_120_0_clk),
    .RESET_B(net1992),
    .D(_02001_),
    .Q_N(_12175_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[18]$_DFFE_PP_  (.CLK(clknet_leaf_375_clk),
    .RESET_B(net1993),
    .D(_02002_),
    .Q_N(_12174_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[19]$_DFFE_PP_  (.CLK(clknet_leaf_380_clk),
    .RESET_B(net1994),
    .D(_02003_),
    .Q_N(_12173_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[1]$_DFFE_PP_  (.CLK(clknet_leaf_406_clk),
    .RESET_B(net1995),
    .D(_02004_),
    .Q_N(_12172_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[20]$_DFFE_PP_  (.CLK(clknet_leaf_398_clk),
    .RESET_B(net1996),
    .D(_02005_),
    .Q_N(_12171_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[21]$_DFFE_PP_  (.CLK(clknet_leaf_395_clk),
    .RESET_B(net1997),
    .D(_02006_),
    .Q_N(_12170_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[22]$_DFFE_PP_  (.CLK(clknet_leaf_375_clk),
    .RESET_B(net1998),
    .D(_02007_),
    .Q_N(_12169_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[23]$_DFFE_PP_  (.CLK(clknet_leaf_380_clk),
    .RESET_B(net1999),
    .D(_02008_),
    .Q_N(_12168_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[2]$_DFFE_PP_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2000),
    .D(_02009_),
    .Q_N(_12167_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[3]$_DFFE_PP_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2001),
    .D(_02010_),
    .Q_N(_12166_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[4]$_DFFE_PP_  (.CLK(clknet_8_112_0_clk),
    .RESET_B(net2002),
    .D(_02011_),
    .Q_N(_12165_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[5]$_DFFE_PP_  (.CLK(clknet_8_112_0_clk),
    .RESET_B(net2003),
    .D(_02012_),
    .Q_N(_12164_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[6]$_DFFE_PP_  (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2004),
    .D(_02013_),
    .Q_N(_12163_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[7]$_DFFE_PP_  (.CLK(clknet_leaf_403_clk),
    .RESET_B(net2005),
    .D(_02014_),
    .Q_N(_12162_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[8]$_DFFE_PP_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2006),
    .D(_02015_),
    .Q_N(_12161_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[9]$_DFFE_PP_  (.CLK(clknet_leaf_407_clk),
    .RESET_B(net2007),
    .D(_02016_),
    .Q_N(_12160_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.buffer[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_clk$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2008),
    .D(_02017_),
    .Q_N(_12159_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.config_clk ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_cont$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2009),
    .D(_02018_),
    .Q_N(_00098_),
    .Q(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_csb$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2010),
    .D(_02019_),
    .Q_N(_12158_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.config_csb ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_ddr$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2011),
    .D(_02020_),
    .Q_N(_12157_),
    .Q(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2012),
    .D(_02021_),
    .Q_N(_12156_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2013),
    .D(_02022_),
    .Q_N(_12155_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[2]$_SDFFE_PN0P_  (.CLK(clknet_8_68_0_clk),
    .RESET_B(net2014),
    .D(_02023_),
    .Q_N(_12154_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2015),
    .D(_02024_),
    .Q_N(_12153_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.config_do[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_dummy[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2016),
    .D(_02025_),
    .Q_N(_12152_),
    .Q(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_dummy[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2017),
    .D(_02026_),
    .Q_N(_12151_),
    .Q(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_dummy[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2018),
    .D(_02027_),
    .Q_N(_12150_),
    .Q(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_dummy[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2019),
    .D(_02028_),
    .Q_N(_12149_),
    .Q(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_en$_SDFFE_PN1P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2020),
    .D(_02029_),
    .Q_N(_00120_),
    .Q(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2021),
    .D(_02030_),
    .Q_N(_12148_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2022),
    .D(_02031_),
    .Q_N(_12147_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2023),
    .D(_02032_),
    .Q_N(_12146_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2024),
    .D(_02033_),
    .Q_N(_12145_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.config_qspi$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2025),
    .D(_02034_),
    .Q_N(_12144_),
    .Q(\u_ac_controller_soc_inst.spi_flash_cfg_rdata[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[0]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2026),
    .D(_02035_),
    .Q_N(_12143_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[1]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2027),
    .D(_02036_),
    .Q_N(_12142_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2028),
    .D(_02037_),
    .Q_N(_12141_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[3]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2029),
    .D(_02038_),
    .Q_N(_12140_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[4]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2030),
    .D(_02039_),
    .Q_N(_12139_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[5]$_SDFFCE_PN1P_  (.CLK(clknet_8_66_0_clk),
    .RESET_B(net2031),
    .D(_02040_),
    .Q_N(_12138_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[6]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2032),
    .D(_02041_),
    .Q_N(_12137_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[7]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2033),
    .D(_02042_),
    .Q_N(_12136_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_data[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_ddr$_SDFF_PP0_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2034),
    .D(_02043_),
    .Q_N(_12135_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_ddr ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_qspi$_SDFF_PP0_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2035),
    .D(_02044_),
    .Q_N(_12134_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_qspi ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_rd$_SDFFE_PP0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2036),
    .D(_02045_),
    .Q_N(_12133_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_rd ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2037),
    .D(_02046_),
    .Q_N(_12132_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2038),
    .D(_02047_),
    .Q_N(_12131_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2039),
    .D(_02048_),
    .Q_N(_12130_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.din_valid$_SDFF_PP0_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2040),
    .D(_02049_),
    .Q_N(_12129_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.din_valid ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[10]$_DFFE_PP_  (.CLK(clknet_8_22_0_clk),
    .RESET_B(net2041),
    .D(_02050_),
    .Q_N(_12128_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[11]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2042),
    .D(_02051_),
    .Q_N(_12127_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[12]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2043),
    .D(_02052_),
    .Q_N(_12126_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[13]$_DFFE_PP_  (.CLK(clknet_8_22_0_clk),
    .RESET_B(net2044),
    .D(_02053_),
    .Q_N(_12125_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[14]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2045),
    .D(_02054_),
    .Q_N(_12124_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2046),
    .D(_02055_),
    .Q_N(_12123_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[16]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2047),
    .D(_02056_),
    .Q_N(_12122_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[17]$_DFFE_PP_  (.CLK(clknet_8_25_0_clk),
    .RESET_B(net2048),
    .D(_02057_),
    .Q_N(_12121_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[18]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2049),
    .D(_02058_),
    .Q_N(_12120_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2050),
    .D(_02059_),
    .Q_N(_12119_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20]$_DFFE_PP_  (.CLK(clknet_8_74_0_clk),
    .RESET_B(net2051),
    .D(_02060_),
    .Q_N(_12118_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2052),
    .D(_02061_),
    .Q_N(_12117_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[22]$_DFFE_PP_  (.CLK(clknet_8_75_0_clk),
    .RESET_B(net2053),
    .D(_02062_),
    .Q_N(_12116_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23]$_DFFE_PP_  (.CLK(clknet_8_74_0_clk),
    .RESET_B(net2054),
    .D(_02063_),
    .Q_N(_12115_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2055),
    .D(_02064_),
    .Q_N(_00125_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2056),
    .D(_02065_),
    .Q_N(_12114_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[4]$_DFFE_PP_  (.CLK(clknet_8_22_0_clk),
    .RESET_B(net2057),
    .D(_02066_),
    .Q_N(_12113_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[5]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2058),
    .D(_02067_),
    .Q_N(_12112_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[6]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2059),
    .D(_02068_),
    .Q_N(_12111_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[7]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2060),
    .D(_02069_),
    .Q_N(_12110_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[8]$_DFFE_PP_  (.CLK(clknet_8_78_0_clk),
    .RESET_B(net2061),
    .D(_02070_),
    .Q_N(_12109_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[9]$_DFFE_PP_  (.CLK(clknet_8_78_0_clk),
    .RESET_B(net2062),
    .D(_02071_),
    .Q_N(_12108_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_inc$_SDFFCE_PP0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2063),
    .D(_02072_),
    .Q_N(_12107_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_inc ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_valid$_SDFFE_PP0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2064),
    .D(_02073_),
    .Q_N(_12106_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_valid ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rd_wait$_SDFFCE_PP0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2065),
    .D(_02074_),
    .Q_N(_12105_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.rd_wait ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_414_clk),
    .RESET_B(net2066),
    .D(_02075_),
    .Q_N(_12104_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_399_clk),
    .RESET_B(net2067),
    .D(_02076_),
    .Q_N(_12103_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_400_clk),
    .RESET_B(net2068),
    .D(_02077_),
    .Q_N(_12102_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_399_clk),
    .RESET_B(net2069),
    .D(_02078_),
    .Q_N(_12101_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_396_clk),
    .RESET_B(net2070),
    .D(_02079_),
    .Q_N(_12100_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[13] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_376_clk),
    .RESET_B(net2071),
    .D(_02080_),
    .Q_N(_12099_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[14] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_378_clk),
    .RESET_B(net2072),
    .D(_02081_),
    .Q_N(_12098_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[15] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[16]$_DFFE_PP_  (.CLK(clknet_8_112_0_clk),
    .RESET_B(net2073),
    .D(_02082_),
    .Q_N(_12097_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[16] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[17]$_DFFE_PP_  (.CLK(clknet_leaf_382_clk),
    .RESET_B(net2074),
    .D(_02083_),
    .Q_N(_12096_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[17] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[18]$_DFFE_PP_  (.CLK(clknet_leaf_379_clk),
    .RESET_B(net2075),
    .D(_02084_),
    .Q_N(_12095_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[18] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[19]$_DFFE_PP_  (.CLK(clknet_leaf_382_clk),
    .RESET_B(net2076),
    .D(_02085_),
    .Q_N(_12094_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[19] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_412_clk),
    .RESET_B(net2077),
    .D(_02086_),
    .Q_N(_12093_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[20]$_DFFE_PP_  (.CLK(clknet_leaf_377_clk),
    .RESET_B(net2078),
    .D(_02087_),
    .Q_N(_12092_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[20] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[21]$_DFFE_PP_  (.CLK(clknet_leaf_394_clk),
    .RESET_B(net2079),
    .D(_02088_),
    .Q_N(_12091_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[21] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[22]$_DFFE_PP_  (.CLK(clknet_leaf_379_clk),
    .RESET_B(net2080),
    .D(_02089_),
    .Q_N(_12090_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[22] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[23]$_DFFE_PP_  (.CLK(clknet_leaf_382_clk),
    .RESET_B(net2081),
    .D(_02090_),
    .Q_N(_12089_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[23] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[24]$_DFFE_PP_  (.CLK(clknet_leaf_414_clk),
    .RESET_B(net2082),
    .D(_02091_),
    .Q_N(_12088_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[24] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[25]$_DFFE_PP_  (.CLK(clknet_leaf_394_clk),
    .RESET_B(net2083),
    .D(_02092_),
    .Q_N(_12087_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[25] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[26]$_DFFE_PP_  (.CLK(clknet_leaf_398_clk),
    .RESET_B(net2084),
    .D(_02093_),
    .Q_N(_12086_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[26] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[27]$_DFFE_PP_  (.CLK(clknet_leaf_378_clk),
    .RESET_B(net2085),
    .D(_02094_),
    .Q_N(_12085_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[27] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[28]$_DFFE_PP_  (.CLK(clknet_leaf_398_clk),
    .RESET_B(net2086),
    .D(_02095_),
    .Q_N(_12084_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[28] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[29]$_DFFE_PP_  (.CLK(clknet_leaf_394_clk),
    .RESET_B(net2087),
    .D(_02096_),
    .Q_N(_12083_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[29] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2088),
    .D(_02097_),
    .Q_N(_12082_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[30]$_DFFE_PP_  (.CLK(clknet_leaf_399_clk),
    .RESET_B(net2089),
    .D(_02098_),
    .Q_N(_12081_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[30] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[31]$_DFFE_PP_  (.CLK(clknet_leaf_377_clk),
    .RESET_B(net2090),
    .D(_02099_),
    .Q_N(_00127_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[31] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2091),
    .D(_02100_),
    .Q_N(_12080_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_406_clk),
    .RESET_B(net2092),
    .D(_02101_),
    .Q_N(_12079_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_404_clk),
    .RESET_B(net2093),
    .D(_02102_),
    .Q_N(_12078_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2094),
    .D(_02103_),
    .Q_N(_12077_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_403_clk),
    .RESET_B(net2095),
    .D(_02104_),
    .Q_N(_00126_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_407_clk),
    .RESET_B(net2096),
    .D(_02105_),
    .Q_N(_12076_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_408_clk),
    .RESET_B(net2097),
    .D(_02106_),
    .Q_N(_12075_),
    .Q(\u_ac_controller_soc_inst.spi_flash_rdata[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.softreset$_SDFF_PN1_  (.CLK(clknet_8_73_0_clk),
    .RESET_B(net2098),
    .D(_02107_),
    .Q_N(_14096_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.softreset ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[0]$_DFF_P_  (.CLK(clknet_8_77_0_clk),
    .RESET_B(net2099),
    .D(_00020_),
    .Q_N(_14097_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[10]$_DFF_P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2100),
    .D(_00021_),
    .Q_N(_14098_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[10] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[11]$_DFF_P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2101),
    .D(_00022_),
    .Q_N(_14099_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[11] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[12]$_DFF_P_  (.CLK(clknet_8_76_0_clk),
    .RESET_B(net2102),
    .D(_00023_),
    .Q_N(_14100_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[12] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[1]$_DFF_P_  (.CLK(clknet_8_76_0_clk),
    .RESET_B(net2103),
    .D(_00024_),
    .Q_N(_14101_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[2]$_DFF_P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2104),
    .D(_00025_),
    .Q_N(_14102_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[3]$_DFF_P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2105),
    .D(_00026_),
    .Q_N(_00100_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[4]$_DFF_P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2106),
    .D(_00027_),
    .Q_N(_14103_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[5]$_DFF_P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2107),
    .D(_00028_),
    .Q_N(_14104_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[6]$_DFF_P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2108),
    .D(_00029_),
    .Q_N(_14105_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[7]$_DFF_P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2109),
    .D(_00030_),
    .Q_N(_14106_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[8]$_DFF_P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2110),
    .D(_00031_),
    .Q_N(_14107_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[8] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.state[9]$_DFF_P_  (.CLK(clknet_8_76_0_clk),
    .RESET_B(net2111),
    .D(_00032_),
    .Q_N(_00099_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.state[9] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2112),
    .D(_02108_),
    .Q_N(_00094_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2113),
    .D(_02109_),
    .Q_N(_00091_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2114),
    .D(_02110_),
    .Q_N(_00093_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[3]$_SDFFE_PN0P_  (.CLK(clknet_8_68_0_clk),
    .RESET_B(net2115),
    .D(_02111_),
    .Q_N(_00092_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[0]$_SDFFE_PN0N_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2116),
    .D(_02112_),
    .Q_N(_12074_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[1]$_SDFFE_PN0N_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2117),
    .D(_02113_),
    .Q_N(_12073_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[2]$_SDFFE_PN0N_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2118),
    .D(_02114_),
    .Q_N(_12072_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[3]$_SDFFE_PN0N_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2119),
    .D(_02115_),
    .Q_N(_12071_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.fetch$_SDFF_PN1_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2120),
    .D(_02116_),
    .Q_N(_12070_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.fetch ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk$_SDFFE_PP0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2121),
    .D(_02117_),
    .Q_N(_00090_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_csb$_SDFFE_PN1P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2122),
    .D(_02118_),
    .Q_N(_12069_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_csb ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[0]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2123),
    .D(_02119_),
    .Q_N(_12068_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[1]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2124),
    .D(_02120_),
    .Q_N(_12067_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[2]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2125),
    .D(_02121_),
    .Q_N(_12066_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[3]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2126),
    .D(_02122_),
    .Q_N(_12065_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[4]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2127),
    .D(_02123_),
    .Q_N(_12064_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[5]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2128),
    .D(_02124_),
    .Q_N(_12063_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[6]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2129),
    .D(_02125_),
    .Q_N(_12062_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[7]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2130),
    .D(_02126_),
    .Q_N(_12061_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_data[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.last_fetch$_SDFF_PN1_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2131),
    .D(_02127_),
    .Q_N(_12060_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.last_fetch ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2132),
    .D(_02128_),
    .Q_N(_12059_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[1]$_DFFE_PP_  (.CLK(clknet_8_71_0_clk),
    .RESET_B(net2133),
    .D(_02129_),
    .Q_N(_12058_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[2]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2134),
    .D(_02130_),
    .Q_N(_12057_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2135),
    .D(_02131_),
    .Q_N(_12056_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[3] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[4]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2136),
    .D(_02132_),
    .Q_N(_12055_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[4] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[5]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2137),
    .D(_02133_),
    .Q_N(_12054_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[5] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[6]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2138),
    .D(_02134_),
    .Q_N(_12053_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[6] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[7]$_DFFE_PP_  (.CLK(clknet_8_69_0_clk),
    .RESET_B(net2139),
    .D(_02135_),
    .Q_N(_00124_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[7] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr$_SDFFE_PN0P_  (.CLK(clknet_8_70_0_clk),
    .RESET_B(net2140),
    .D(_02136_),
    .Q_N(_14108_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr_q$_DFF_P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2141),
    .D(net10466),
    .Q_N(_12052_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr_q ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2142),
    .D(_02137_),
    .Q_N(_12051_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_qspi$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2143),
    .D(_02138_),
    .Q_N(_12050_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_qspi ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_rd$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2144),
    .D(_02139_),
    .Q_N(_12049_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_rd ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2145),
    .D(_02140_),
    .Q_N(_12048_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2146),
    .D(_02141_),
    .Q_N(_12047_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2147),
    .D(_02142_),
    .Q_N(_14109_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag_q[0]$_DFF_P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2148),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[0] ),
    .Q_N(_14110_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[0] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag_q[1]$_DFF_P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2149),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[1] ),
    .Q_N(_14111_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[1] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag_q[2]$_DFF_P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2150),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[2] ),
    .Q_N(_12046_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.dout_tag[2] ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io0_90$_DFF_N_  (.CLK(net11061),
    .RESET_B(net2151),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io0_do ),
    .Q_N(_12045_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io0_90 ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io1_90$_DFF_N_  (.CLK(net11060),
    .RESET_B(net2152),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io1_do ),
    .Q_N(_12044_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io1_90 ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io2_90$_DFF_N_  (.CLK(net11059),
    .RESET_B(net2153),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io2_do ),
    .Q_N(_12043_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io2_90 ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io3_90$_DFF_N_  (.CLK(net11058),
    .RESET_B(net2154),
    .D(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_io3_do ),
    .Q_N(_12042_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io3_90 ));
 sg13g2_dfrbp_1 \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_resetn$_SDFF_PP0_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2155),
    .D(_02143_),
    .Q_N(_00095_),
    .Q(\u_ac_controller_soc_inst.u_spi_flash_mem.xfer.resetn ));
 sg13g2_IOPadVdd sg13g2_IOPadVdd_north_0 ();
 sg13g2_IOPadVss sg13g2_IOPadVss_north_1 ();
 sg13g2_IOPadOut16mA sg13g2_IOPadInOut16mA_x1 ();
 sg13g2_IOPadOut16mA sg13g2_IOPadOut16mA_x2 ();
 sg13g2_IOPadOut16mA sg13g2_IOPadOut16mA_x3 ();
 sg13g2_IOPadVdd sg13g2_IOPadVdd_south_0 ();
 sg13g2_IOPadVss sg13g2_IOPadVss_south_1 ();
 sg13g2_Corner IO_CORNER_NORTH_WEST_INST ();
 sg13g2_Corner IO_CORNER_NORTH_EAST_INST ();
 sg13g2_Corner IO_CORNER_SOUTH_WEST_INST ();
 sg13g2_Corner IO_CORNER_SOUTH_EAST_INST ();
 sg13g2_Filler4000 IO_FILL_IO_NORTH_0_0 ();
 sg13g2_Filler2000 IO_FILL_IO_NORTH_0_20 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_0_30 ();
 sg13g2_Filler10000 IO_FILL_IO_NORTH_1_0 ();
 sg13g2_Filler2000 IO_FILL_IO_NORTH_1_50 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_1_60 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_62 ();
 sg13g2_Filler10000 IO_FILL_IO_NORTH_2_0 ();
 sg13g2_Filler2000 IO_FILL_IO_NORTH_2_50 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_2_60 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_62 ();
 sg13g2_Filler10000 IO_FILL_IO_NORTH_3_0 ();
 sg13g2_Filler2000 IO_FILL_IO_NORTH_3_50 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_3_60 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_3_62 ();
 sg13g2_Filler10000 IO_FILL_IO_NORTH_4_0 ();
 sg13g2_Filler2000 IO_FILL_IO_NORTH_4_50 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_4_60 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_62 ();
 sg13g2_Filler10000 IO_FILL_IO_NORTH_5_0 ();
 sg13g2_Filler2000 IO_FILL_IO_NORTH_5_50 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_5_60 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_62 ();
 sg13g2_Filler4000 IO_FILL_IO_NORTH_6_0 ();
 sg13g2_Filler2000 IO_FILL_IO_NORTH_6_20 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_6_30 ();
 sg13g2_Filler4000 IO_FILL_IO_SOUTH_0_0 ();
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_0_20 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_0_30 ();
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_1_0 ();
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_1_50 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_1_60 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_62 ();
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_2_0 ();
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_2_50 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_2_60 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_62 ();
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_3_0 ();
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_3_50 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_3_60 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_3_62 ();
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_4_0 ();
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_4_50 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_4_60 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_62 ();
 sg13g2_Filler10000 IO_FILL_IO_SOUTH_5_0 ();
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_5_50 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_5_60 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_62 ();
 sg13g2_Filler4000 IO_FILL_IO_SOUTH_6_0 ();
 sg13g2_Filler2000 IO_FILL_IO_SOUTH_6_20 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_6_30 ();
 sg13g2_Filler4000 IO_FILL_IO_WEST_0_0 ();
 sg13g2_Filler2000 IO_FILL_IO_WEST_0_20 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_0_30 ();
 sg13g2_Filler10000 IO_FILL_IO_WEST_1_0 ();
 sg13g2_Filler2000 IO_FILL_IO_WEST_1_50 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_1_60 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_62 ();
 sg13g2_Filler10000 IO_FILL_IO_WEST_2_0 ();
 sg13g2_Filler2000 IO_FILL_IO_WEST_2_50 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_2_60 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_62 ();
 sg13g2_Filler10000 IO_FILL_IO_WEST_3_0 ();
 sg13g2_Filler2000 IO_FILL_IO_WEST_3_50 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_3_60 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_3_62 ();
 sg13g2_Filler10000 IO_FILL_IO_WEST_4_0 ();
 sg13g2_Filler2000 IO_FILL_IO_WEST_4_50 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_4_60 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_62 ();
 sg13g2_Filler10000 IO_FILL_IO_WEST_5_0 ();
 sg13g2_Filler2000 IO_FILL_IO_WEST_5_50 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_5_60 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_62 ();
 sg13g2_Filler4000 IO_FILL_IO_WEST_6_0 ();
 sg13g2_Filler2000 IO_FILL_IO_WEST_6_20 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_6_30 ();
 sg13g2_Filler4000 IO_FILL_IO_EAST_0_0 ();
 sg13g2_Filler2000 IO_FILL_IO_EAST_0_20 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_0_30 ();
 sg13g2_Filler10000 IO_FILL_IO_EAST_1_0 ();
 sg13g2_Filler2000 IO_FILL_IO_EAST_1_50 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_1_60 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_62 ();
 sg13g2_Filler10000 IO_FILL_IO_EAST_2_0 ();
 sg13g2_Filler2000 IO_FILL_IO_EAST_2_50 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_2_60 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_62 ();
 sg13g2_Filler10000 IO_FILL_IO_EAST_3_0 ();
 sg13g2_Filler2000 IO_FILL_IO_EAST_3_50 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_3_60 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_3_62 ();
 sg13g2_Filler10000 IO_FILL_IO_EAST_4_0 ();
 sg13g2_Filler2000 IO_FILL_IO_EAST_4_50 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_4_60 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_62 ();
 sg13g2_Filler10000 IO_FILL_IO_EAST_5_0 ();
 sg13g2_Filler2000 IO_FILL_IO_EAST_5_50 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_5_60 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_62 ();
 sg13g2_Filler4000 IO_FILL_IO_EAST_6_0 ();
 sg13g2_Filler2000 IO_FILL_IO_EAST_6_20 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_6_30 ();
 bondpad_70x70 IO_BOND_sg13g2_IOPadInOut16mA_gpio_1_pad_inst (.pad(gpio_1_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadInOut16mA_gpio_2_pad_inst (.pad(gpio_2_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadInOut16mA_spi_flash_io0_pad_inst (.pad(spi_flash_io0_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadInOut16mA_spi_flash_io1_pad_inst (.pad(spi_flash_io1_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadInOut16mA_spi_flash_io2_pad_inst (.pad(spi_flash_io2_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadInOut16mA_spi_flash_io3_pad_inst (.pad(spi_flash_io3_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadIn_clk_pad_inst (.pad(clk_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadIn_resetn_pad_inst (.pad(resetn_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadIn_ser_rx_pad_inst (.pad(ser_rx_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadIn_spi_sensor_miso_pad_inst (.pad(spi_sensor_miso_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadOut16mA_pwm_out_pad_inst (.pad(pwm_out_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadOut16mA_ser_tx_pad_inst (.pad(ser_tx_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadOut16mA_spi_flash_clk_pad_inst (.pad(spi_flash_clk_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadOut16mA_spi_flash_cs_n_pad_inst (.pad(spi_flash_cs_n_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadOut16mA_spi_sensor_clk_pad_inst (.pad(spi_sensor_clk_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadOut16mA_spi_sensor_cs_n_pad_inst (.pad(spi_sensor_cs_n_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadOut16mA_spi_sensor_mosi_pad_inst (.pad(spi_sensor_mosi_pad));
 bondpad_70x70 IO_BOND_sg13g2_IOPadVdd_north_0 (.pad(\IO_CORNER_NORTH_WEST_INST.vdd_RING ));
 bondpad_70x70 IO_BOND_sg13g2_IOPadVss_north_1 (.pad(\IO_CORNER_NORTH_WEST_INST.vss_RING ));
 bondpad_70x70 IO_BOND_sg13g2_IOPadInOut16mA_x1 ();
 bondpad_70x70 IO_BOND_sg13g2_IOPadOut16mA_x2 ();
 bondpad_70x70 IO_BOND_sg13g2_IOPadOut16mA_x3 ();
 bondpad_70x70 IO_BOND_sg13g2_IOPadVdd_south_0 (.pad(\IO_CORNER_NORTH_WEST_INST.vdd_RING ));
 bondpad_70x70 IO_BOND_sg13g2_IOPadVss_south_1 (.pad(\IO_CORNER_NORTH_WEST_INST.vss_RING ));
 sg13g2_tiehi _26132__1 (.L_HI(net1));
 sg13g2_tiehi _26133__2 (.L_HI(net2));
 sg13g2_tiehi _26134__3 (.L_HI(net3));
 sg13g2_tiehi _26135__4 (.L_HI(net4));
 sg13g2_tiehi _26136__5 (.L_HI(net5));
 sg13g2_tiehi _26137__6 (.L_HI(net6));
 sg13g2_tiehi _26138__7 (.L_HI(net7));
 sg13g2_tiehi _26139__8 (.L_HI(net8));
 sg13g2_tiehi _26140__9 (.L_HI(net9));
 sg13g2_tiehi _26141__10 (.L_HI(net10));
 sg13g2_tiehi \u_ac_controller_soc_inst.sram_wrapper_inst.ready_state$_SDFF_PP0__11  (.L_HI(net11));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[0]$_SDFF_PP0__12  (.L_HI(net12));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[10]$_SDFF_PP0__13  (.L_HI(net13));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[11]$_SDFF_PP0__14  (.L_HI(net14));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[12]$_SDFF_PP0__15  (.L_HI(net15));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[13]$_SDFF_PP0__16  (.L_HI(net16));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[14]$_SDFF_PP0__17  (.L_HI(net17));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[15]$_SDFF_PP0__18  (.L_HI(net18));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[16]$_SDFF_PP0__19  (.L_HI(net19));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[17]$_SDFF_PP0__20  (.L_HI(net20));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[18]$_SDFF_PP0__21  (.L_HI(net21));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[19]$_SDFF_PP0__22  (.L_HI(net22));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[1]$_SDFF_PP0__23  (.L_HI(net23));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[20]$_SDFF_PP0__24  (.L_HI(net24));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[21]$_SDFF_PP0__25  (.L_HI(net25));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[22]$_SDFF_PP0__26  (.L_HI(net26));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[23]$_SDFF_PP0__27  (.L_HI(net27));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[24]$_SDFF_PP0__28  (.L_HI(net28));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[25]$_SDFF_PP0__29  (.L_HI(net29));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[26]$_SDFF_PP0__30  (.L_HI(net30));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[27]$_SDFF_PP0__31  (.L_HI(net31));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[28]$_SDFF_PP0__32  (.L_HI(net32));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[29]$_SDFF_PP0__33  (.L_HI(net33));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[2]$_SDFF_PP0__34  (.L_HI(net34));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[30]$_SDFF_PP0__35  (.L_HI(net35));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[31]$_SDFF_PP0__36  (.L_HI(net36));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[3]$_SDFF_PP0__37  (.L_HI(net37));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[4]$_SDFF_PP0__38  (.L_HI(net38));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[5]$_SDFF_PP0__39  (.L_HI(net39));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[6]$_SDFF_PP0__40  (.L_HI(net40));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[7]$_SDFF_PP0__41  (.L_HI(net41));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[8]$_SDFF_PP0__42  (.L_HI(net42));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.counter[9]$_SDFF_PP0__43  (.L_HI(net43));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[0]$_SDFFE_PN0P__44  (.L_HI(net44));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[10]$_SDFFE_PN0P__45  (.L_HI(net45));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[11]$_SDFFE_PN0P__46  (.L_HI(net46));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[12]$_SDFFE_PN0P__47  (.L_HI(net47));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[13]$_SDFFE_PN0P__48  (.L_HI(net48));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[14]$_SDFFE_PN0P__49  (.L_HI(net49));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[15]$_SDFFE_PN0P__50  (.L_HI(net50));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[16]$_SDFFE_PN0P__51  (.L_HI(net51));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[17]$_SDFFE_PN0P__52  (.L_HI(net52));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[18]$_SDFFE_PN0P__53  (.L_HI(net53));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[19]$_SDFFE_PN0P__54  (.L_HI(net54));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[1]$_SDFFE_PN0P__55  (.L_HI(net55));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[20]$_SDFFE_PN0P__56  (.L_HI(net56));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[21]$_SDFFE_PN0P__57  (.L_HI(net57));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[22]$_SDFFE_PN0P__58  (.L_HI(net58));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[23]$_SDFFE_PN0P__59  (.L_HI(net59));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[24]$_SDFFE_PN0P__60  (.L_HI(net60));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[25]$_SDFFE_PN0P__61  (.L_HI(net61));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[26]$_SDFFE_PN0P__62  (.L_HI(net62));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[27]$_SDFFE_PN0P__63  (.L_HI(net63));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[28]$_SDFFE_PN0P__64  (.L_HI(net64));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[29]$_SDFFE_PN0P__65  (.L_HI(net65));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[2]$_SDFFE_PN0P__66  (.L_HI(net66));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[30]$_SDFFE_PN0P__67  (.L_HI(net67));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[31]$_SDFFE_PN0P__68  (.L_HI(net68));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[3]$_SDFFE_PN0P__69  (.L_HI(net69));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[4]$_SDFFE_PN0P__70  (.L_HI(net70));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[5]$_SDFFE_PN0P__71  (.L_HI(net71));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[6]$_SDFFE_PN0P__72  (.L_HI(net72));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[7]$_SDFFE_PN0P__73  (.L_HI(net73));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[8]$_SDFFE_PN0P__74  (.L_HI(net74));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.device_address_reg[9]$_SDFFE_PN0P__75  (.L_HI(net75));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in1_sync1$_SDFF_PN0__76  (.L_HI(net76));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in1_sync2$_SDFF_PN0__77  (.L_HI(net77));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in2_sync1$_SDFF_PN0__78  (.L_HI(net78));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_in2_sync2$_SDFF_PN0__79  (.L_HI(net79));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_io1_oe$_SDFFE_PN0P__80  (.L_HI(net80));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_io2_oe$_SDFFE_PN0P__81  (.L_HI(net81));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_out1$_SDFFE_PN0P__82  (.L_HI(net82));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.gpio_out2$_SDFFE_PN0P__83  (.L_HI(net83));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[0]$_SDFFE_PN0P__84  (.L_HI(net84));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[10]$_SDFFE_PN0P__85  (.L_HI(net85));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[11]$_SDFFE_PN0P__86  (.L_HI(net86));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[12]$_SDFFE_PN0P__87  (.L_HI(net87));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[13]$_SDFFE_PN0P__88  (.L_HI(net88));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[14]$_SDFFE_PN0P__89  (.L_HI(net89));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[15]$_SDFFE_PN0P__90  (.L_HI(net90));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[16]$_SDFFE_PN0P__91  (.L_HI(net91));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[17]$_SDFFE_PN0P__92  (.L_HI(net92));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[18]$_SDFFE_PN0P__93  (.L_HI(net93));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[19]$_SDFFE_PN0P__94  (.L_HI(net94));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[1]$_SDFFE_PN0P__95  (.L_HI(net95));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[20]$_SDFFE_PN0P__96  (.L_HI(net96));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[21]$_SDFFE_PN0P__97  (.L_HI(net97));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[22]$_SDFFE_PN0P__98  (.L_HI(net98));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[23]$_SDFFE_PN0P__99  (.L_HI(net99));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[24]$_SDFFE_PN0P__100  (.L_HI(net100));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[25]$_SDFFE_PN0P__101  (.L_HI(net101));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[26]$_SDFFE_PN0P__102  (.L_HI(net102));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[27]$_SDFFE_PN0P__103  (.L_HI(net103));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[28]$_SDFFE_PN0P__104  (.L_HI(net104));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[29]$_SDFFE_PN0P__105  (.L_HI(net105));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[2]$_SDFFE_PN0P__106  (.L_HI(net106));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[30]$_SDFFE_PN0P__107  (.L_HI(net107));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[31]$_SDFFE_PN0P__108  (.L_HI(net108));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[3]$_SDFFE_PN0P__109  (.L_HI(net109));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[4]$_SDFFE_PN0P__110  (.L_HI(net110));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[5]$_SDFFE_PN0P__111  (.L_HI(net111));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[6]$_SDFFE_PN0P__112  (.L_HI(net112));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[7]$_SDFFE_PN0P__113  (.L_HI(net113));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[8]$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_rdata[9]$_SDFFE_PN0P__115  (.L_HI(net115));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.io_ready$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[0]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[10]$_SDFFE_PN0P__118  (.L_HI(net118));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[11]$_SDFFE_PN0P__119  (.L_HI(net119));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[12]$_SDFFE_PN0P__120  (.L_HI(net120));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[13]$_SDFFE_PN0P__121  (.L_HI(net121));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[14]$_SDFFE_PN0P__122  (.L_HI(net122));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[15]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[16]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[17]$_SDFFE_PN0P__125  (.L_HI(net125));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[18]$_SDFFE_PN0P__126  (.L_HI(net126));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[19]$_SDFFE_PN0P__127  (.L_HI(net127));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[1]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[20]$_SDFFE_PN0P__129  (.L_HI(net129));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[21]$_SDFFE_PN0P__130  (.L_HI(net130));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[22]$_SDFFE_PN0P__131  (.L_HI(net131));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[23]$_SDFFE_PN0P__132  (.L_HI(net132));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[24]$_SDFFE_PN0P__133  (.L_HI(net133));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[25]$_SDFFE_PN0P__134  (.L_HI(net134));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[26]$_SDFFE_PN0P__135  (.L_HI(net135));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[27]$_SDFFE_PN0P__136  (.L_HI(net136));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[28]$_SDFFE_PN0P__137  (.L_HI(net137));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[29]$_SDFFE_PN0P__138  (.L_HI(net138));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[2]$_SDFFE_PN0P__139  (.L_HI(net139));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[30]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[31]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[3]$_SDFFE_PN0P__142  (.L_HI(net142));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[4]$_SDFFE_PN0P__143  (.L_HI(net143));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[5]$_SDFFE_PN0P__144  (.L_HI(net144));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[6]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[7]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[8]$_SDFFE_PN0P__147  (.L_HI(net147));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_duty[9]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_enable$_SDFFE_PN1P__149  (.L_HI(net149));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_out$_SDFF_PN0__150  (.L_HI(net150));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[0]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[10]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[11]$_SDFFE_PN0P__153  (.L_HI(net153));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[12]$_SDFFE_PN0P__154  (.L_HI(net154));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[13]$_SDFFE_PN0P__155  (.L_HI(net155));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[14]$_SDFFE_PN0P__156  (.L_HI(net156));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[15]$_SDFFE_PN0P__157  (.L_HI(net157));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[16]$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[17]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[18]$_SDFFE_PN0P__160  (.L_HI(net160));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[19]$_SDFFE_PN0P__161  (.L_HI(net161));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[1]$_SDFFE_PN0P__162  (.L_HI(net162));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[20]$_SDFFE_PN0P__163  (.L_HI(net163));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[21]$_SDFFE_PN0P__164  (.L_HI(net164));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[22]$_SDFFE_PN0P__165  (.L_HI(net165));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[23]$_SDFFE_PN0P__166  (.L_HI(net166));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[24]$_SDFFE_PN0P__167  (.L_HI(net167));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[25]$_SDFFE_PN0P__168  (.L_HI(net168));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[26]$_SDFFE_PN0P__169  (.L_HI(net169));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[27]$_SDFFE_PN0P__170  (.L_HI(net170));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[28]$_SDFFE_PN0P__171  (.L_HI(net171));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[29]$_SDFFE_PN0P__172  (.L_HI(net172));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[2]$_SDFFE_PN0P__173  (.L_HI(net173));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[30]$_SDFFE_PN0P__174  (.L_HI(net174));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[31]$_SDFFE_PN0P__175  (.L_HI(net175));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[3]$_SDFFE_PN0P__176  (.L_HI(net176));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[4]$_SDFFE_PN0P__177  (.L_HI(net177));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[5]$_SDFFE_PN0P__178  (.L_HI(net178));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[6]$_SDFFE_PN0P__179  (.L_HI(net179));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[7]$_SDFFE_PN0P__180  (.L_HI(net180));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[8]$_SDFFE_PN0P__181  (.L_HI(net181));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_io_controller_bridge.pwm_period[9]$_SDFFE_PN0P__182  (.L_HI(net182));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[0]$_SDFFE_PN0P__183  (.L_HI(net183));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[1]$_SDFFE_PN0P__184  (.L_HI(net184));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[2]$_SDFFE_PN0P__185  (.L_HI(net185));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[3]$_SDFFE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[4]$_SDFFE_PN0P__187  (.L_HI(net187));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.current_bit_count[5]$_SDFFE_PN0P__188  (.L_HI(net188));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[0]$_SDFFE_PN0P__189  (.L_HI(net189));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[10]$_SDFFE_PN0P__190  (.L_HI(net190));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[11]$_SDFFE_PN0P__191  (.L_HI(net191));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[12]$_SDFFE_PN0P__192  (.L_HI(net192));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[13]$_SDFFE_PN0P__193  (.L_HI(net193));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[14]$_SDFFE_PN0P__194  (.L_HI(net194));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[15]$_SDFFE_PN0P__195  (.L_HI(net195));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[16]$_SDFFE_PN0P__196  (.L_HI(net196));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[17]$_SDFFE_PN0P__197  (.L_HI(net197));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[18]$_SDFFE_PN0P__198  (.L_HI(net198));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[19]$_SDFFE_PN0P__199  (.L_HI(net199));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[1]$_SDFFE_PN0P__200  (.L_HI(net200));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[20]$_SDFFE_PN0P__201  (.L_HI(net201));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[21]$_SDFFE_PN0P__202  (.L_HI(net202));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[22]$_SDFFE_PN0P__203  (.L_HI(net203));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[23]$_SDFFE_PN0P__204  (.L_HI(net204));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[24]$_SDFFE_PN0P__205  (.L_HI(net205));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[25]$_SDFFE_PN0P__206  (.L_HI(net206));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[26]$_SDFFE_PN0P__207  (.L_HI(net207));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[27]$_SDFFE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[28]$_SDFFE_PN0P__209  (.L_HI(net209));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[29]$_SDFFE_PN0P__210  (.L_HI(net210));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[2]$_SDFFE_PN0P__211  (.L_HI(net211));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[30]$_SDFFE_PN0P__212  (.L_HI(net212));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[31]$_SDFFE_PN0P__213  (.L_HI(net213));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[3]$_SDFFE_PN0P__214  (.L_HI(net214));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[4]$_SDFFE_PN0P__215  (.L_HI(net215));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[5]$_SDFFE_PN0P__216  (.L_HI(net216));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[6]$_SDFFE_PN0P__217  (.L_HI(net217));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[7]$_SDFFE_PN0P__218  (.L_HI(net218));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[8]$_SDFFE_PN0P__219  (.L_HI(net219));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_capture[9]$_SDFFE_PN0P__220  (.L_HI(net220));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[0]$_SDFFE_PN0P__221  (.L_HI(net221));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[10]$_SDFFE_PN0P__222  (.L_HI(net222));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[11]$_SDFFE_PN0P__223  (.L_HI(net223));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[12]$_SDFFE_PN0P__224  (.L_HI(net224));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[13]$_SDFFE_PN0P__225  (.L_HI(net225));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[14]$_SDFFE_PN0P__226  (.L_HI(net226));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[15]$_SDFFE_PN0P__227  (.L_HI(net227));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[16]$_SDFFE_PN0P__228  (.L_HI(net228));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[17]$_SDFFE_PN0P__229  (.L_HI(net229));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[18]$_SDFFE_PN0P__230  (.L_HI(net230));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[19]$_SDFFE_PN0P__231  (.L_HI(net231));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[1]$_SDFFE_PN0P__232  (.L_HI(net232));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[20]$_SDFFE_PN0P__233  (.L_HI(net233));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[21]$_SDFFE_PN0P__234  (.L_HI(net234));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[22]$_SDFFE_PN0P__235  (.L_HI(net235));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[23]$_SDFFE_PN0P__236  (.L_HI(net236));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[24]$_SDFFE_PN0P__237  (.L_HI(net237));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[25]$_SDFFE_PN0P__238  (.L_HI(net238));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[26]$_SDFFE_PN0P__239  (.L_HI(net239));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[27]$_SDFFE_PN0P__240  (.L_HI(net240));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[28]$_SDFFE_PN0P__241  (.L_HI(net241));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[29]$_SDFFE_PN0P__242  (.L_HI(net242));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[2]$_SDFFE_PN0P__243  (.L_HI(net243));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[30]$_SDFFE_PN0P__244  (.L_HI(net244));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[31]$_SDFFE_PN0P__245  (.L_HI(net245));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[32]$_SDFFE_PN0P__246  (.L_HI(net246));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[33]$_SDFFE_PN0P__247  (.L_HI(net247));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[34]$_SDFFE_PP0P__248  (.L_HI(net248));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[35]$_SDFFE_PP0P__249  (.L_HI(net249));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[36]$_SDFFE_PN0P__250  (.L_HI(net250));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[37]$_SDFFE_PN0P__251  (.L_HI(net251));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[38]$_SDFFE_PN0P__252  (.L_HI(net252));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[39]$_SDFFE_PN0P__253  (.L_HI(net253));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[3]$_SDFFE_PN0P__254  (.L_HI(net254));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[4]$_SDFFE_PN0P__255  (.L_HI(net255));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[5]$_SDFFE_PN0P__256  (.L_HI(net256));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[6]$_SDFFE_PN0P__257  (.L_HI(net257));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[7]$_SDFFE_PN0P__258  (.L_HI(net258));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[8]$_SDFFE_PN0P__259  (.L_HI(net259));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.data_to_send[9]$_SDFFE_PN0P__260  (.L_HI(net260));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.spi_clk_reg$_SDFF_PN0__261  (.L_HI(net261));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.spi_cs_n_reg$_SDFFE_PP1P__262  (.L_HI(net262));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.spi_sensor_ready_reg$_SDFF_PN0__263  (.L_HI(net263));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[3]$_SDFF_PN0__264  (.L_HI(net264));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[4]$_SDFF_PN1__265  (.L_HI(net265));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_bit_count[5]$_SDFF_PN0__266  (.L_HI(net266));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[0]$_SDFFE_PN0P__267  (.L_HI(net267));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_spi_bridge.write_read_byte_count[1]$_SDFFE_PN0P__268  (.L_HI(net268));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[0]$_SDFFE_PP0P__269  (.L_HI(net269));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[1]$_SDFFE_PP0P__270  (.L_HI(net270));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_bit_count[2]$_SDFFE_PP0P__271  (.L_HI(net271));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[0]$_SDFFE_PP0P__272  (.L_HI(net272));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[10]$_SDFFE_PP0P__273  (.L_HI(net273));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[11]$_SDFFE_PP0P__274  (.L_HI(net274));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[12]$_SDFFE_PP0P__275  (.L_HI(net275));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[13]$_SDFFE_PP0P__276  (.L_HI(net276));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[14]$_SDFFE_PP0P__277  (.L_HI(net277));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[15]$_SDFFE_PP0P__278  (.L_HI(net278));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[16]$_SDFFE_PP0P__279  (.L_HI(net279));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[17]$_SDFFE_PP0P__280  (.L_HI(net280));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[18]$_SDFFE_PP0P__281  (.L_HI(net281));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[19]$_SDFFE_PP0P__282  (.L_HI(net282));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[1]$_SDFFE_PP0P__283  (.L_HI(net283));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[20]$_SDFFE_PP0P__284  (.L_HI(net284));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[21]$_SDFFE_PP0P__285  (.L_HI(net285));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[22]$_SDFFE_PP0P__286  (.L_HI(net286));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[23]$_SDFFE_PP0P__287  (.L_HI(net287));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[24]$_SDFFE_PP0P__288  (.L_HI(net288));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[25]$_SDFFE_PP0P__289  (.L_HI(net289));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[26]$_SDFFE_PP0P__290  (.L_HI(net290));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[27]$_SDFFE_PP0P__291  (.L_HI(net291));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[28]$_SDFFE_PP0P__292  (.L_HI(net292));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[29]$_SDFFE_PP0P__293  (.L_HI(net293));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[2]$_SDFFE_PP0P__294  (.L_HI(net294));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[30]$_SDFFE_PP0P__295  (.L_HI(net295));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[31]$_SDFFE_PP0P__296  (.L_HI(net296));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[3]$_SDFFE_PP0P__297  (.L_HI(net297));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[4]$_SDFFE_PP0P__298  (.L_HI(net298));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[5]$_SDFFE_PP0P__299  (.L_HI(net299));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[6]$_SDFFE_PP0P__300  (.L_HI(net300));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[7]$_SDFFE_PP0P__301  (.L_HI(net301));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[8]$_SDFFE_PP0P__302  (.L_HI(net302));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.actual_clk_div_count[9]$_SDFFE_PP0P__303  (.L_HI(net303));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[0]$_SDFFE_PN0P__304  (.L_HI(net304));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[1]$_SDFFE_PN0P__305  (.L_HI(net305));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[2]$_SDFFE_PN0P__306  (.L_HI(net306));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[3]$_SDFFE_PN0P__307  (.L_HI(net307));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[4]$_SDFFE_PN0P__308  (.L_HI(net308));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[5]$_SDFFE_PN0P__309  (.L_HI(net309));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[6]$_SDFFE_PN0P__310  (.L_HI(net310));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[7]$_SDFFE_PN0P__311  (.L_HI(net311));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.received_data[8]$_SDFFE_PN0P__312  (.L_HI(net312));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync1$_SDFF_PN1__313  (.L_HI(net313));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_rx_sync2$_SDFF_PN1__314  (.L_HI(net314));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.ser_tx$_SDFFE_PP1P__315  (.L_HI(net315));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.start_bit$_SDFFE_PP0P__316  (.L_HI(net316));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.stop_bit$_SDFFE_PP0P__317  (.L_HI(net317));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[0]$_SDFFE_PN0P__318  (.L_HI(net318));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[1]$_SDFFE_PN0P__319  (.L_HI(net319));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[2]$_SDFFE_PN0P__320  (.L_HI(net320));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[3]$_SDFFE_PN0P__321  (.L_HI(net321));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[4]$_SDFFE_PN0P__322  (.L_HI(net322));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[5]$_SDFFE_PN0P__323  (.L_HI(net323));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[6]$_SDFFE_PN0P__324  (.L_HI(net324));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[7]$_SDFFE_PN0P__325  (.L_HI(net325));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_rdata[8]$_SDFFE_PN0P__326  (.L_HI(net326));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.uart_ready$_SDFF_PN0__327  (.L_HI(net327));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[0]$_SDFFE_PN0P__328  (.L_HI(net328));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[1]$_SDFFE_PN0P__329  (.L_HI(net329));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_bit_count[2]$_SDFFE_PN0P__330  (.L_HI(net330));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[0]$_SDFFE_PN0P__331  (.L_HI(net331));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[10]$_SDFFE_PN0P__332  (.L_HI(net332));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[11]$_SDFFE_PN0P__333  (.L_HI(net333));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[12]$_SDFFE_PN0P__334  (.L_HI(net334));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[13]$_SDFFE_PN0P__335  (.L_HI(net335));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[14]$_SDFFE_PN0P__336  (.L_HI(net336));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[15]$_SDFFE_PN0P__337  (.L_HI(net337));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[16]$_SDFFE_PN0P__338  (.L_HI(net338));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[17]$_SDFFE_PN0P__339  (.L_HI(net339));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[18]$_SDFFE_PN0P__340  (.L_HI(net340));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[19]$_SDFFE_PN0P__341  (.L_HI(net341));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[1]$_SDFFE_PN0P__342  (.L_HI(net342));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[20]$_SDFFE_PN0P__343  (.L_HI(net343));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[21]$_SDFFE_PN0P__344  (.L_HI(net344));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[22]$_SDFFE_PN0P__345  (.L_HI(net345));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[23]$_SDFFE_PN0P__346  (.L_HI(net346));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[24]$_SDFFE_PN0P__347  (.L_HI(net347));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[25]$_SDFFE_PN0P__348  (.L_HI(net348));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[26]$_SDFFE_PN0P__349  (.L_HI(net349));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[27]$_SDFFE_PN0P__350  (.L_HI(net350));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[28]$_SDFFE_PN0P__351  (.L_HI(net351));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[29]$_SDFFE_PN0P__352  (.L_HI(net352));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[2]$_SDFFE_PN0P__353  (.L_HI(net353));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[30]$_SDFFE_PN0P__354  (.L_HI(net354));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[31]$_SDFFE_PN0P__355  (.L_HI(net355));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[3]$_SDFFE_PN0P__356  (.L_HI(net356));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[4]$_SDFFE_PN0P__357  (.L_HI(net357));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[5]$_SDFFE_PN0P__358  (.L_HI(net358));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[6]$_SDFFE_PN0P__359  (.L_HI(net359));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[7]$_SDFFE_PN0P__360  (.L_HI(net360));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[8]$_SDFFE_PN0P__361  (.L_HI(net361));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_clk_div_count[9]$_SDFFE_PN0P__362  (.L_HI(net362));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_done$_SDFF_PN0__363  (.L_HI(net363));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout$_SDFF_PP0__364  (.L_HI(net364));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[0]$_SDFFE_PN0P__365  (.L_HI(net365));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[10]$_SDFFE_PN0P__366  (.L_HI(net366));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[11]$_SDFFE_PN0P__367  (.L_HI(net367));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[12]$_SDFFE_PN0P__368  (.L_HI(net368));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[13]$_SDFFE_PN0P__369  (.L_HI(net369));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[14]$_SDFFE_PN0P__370  (.L_HI(net370));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[15]$_SDFFE_PN0P__371  (.L_HI(net371));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[16]$_SDFFE_PN0P__372  (.L_HI(net372));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[17]$_SDFFE_PN0P__373  (.L_HI(net373));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[18]$_SDFFE_PN0P__374  (.L_HI(net374));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[19]$_SDFFE_PN0P__375  (.L_HI(net375));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[1]$_SDFFE_PN0P__376  (.L_HI(net376));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[20]$_SDFFE_PN0P__377  (.L_HI(net377));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[21]$_SDFFE_PN0P__378  (.L_HI(net378));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[22]$_SDFFE_PN0P__379  (.L_HI(net379));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[23]$_SDFFE_PN0P__380  (.L_HI(net380));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[24]$_SDFFE_PN0P__381  (.L_HI(net381));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[25]$_SDFFE_PN0P__382  (.L_HI(net382));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[26]$_SDFFE_PN0P__383  (.L_HI(net383));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[27]$_SDFFE_PN0P__384  (.L_HI(net384));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[28]$_SDFFE_PN0P__385  (.L_HI(net385));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[29]$_SDFFE_PN0P__386  (.L_HI(net386));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[2]$_SDFFE_PN0P__387  (.L_HI(net387));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[30]$_SDFFE_PN0P__388  (.L_HI(net388));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[31]$_SDFFE_PN0P__389  (.L_HI(net389));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[3]$_SDFFE_PN0P__390  (.L_HI(net390));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[4]$_SDFFE_PN0P__391  (.L_HI(net391));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[5]$_SDFFE_PN0P__392  (.L_HI(net392));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[6]$_SDFFE_PN0P__393  (.L_HI(net393));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[7]$_SDFFE_PN0P__394  (.L_HI(net394));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[8]$_SDFFE_PN0P__395  (.L_HI(net395));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfer_timeout_counter[9]$_SDFFE_PN0P__396  (.L_HI(net396));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_cbus_to_uart_bridge.xfering$_SDFFE_PN0P__397  (.L_HI(net397));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[0]$_DFF_P__398  (.L_HI(net398));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[10]$_DFF_P__399  (.L_HI(net399));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[11]$_DFF_P__400  (.L_HI(net400));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[12]$_DFF_P__401  (.L_HI(net401));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[13]$_DFF_P__402  (.L_HI(net402));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[14]$_DFF_P__403  (.L_HI(net403));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[15]$_DFF_P__404  (.L_HI(net404));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[16]$_DFF_P__405  (.L_HI(net405));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[17]$_DFF_P__406  (.L_HI(net406));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[18]$_DFF_P__407  (.L_HI(net407));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[19]$_DFF_P__408  (.L_HI(net408));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[1]$_DFF_P__409  (.L_HI(net409));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[20]$_DFF_P__410  (.L_HI(net410));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[21]$_DFF_P__411  (.L_HI(net411));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[22]$_DFF_P__412  (.L_HI(net412));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[23]$_DFF_P__413  (.L_HI(net413));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[24]$_DFF_P__414  (.L_HI(net414));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[25]$_DFF_P__415  (.L_HI(net415));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[26]$_DFF_P__416  (.L_HI(net416));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[27]$_DFF_P__417  (.L_HI(net417));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[28]$_DFF_P__418  (.L_HI(net418));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[29]$_DFF_P__419  (.L_HI(net419));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[2]$_DFF_P__420  (.L_HI(net420));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[30]$_DFF_P__421  (.L_HI(net421));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[31]$_DFF_P__422  (.L_HI(net422));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[3]$_DFF_P__423  (.L_HI(net423));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[4]$_DFF_P__424  (.L_HI(net424));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[5]$_DFF_P__425  (.L_HI(net425));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[6]$_DFF_P__426  (.L_HI(net426));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[7]$_DFF_P__427  (.L_HI(net427));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[8]$_DFF_P__428  (.L_HI(net428));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.alu_out_q[9]$_DFF_P__429  (.L_HI(net429));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[0]$_SDFF_PN0__430  (.L_HI(net430));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[10]$_SDFF_PN0__431  (.L_HI(net431));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[11]$_SDFF_PN0__432  (.L_HI(net432));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[12]$_SDFF_PN0__433  (.L_HI(net433));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[13]$_SDFF_PN0__434  (.L_HI(net434));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[14]$_SDFF_PN0__435  (.L_HI(net435));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[15]$_SDFF_PN0__436  (.L_HI(net436));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[16]$_SDFF_PN0__437  (.L_HI(net437));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[17]$_SDFF_PN0__438  (.L_HI(net438));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[18]$_SDFF_PN0__439  (.L_HI(net439));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[19]$_SDFF_PN0__440  (.L_HI(net440));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[1]$_SDFF_PN0__441  (.L_HI(net441));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[20]$_SDFF_PN0__442  (.L_HI(net442));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[21]$_SDFF_PN0__443  (.L_HI(net443));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[22]$_SDFF_PN0__444  (.L_HI(net444));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[23]$_SDFF_PN0__445  (.L_HI(net445));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[24]$_SDFF_PN0__446  (.L_HI(net446));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[25]$_SDFF_PN0__447  (.L_HI(net447));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[26]$_SDFF_PN0__448  (.L_HI(net448));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[27]$_SDFF_PN0__449  (.L_HI(net449));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[28]$_SDFF_PN0__450  (.L_HI(net450));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[29]$_SDFF_PN0__451  (.L_HI(net451));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[2]$_SDFF_PN0__452  (.L_HI(net452));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[30]$_SDFF_PN0__453  (.L_HI(net453));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[31]$_SDFF_PN0__454  (.L_HI(net454));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[32]$_SDFF_PN0__455  (.L_HI(net455));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[33]$_SDFF_PN0__456  (.L_HI(net456));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[34]$_SDFF_PN0__457  (.L_HI(net457));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[35]$_SDFF_PN0__458  (.L_HI(net458));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[36]$_SDFF_PN0__459  (.L_HI(net459));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[37]$_SDFF_PN0__460  (.L_HI(net460));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[38]$_SDFF_PN0__461  (.L_HI(net461));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[39]$_SDFF_PN0__462  (.L_HI(net462));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[3]$_SDFF_PN0__463  (.L_HI(net463));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[40]$_SDFF_PN0__464  (.L_HI(net464));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[41]$_SDFF_PN0__465  (.L_HI(net465));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[42]$_SDFF_PN0__466  (.L_HI(net466));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[43]$_SDFF_PN0__467  (.L_HI(net467));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[44]$_SDFF_PN0__468  (.L_HI(net468));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[45]$_SDFF_PN0__469  (.L_HI(net469));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[46]$_SDFF_PN0__470  (.L_HI(net470));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[47]$_SDFF_PN0__471  (.L_HI(net471));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[48]$_SDFF_PN0__472  (.L_HI(net472));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[49]$_SDFF_PN0__473  (.L_HI(net473));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[4]$_SDFF_PN0__474  (.L_HI(net474));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[50]$_SDFF_PN0__475  (.L_HI(net475));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[51]$_SDFF_PN0__476  (.L_HI(net476));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[52]$_SDFF_PN0__477  (.L_HI(net477));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[53]$_SDFF_PN0__478  (.L_HI(net478));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[54]$_SDFF_PN0__479  (.L_HI(net479));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[55]$_SDFF_PN0__480  (.L_HI(net480));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[56]$_SDFF_PN0__481  (.L_HI(net481));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[57]$_SDFF_PN0__482  (.L_HI(net482));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[58]$_SDFF_PN0__483  (.L_HI(net483));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[59]$_SDFF_PN0__484  (.L_HI(net484));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[5]$_SDFF_PN0__485  (.L_HI(net485));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[60]$_SDFF_PN0__486  (.L_HI(net486));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[61]$_SDFF_PN0__487  (.L_HI(net487));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[62]$_SDFF_PN0__488  (.L_HI(net488));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[63]$_SDFF_PN0__489  (.L_HI(net489));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[6]$_SDFF_PN0__490  (.L_HI(net490));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[7]$_SDFF_PN0__491  (.L_HI(net491));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[8]$_SDFF_PN0__492  (.L_HI(net492));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_cycle[9]$_SDFF_PN0__493  (.L_HI(net493));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[0]$_SDFFE_PN0P__494  (.L_HI(net494));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[10]$_SDFFE_PN0P__495  (.L_HI(net495));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[11]$_SDFFE_PN0P__496  (.L_HI(net496));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[12]$_SDFFE_PN0P__497  (.L_HI(net497));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[13]$_SDFFE_PN0P__498  (.L_HI(net498));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[14]$_SDFFE_PN0P__499  (.L_HI(net499));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[15]$_SDFFE_PN0P__500  (.L_HI(net500));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[16]$_SDFFE_PN0P__501  (.L_HI(net501));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[17]$_SDFFE_PN0P__502  (.L_HI(net502));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[18]$_SDFFE_PN0P__503  (.L_HI(net503));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[19]$_SDFFE_PN0P__504  (.L_HI(net504));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[1]$_SDFFE_PN0P__505  (.L_HI(net505));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[20]$_SDFFE_PN0P__506  (.L_HI(net506));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[21]$_SDFFE_PN0P__507  (.L_HI(net507));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[22]$_SDFFE_PN0P__508  (.L_HI(net508));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[23]$_SDFFE_PN0P__509  (.L_HI(net509));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[24]$_SDFFE_PN0P__510  (.L_HI(net510));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[25]$_SDFFE_PN0P__511  (.L_HI(net511));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[26]$_SDFFE_PN0P__512  (.L_HI(net512));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[27]$_SDFFE_PN0P__513  (.L_HI(net513));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[28]$_SDFFE_PN0P__514  (.L_HI(net514));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[29]$_SDFFE_PN0P__515  (.L_HI(net515));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[2]$_SDFFE_PN0P__516  (.L_HI(net516));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[30]$_SDFFE_PN0P__517  (.L_HI(net517));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[31]$_SDFFE_PN0P__518  (.L_HI(net518));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[32]$_SDFFE_PN0P__519  (.L_HI(net519));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[33]$_SDFFE_PN0P__520  (.L_HI(net520));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[34]$_SDFFE_PN0P__521  (.L_HI(net521));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[35]$_SDFFE_PN0P__522  (.L_HI(net522));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[36]$_SDFFE_PN0P__523  (.L_HI(net523));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[37]$_SDFFE_PN0P__524  (.L_HI(net524));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[38]$_SDFFE_PN0P__525  (.L_HI(net525));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[39]$_SDFFE_PN0P__526  (.L_HI(net526));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[3]$_SDFFE_PN0P__527  (.L_HI(net527));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[40]$_SDFFE_PN0P__528  (.L_HI(net528));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[41]$_SDFFE_PN0P__529  (.L_HI(net529));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[42]$_SDFFE_PN0P__530  (.L_HI(net530));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[43]$_SDFFE_PN0P__531  (.L_HI(net531));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[44]$_SDFFE_PN0P__532  (.L_HI(net532));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[45]$_SDFFE_PN0P__533  (.L_HI(net533));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[46]$_SDFFE_PN0P__534  (.L_HI(net534));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[47]$_SDFFE_PN0P__535  (.L_HI(net535));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[48]$_SDFFE_PN0P__536  (.L_HI(net536));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[49]$_SDFFE_PN0P__537  (.L_HI(net537));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[4]$_SDFFE_PN0P__538  (.L_HI(net538));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[50]$_SDFFE_PN0P__539  (.L_HI(net539));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[51]$_SDFFE_PN0P__540  (.L_HI(net540));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[52]$_SDFFE_PN0P__541  (.L_HI(net541));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[53]$_SDFFE_PN0P__542  (.L_HI(net542));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[54]$_SDFFE_PN0P__543  (.L_HI(net543));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[55]$_SDFFE_PN0P__544  (.L_HI(net544));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[56]$_SDFFE_PN0P__545  (.L_HI(net545));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[57]$_SDFFE_PN0P__546  (.L_HI(net546));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[58]$_SDFFE_PN0P__547  (.L_HI(net547));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[59]$_SDFFE_PN0P__548  (.L_HI(net548));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[5]$_SDFFE_PN0P__549  (.L_HI(net549));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[60]$_SDFFE_PN0P__550  (.L_HI(net550));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[61]$_SDFFE_PN0P__551  (.L_HI(net551));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[62]$_SDFFE_PN0P__552  (.L_HI(net552));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[63]$_SDFFE_PN0P__553  (.L_HI(net553));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[6]$_SDFFE_PN0P__554  (.L_HI(net554));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[7]$_SDFFE_PN0P__555  (.L_HI(net555));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[8]$_SDFFE_PN0P__556  (.L_HI(net556));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.count_instr[9]$_SDFFE_PN0P__557  (.L_HI(net557));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpu_state[0]$_DFF_P__558  (.L_HI(net558));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpu_state[1]$_DFF_P__559  (.L_HI(net559));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpu_state[2]$_DFF_P__560  (.L_HI(net560));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpu_state[3]$_DFF_P__561  (.L_HI(net561));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpu_state[4]$_DFF_P__562  (.L_HI(net562));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpu_state[5]$_DFF_P__563  (.L_HI(net563));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpu_state[6]$_DFF_P__564  (.L_HI(net564));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][0]$_DFFE_PP__565  (.L_HI(net565));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][10]$_DFFE_PP__566  (.L_HI(net566));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][11]$_DFFE_PP__567  (.L_HI(net567));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][12]$_DFFE_PP__568  (.L_HI(net568));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][13]$_DFFE_PP__569  (.L_HI(net569));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][14]$_DFFE_PP__570  (.L_HI(net570));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][15]$_DFFE_PP__571  (.L_HI(net571));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][16]$_DFFE_PP__572  (.L_HI(net572));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][17]$_DFFE_PP__573  (.L_HI(net573));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][18]$_DFFE_PP__574  (.L_HI(net574));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][19]$_DFFE_PP__575  (.L_HI(net575));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][1]$_DFFE_PP__576  (.L_HI(net576));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][20]$_DFFE_PP__577  (.L_HI(net577));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][21]$_DFFE_PP__578  (.L_HI(net578));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][22]$_DFFE_PP__579  (.L_HI(net579));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][23]$_DFFE_PP__580  (.L_HI(net580));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][24]$_DFFE_PP__581  (.L_HI(net581));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][25]$_DFFE_PP__582  (.L_HI(net582));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][26]$_DFFE_PP__583  (.L_HI(net583));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][27]$_DFFE_PP__584  (.L_HI(net584));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][28]$_DFFE_PP__585  (.L_HI(net585));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][29]$_DFFE_PP__586  (.L_HI(net586));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][2]$_DFFE_PP__587  (.L_HI(net587));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][30]$_DFFE_PP__588  (.L_HI(net588));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][31]$_DFFE_PP__589  (.L_HI(net589));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][3]$_DFFE_PP__590  (.L_HI(net590));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][4]$_DFFE_PP__591  (.L_HI(net591));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][5]$_DFFE_PP__592  (.L_HI(net592));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][6]$_DFFE_PP__593  (.L_HI(net593));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][7]$_DFFE_PP__594  (.L_HI(net594));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][8]$_DFFE_PP__595  (.L_HI(net595));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[0][9]$_DFFE_PP__596  (.L_HI(net596));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][0]$_DFFE_PP__597  (.L_HI(net597));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][10]$_DFFE_PP__598  (.L_HI(net598));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][11]$_DFFE_PP__599  (.L_HI(net599));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][12]$_DFFE_PP__600  (.L_HI(net600));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][13]$_DFFE_PP__601  (.L_HI(net601));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][14]$_DFFE_PP__602  (.L_HI(net602));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][15]$_DFFE_PP__603  (.L_HI(net603));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][16]$_DFFE_PP__604  (.L_HI(net604));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][17]$_DFFE_PP__605  (.L_HI(net605));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][18]$_DFFE_PP__606  (.L_HI(net606));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][19]$_DFFE_PP__607  (.L_HI(net607));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][1]$_DFFE_PP__608  (.L_HI(net608));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][20]$_DFFE_PP__609  (.L_HI(net609));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][21]$_DFFE_PP__610  (.L_HI(net610));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][22]$_DFFE_PP__611  (.L_HI(net611));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][23]$_DFFE_PP__612  (.L_HI(net612));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][24]$_DFFE_PP__613  (.L_HI(net613));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][25]$_DFFE_PP__614  (.L_HI(net614));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][26]$_DFFE_PP__615  (.L_HI(net615));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][27]$_DFFE_PP__616  (.L_HI(net616));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][28]$_DFFE_PP__617  (.L_HI(net617));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][29]$_DFFE_PP__618  (.L_HI(net618));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][2]$_DFFE_PP__619  (.L_HI(net619));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][30]$_DFFE_PP__620  (.L_HI(net620));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][31]$_DFFE_PP__621  (.L_HI(net621));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][3]$_DFFE_PP__622  (.L_HI(net622));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][4]$_DFFE_PP__623  (.L_HI(net623));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][5]$_DFFE_PP__624  (.L_HI(net624));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][6]$_DFFE_PP__625  (.L_HI(net625));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][7]$_DFFE_PP__626  (.L_HI(net626));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][8]$_DFFE_PP__627  (.L_HI(net627));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[10][9]$_DFFE_PP__628  (.L_HI(net628));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][0]$_DFFE_PP__629  (.L_HI(net629));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][10]$_DFFE_PP__630  (.L_HI(net630));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][11]$_DFFE_PP__631  (.L_HI(net631));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][12]$_DFFE_PP__632  (.L_HI(net632));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][13]$_DFFE_PP__633  (.L_HI(net633));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][14]$_DFFE_PP__634  (.L_HI(net634));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][15]$_DFFE_PP__635  (.L_HI(net635));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][16]$_DFFE_PP__636  (.L_HI(net636));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][17]$_DFFE_PP__637  (.L_HI(net637));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][18]$_DFFE_PP__638  (.L_HI(net638));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][19]$_DFFE_PP__639  (.L_HI(net639));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][1]$_DFFE_PP__640  (.L_HI(net640));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][20]$_DFFE_PP__641  (.L_HI(net641));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][21]$_DFFE_PP__642  (.L_HI(net642));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][22]$_DFFE_PP__643  (.L_HI(net643));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][23]$_DFFE_PP__644  (.L_HI(net644));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][24]$_DFFE_PP__645  (.L_HI(net645));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][25]$_DFFE_PP__646  (.L_HI(net646));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][26]$_DFFE_PP__647  (.L_HI(net647));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][27]$_DFFE_PP__648  (.L_HI(net648));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][28]$_DFFE_PP__649  (.L_HI(net649));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][29]$_DFFE_PP__650  (.L_HI(net650));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][2]$_DFFE_PP__651  (.L_HI(net651));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][30]$_DFFE_PP__652  (.L_HI(net652));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][31]$_DFFE_PP__653  (.L_HI(net653));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][3]$_DFFE_PP__654  (.L_HI(net654));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][4]$_DFFE_PP__655  (.L_HI(net655));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][5]$_DFFE_PP__656  (.L_HI(net656));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][6]$_DFFE_PP__657  (.L_HI(net657));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][7]$_DFFE_PP__658  (.L_HI(net658));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][8]$_DFFE_PP__659  (.L_HI(net659));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[11][9]$_DFFE_PP__660  (.L_HI(net660));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][0]$_DFFE_PP__661  (.L_HI(net661));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][10]$_DFFE_PP__662  (.L_HI(net662));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][11]$_DFFE_PP__663  (.L_HI(net663));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][12]$_DFFE_PP__664  (.L_HI(net664));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][13]$_DFFE_PP__665  (.L_HI(net665));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][14]$_DFFE_PP__666  (.L_HI(net666));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][15]$_DFFE_PP__667  (.L_HI(net667));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][16]$_DFFE_PP__668  (.L_HI(net668));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][17]$_DFFE_PP__669  (.L_HI(net669));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][18]$_DFFE_PP__670  (.L_HI(net670));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][19]$_DFFE_PP__671  (.L_HI(net671));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][1]$_DFFE_PP__672  (.L_HI(net672));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][20]$_DFFE_PP__673  (.L_HI(net673));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][21]$_DFFE_PP__674  (.L_HI(net674));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][22]$_DFFE_PP__675  (.L_HI(net675));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][23]$_DFFE_PP__676  (.L_HI(net676));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][24]$_DFFE_PP__677  (.L_HI(net677));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][25]$_DFFE_PP__678  (.L_HI(net678));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][26]$_DFFE_PP__679  (.L_HI(net679));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][27]$_DFFE_PP__680  (.L_HI(net680));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][28]$_DFFE_PP__681  (.L_HI(net681));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][29]$_DFFE_PP__682  (.L_HI(net682));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][2]$_DFFE_PP__683  (.L_HI(net683));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][30]$_DFFE_PP__684  (.L_HI(net684));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][31]$_DFFE_PP__685  (.L_HI(net685));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][3]$_DFFE_PP__686  (.L_HI(net686));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][4]$_DFFE_PP__687  (.L_HI(net687));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][5]$_DFFE_PP__688  (.L_HI(net688));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][6]$_DFFE_PP__689  (.L_HI(net689));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][7]$_DFFE_PP__690  (.L_HI(net690));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][8]$_DFFE_PP__691  (.L_HI(net691));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[12][9]$_DFFE_PP__692  (.L_HI(net692));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][0]$_DFFE_PP__693  (.L_HI(net693));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][10]$_DFFE_PP__694  (.L_HI(net694));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][11]$_DFFE_PP__695  (.L_HI(net695));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][12]$_DFFE_PP__696  (.L_HI(net696));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][13]$_DFFE_PP__697  (.L_HI(net697));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][14]$_DFFE_PP__698  (.L_HI(net698));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][15]$_DFFE_PP__699  (.L_HI(net699));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][16]$_DFFE_PP__700  (.L_HI(net700));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][17]$_DFFE_PP__701  (.L_HI(net701));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][18]$_DFFE_PP__702  (.L_HI(net702));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][19]$_DFFE_PP__703  (.L_HI(net703));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][1]$_DFFE_PP__704  (.L_HI(net704));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][20]$_DFFE_PP__705  (.L_HI(net705));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][21]$_DFFE_PP__706  (.L_HI(net706));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][22]$_DFFE_PP__707  (.L_HI(net707));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][23]$_DFFE_PP__708  (.L_HI(net708));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][24]$_DFFE_PP__709  (.L_HI(net709));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][25]$_DFFE_PP__710  (.L_HI(net710));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][26]$_DFFE_PP__711  (.L_HI(net711));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][27]$_DFFE_PP__712  (.L_HI(net712));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][28]$_DFFE_PP__713  (.L_HI(net713));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][29]$_DFFE_PP__714  (.L_HI(net714));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][2]$_DFFE_PP__715  (.L_HI(net715));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][30]$_DFFE_PP__716  (.L_HI(net716));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][31]$_DFFE_PP__717  (.L_HI(net717));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][3]$_DFFE_PP__718  (.L_HI(net718));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][4]$_DFFE_PP__719  (.L_HI(net719));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][5]$_DFFE_PP__720  (.L_HI(net720));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][6]$_DFFE_PP__721  (.L_HI(net721));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][7]$_DFFE_PP__722  (.L_HI(net722));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][8]$_DFFE_PP__723  (.L_HI(net723));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[13][9]$_DFFE_PP__724  (.L_HI(net724));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][0]$_DFFE_PP__725  (.L_HI(net725));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][10]$_DFFE_PP__726  (.L_HI(net726));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][11]$_DFFE_PP__727  (.L_HI(net727));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][12]$_DFFE_PP__728  (.L_HI(net728));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][13]$_DFFE_PP__729  (.L_HI(net729));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][14]$_DFFE_PP__730  (.L_HI(net730));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][15]$_DFFE_PP__731  (.L_HI(net731));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][16]$_DFFE_PP__732  (.L_HI(net732));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][17]$_DFFE_PP__733  (.L_HI(net733));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][18]$_DFFE_PP__734  (.L_HI(net734));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][19]$_DFFE_PP__735  (.L_HI(net735));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][1]$_DFFE_PP__736  (.L_HI(net736));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][20]$_DFFE_PP__737  (.L_HI(net737));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][21]$_DFFE_PP__738  (.L_HI(net738));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][22]$_DFFE_PP__739  (.L_HI(net739));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][23]$_DFFE_PP__740  (.L_HI(net740));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][24]$_DFFE_PP__741  (.L_HI(net741));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][25]$_DFFE_PP__742  (.L_HI(net742));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][26]$_DFFE_PP__743  (.L_HI(net743));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][27]$_DFFE_PP__744  (.L_HI(net744));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][28]$_DFFE_PP__745  (.L_HI(net745));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][29]$_DFFE_PP__746  (.L_HI(net746));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][2]$_DFFE_PP__747  (.L_HI(net747));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][30]$_DFFE_PP__748  (.L_HI(net748));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][31]$_DFFE_PP__749  (.L_HI(net749));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][3]$_DFFE_PP__750  (.L_HI(net750));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][4]$_DFFE_PP__751  (.L_HI(net751));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][5]$_DFFE_PP__752  (.L_HI(net752));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][6]$_DFFE_PP__753  (.L_HI(net753));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][7]$_DFFE_PP__754  (.L_HI(net754));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][8]$_DFFE_PP__755  (.L_HI(net755));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[14][9]$_DFFE_PP__756  (.L_HI(net756));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][0]$_DFFE_PP__757  (.L_HI(net757));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][10]$_DFFE_PP__758  (.L_HI(net758));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][11]$_DFFE_PP__759  (.L_HI(net759));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][12]$_DFFE_PP__760  (.L_HI(net760));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][13]$_DFFE_PP__761  (.L_HI(net761));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][14]$_DFFE_PP__762  (.L_HI(net762));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][15]$_DFFE_PP__763  (.L_HI(net763));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][16]$_DFFE_PP__764  (.L_HI(net764));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][17]$_DFFE_PP__765  (.L_HI(net765));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][18]$_DFFE_PP__766  (.L_HI(net766));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][19]$_DFFE_PP__767  (.L_HI(net767));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][1]$_DFFE_PP__768  (.L_HI(net768));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][20]$_DFFE_PP__769  (.L_HI(net769));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][21]$_DFFE_PP__770  (.L_HI(net770));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][22]$_DFFE_PP__771  (.L_HI(net771));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][23]$_DFFE_PP__772  (.L_HI(net772));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][24]$_DFFE_PP__773  (.L_HI(net773));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][25]$_DFFE_PP__774  (.L_HI(net774));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][26]$_DFFE_PP__775  (.L_HI(net775));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][27]$_DFFE_PP__776  (.L_HI(net776));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][28]$_DFFE_PP__777  (.L_HI(net777));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][29]$_DFFE_PP__778  (.L_HI(net778));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][2]$_DFFE_PP__779  (.L_HI(net779));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][30]$_DFFE_PP__780  (.L_HI(net780));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][31]$_DFFE_PP__781  (.L_HI(net781));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][3]$_DFFE_PP__782  (.L_HI(net782));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][4]$_DFFE_PP__783  (.L_HI(net783));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][5]$_DFFE_PP__784  (.L_HI(net784));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][6]$_DFFE_PP__785  (.L_HI(net785));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][7]$_DFFE_PP__786  (.L_HI(net786));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][8]$_DFFE_PP__787  (.L_HI(net787));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[15][9]$_DFFE_PP__788  (.L_HI(net788));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][0]$_DFFE_PP__789  (.L_HI(net789));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][10]$_DFFE_PP__790  (.L_HI(net790));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][11]$_DFFE_PP__791  (.L_HI(net791));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][12]$_DFFE_PP__792  (.L_HI(net792));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][13]$_DFFE_PP__793  (.L_HI(net793));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][14]$_DFFE_PP__794  (.L_HI(net794));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][15]$_DFFE_PP__795  (.L_HI(net795));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][16]$_DFFE_PP__796  (.L_HI(net796));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][17]$_DFFE_PP__797  (.L_HI(net797));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][18]$_DFFE_PP__798  (.L_HI(net798));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][19]$_DFFE_PP__799  (.L_HI(net799));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][1]$_DFFE_PP__800  (.L_HI(net800));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][20]$_DFFE_PP__801  (.L_HI(net801));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][21]$_DFFE_PP__802  (.L_HI(net802));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][22]$_DFFE_PP__803  (.L_HI(net803));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][23]$_DFFE_PP__804  (.L_HI(net804));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][24]$_DFFE_PP__805  (.L_HI(net805));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][25]$_DFFE_PP__806  (.L_HI(net806));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][26]$_DFFE_PP__807  (.L_HI(net807));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][27]$_DFFE_PP__808  (.L_HI(net808));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][28]$_DFFE_PP__809  (.L_HI(net809));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][29]$_DFFE_PP__810  (.L_HI(net810));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][2]$_DFFE_PP__811  (.L_HI(net811));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][30]$_DFFE_PP__812  (.L_HI(net812));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][31]$_DFFE_PP__813  (.L_HI(net813));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][3]$_DFFE_PP__814  (.L_HI(net814));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][4]$_DFFE_PP__815  (.L_HI(net815));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][5]$_DFFE_PP__816  (.L_HI(net816));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][6]$_DFFE_PP__817  (.L_HI(net817));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][7]$_DFFE_PP__818  (.L_HI(net818));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][8]$_DFFE_PP__819  (.L_HI(net819));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[16][9]$_DFFE_PP__820  (.L_HI(net820));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][0]$_DFFE_PP__821  (.L_HI(net821));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][10]$_DFFE_PP__822  (.L_HI(net822));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][11]$_DFFE_PP__823  (.L_HI(net823));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][12]$_DFFE_PP__824  (.L_HI(net824));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][13]$_DFFE_PP__825  (.L_HI(net825));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][14]$_DFFE_PP__826  (.L_HI(net826));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][15]$_DFFE_PP__827  (.L_HI(net827));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][16]$_DFFE_PP__828  (.L_HI(net828));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][17]$_DFFE_PP__829  (.L_HI(net829));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][18]$_DFFE_PP__830  (.L_HI(net830));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][19]$_DFFE_PP__831  (.L_HI(net831));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][1]$_DFFE_PP__832  (.L_HI(net832));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][20]$_DFFE_PP__833  (.L_HI(net833));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][21]$_DFFE_PP__834  (.L_HI(net834));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][22]$_DFFE_PP__835  (.L_HI(net835));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][23]$_DFFE_PP__836  (.L_HI(net836));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][24]$_DFFE_PP__837  (.L_HI(net837));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][25]$_DFFE_PP__838  (.L_HI(net838));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][26]$_DFFE_PP__839  (.L_HI(net839));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][27]$_DFFE_PP__840  (.L_HI(net840));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][28]$_DFFE_PP__841  (.L_HI(net841));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][29]$_DFFE_PP__842  (.L_HI(net842));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][2]$_DFFE_PP__843  (.L_HI(net843));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][30]$_DFFE_PP__844  (.L_HI(net844));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][31]$_DFFE_PP__845  (.L_HI(net845));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][3]$_DFFE_PP__846  (.L_HI(net846));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][4]$_DFFE_PP__847  (.L_HI(net847));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][5]$_DFFE_PP__848  (.L_HI(net848));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][6]$_DFFE_PP__849  (.L_HI(net849));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][7]$_DFFE_PP__850  (.L_HI(net850));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][8]$_DFFE_PP__851  (.L_HI(net851));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[17][9]$_DFFE_PP__852  (.L_HI(net852));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][0]$_DFFE_PP__853  (.L_HI(net853));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][10]$_DFFE_PP__854  (.L_HI(net854));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][11]$_DFFE_PP__855  (.L_HI(net855));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][12]$_DFFE_PP__856  (.L_HI(net856));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][13]$_DFFE_PP__857  (.L_HI(net857));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][14]$_DFFE_PP__858  (.L_HI(net858));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][15]$_DFFE_PP__859  (.L_HI(net859));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][16]$_DFFE_PP__860  (.L_HI(net860));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][17]$_DFFE_PP__861  (.L_HI(net861));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][18]$_DFFE_PP__862  (.L_HI(net862));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][19]$_DFFE_PP__863  (.L_HI(net863));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][1]$_DFFE_PP__864  (.L_HI(net864));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][20]$_DFFE_PP__865  (.L_HI(net865));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][21]$_DFFE_PP__866  (.L_HI(net866));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][22]$_DFFE_PP__867  (.L_HI(net867));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][23]$_DFFE_PP__868  (.L_HI(net868));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][24]$_DFFE_PP__869  (.L_HI(net869));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][25]$_DFFE_PP__870  (.L_HI(net870));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][26]$_DFFE_PP__871  (.L_HI(net871));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][27]$_DFFE_PP__872  (.L_HI(net872));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][28]$_DFFE_PP__873  (.L_HI(net873));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][29]$_DFFE_PP__874  (.L_HI(net874));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][2]$_DFFE_PP__875  (.L_HI(net875));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][30]$_DFFE_PP__876  (.L_HI(net876));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][31]$_DFFE_PP__877  (.L_HI(net877));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][3]$_DFFE_PP__878  (.L_HI(net878));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][4]$_DFFE_PP__879  (.L_HI(net879));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][5]$_DFFE_PP__880  (.L_HI(net880));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][6]$_DFFE_PP__881  (.L_HI(net881));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][7]$_DFFE_PP__882  (.L_HI(net882));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][8]$_DFFE_PP__883  (.L_HI(net883));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[18][9]$_DFFE_PP__884  (.L_HI(net884));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][0]$_DFFE_PP__885  (.L_HI(net885));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][10]$_DFFE_PP__886  (.L_HI(net886));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][11]$_DFFE_PP__887  (.L_HI(net887));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][12]$_DFFE_PP__888  (.L_HI(net888));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][13]$_DFFE_PP__889  (.L_HI(net889));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][14]$_DFFE_PP__890  (.L_HI(net890));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][15]$_DFFE_PP__891  (.L_HI(net891));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][16]$_DFFE_PP__892  (.L_HI(net892));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][17]$_DFFE_PP__893  (.L_HI(net893));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][18]$_DFFE_PP__894  (.L_HI(net894));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][19]$_DFFE_PP__895  (.L_HI(net895));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][1]$_DFFE_PP__896  (.L_HI(net896));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][20]$_DFFE_PP__897  (.L_HI(net897));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][21]$_DFFE_PP__898  (.L_HI(net898));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][22]$_DFFE_PP__899  (.L_HI(net899));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][23]$_DFFE_PP__900  (.L_HI(net900));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][24]$_DFFE_PP__901  (.L_HI(net901));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][25]$_DFFE_PP__902  (.L_HI(net902));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][26]$_DFFE_PP__903  (.L_HI(net903));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][27]$_DFFE_PP__904  (.L_HI(net904));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][28]$_DFFE_PP__905  (.L_HI(net905));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][29]$_DFFE_PP__906  (.L_HI(net906));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][2]$_DFFE_PP__907  (.L_HI(net907));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][30]$_DFFE_PP__908  (.L_HI(net908));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][31]$_DFFE_PP__909  (.L_HI(net909));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][3]$_DFFE_PP__910  (.L_HI(net910));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][4]$_DFFE_PP__911  (.L_HI(net911));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][5]$_DFFE_PP__912  (.L_HI(net912));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][6]$_DFFE_PP__913  (.L_HI(net913));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][7]$_DFFE_PP__914  (.L_HI(net914));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][8]$_DFFE_PP__915  (.L_HI(net915));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[19][9]$_DFFE_PP__916  (.L_HI(net916));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][0]$_DFFE_PP__917  (.L_HI(net917));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][10]$_DFFE_PP__918  (.L_HI(net918));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][11]$_DFFE_PP__919  (.L_HI(net919));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][12]$_DFFE_PP__920  (.L_HI(net920));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][13]$_DFFE_PP__921  (.L_HI(net921));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][14]$_DFFE_PP__922  (.L_HI(net922));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][15]$_DFFE_PP__923  (.L_HI(net923));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][16]$_DFFE_PP__924  (.L_HI(net924));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][17]$_DFFE_PP__925  (.L_HI(net925));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][18]$_DFFE_PP__926  (.L_HI(net926));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][19]$_DFFE_PP__927  (.L_HI(net927));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][1]$_DFFE_PP__928  (.L_HI(net928));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][20]$_DFFE_PP__929  (.L_HI(net929));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][21]$_DFFE_PP__930  (.L_HI(net930));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][22]$_DFFE_PP__931  (.L_HI(net931));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][23]$_DFFE_PP__932  (.L_HI(net932));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][24]$_DFFE_PP__933  (.L_HI(net933));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][25]$_DFFE_PP__934  (.L_HI(net934));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][26]$_DFFE_PP__935  (.L_HI(net935));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][27]$_DFFE_PP__936  (.L_HI(net936));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][28]$_DFFE_PP__937  (.L_HI(net937));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][29]$_DFFE_PP__938  (.L_HI(net938));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][2]$_DFFE_PP__939  (.L_HI(net939));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][30]$_DFFE_PP__940  (.L_HI(net940));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][31]$_DFFE_PP__941  (.L_HI(net941));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][3]$_DFFE_PP__942  (.L_HI(net942));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][4]$_DFFE_PP__943  (.L_HI(net943));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][5]$_DFFE_PP__944  (.L_HI(net944));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][6]$_DFFE_PP__945  (.L_HI(net945));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][7]$_DFFE_PP__946  (.L_HI(net946));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][8]$_DFFE_PP__947  (.L_HI(net947));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[1][9]$_DFFE_PP__948  (.L_HI(net948));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][0]$_DFFE_PP__949  (.L_HI(net949));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][10]$_DFFE_PP__950  (.L_HI(net950));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][11]$_DFFE_PP__951  (.L_HI(net951));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][12]$_DFFE_PP__952  (.L_HI(net952));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][13]$_DFFE_PP__953  (.L_HI(net953));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][14]$_DFFE_PP__954  (.L_HI(net954));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][15]$_DFFE_PP__955  (.L_HI(net955));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][16]$_DFFE_PP__956  (.L_HI(net956));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][17]$_DFFE_PP__957  (.L_HI(net957));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][18]$_DFFE_PP__958  (.L_HI(net958));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][19]$_DFFE_PP__959  (.L_HI(net959));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][1]$_DFFE_PP__960  (.L_HI(net960));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][20]$_DFFE_PP__961  (.L_HI(net961));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][21]$_DFFE_PP__962  (.L_HI(net962));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][22]$_DFFE_PP__963  (.L_HI(net963));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][23]$_DFFE_PP__964  (.L_HI(net964));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][24]$_DFFE_PP__965  (.L_HI(net965));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][25]$_DFFE_PP__966  (.L_HI(net966));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][26]$_DFFE_PP__967  (.L_HI(net967));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][27]$_DFFE_PP__968  (.L_HI(net968));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][28]$_DFFE_PP__969  (.L_HI(net969));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][29]$_DFFE_PP__970  (.L_HI(net970));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][2]$_DFFE_PP__971  (.L_HI(net971));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][30]$_DFFE_PP__972  (.L_HI(net972));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][31]$_DFFE_PP__973  (.L_HI(net973));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][3]$_DFFE_PP__974  (.L_HI(net974));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][4]$_DFFE_PP__975  (.L_HI(net975));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][5]$_DFFE_PP__976  (.L_HI(net976));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][6]$_DFFE_PP__977  (.L_HI(net977));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][7]$_DFFE_PP__978  (.L_HI(net978));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][8]$_DFFE_PP__979  (.L_HI(net979));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[20][9]$_DFFE_PP__980  (.L_HI(net980));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][0]$_DFFE_PP__981  (.L_HI(net981));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][10]$_DFFE_PP__982  (.L_HI(net982));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][11]$_DFFE_PP__983  (.L_HI(net983));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][12]$_DFFE_PP__984  (.L_HI(net984));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][13]$_DFFE_PP__985  (.L_HI(net985));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][14]$_DFFE_PP__986  (.L_HI(net986));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][15]$_DFFE_PP__987  (.L_HI(net987));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][16]$_DFFE_PP__988  (.L_HI(net988));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][17]$_DFFE_PP__989  (.L_HI(net989));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][18]$_DFFE_PP__990  (.L_HI(net990));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][19]$_DFFE_PP__991  (.L_HI(net991));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][1]$_DFFE_PP__992  (.L_HI(net992));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][20]$_DFFE_PP__993  (.L_HI(net993));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][21]$_DFFE_PP__994  (.L_HI(net994));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][22]$_DFFE_PP__995  (.L_HI(net995));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][23]$_DFFE_PP__996  (.L_HI(net996));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][24]$_DFFE_PP__997  (.L_HI(net997));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][25]$_DFFE_PP__998  (.L_HI(net998));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][26]$_DFFE_PP__999  (.L_HI(net999));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][27]$_DFFE_PP__1000  (.L_HI(net1000));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][28]$_DFFE_PP__1001  (.L_HI(net1001));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][29]$_DFFE_PP__1002  (.L_HI(net1002));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][2]$_DFFE_PP__1003  (.L_HI(net1003));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][30]$_DFFE_PP__1004  (.L_HI(net1004));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][31]$_DFFE_PP__1005  (.L_HI(net1005));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][3]$_DFFE_PP__1006  (.L_HI(net1006));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][4]$_DFFE_PP__1007  (.L_HI(net1007));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][5]$_DFFE_PP__1008  (.L_HI(net1008));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][6]$_DFFE_PP__1009  (.L_HI(net1009));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][7]$_DFFE_PP__1010  (.L_HI(net1010));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][8]$_DFFE_PP__1011  (.L_HI(net1011));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[21][9]$_DFFE_PP__1012  (.L_HI(net1012));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][0]$_DFFE_PP__1013  (.L_HI(net1013));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][10]$_DFFE_PP__1014  (.L_HI(net1014));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][11]$_DFFE_PP__1015  (.L_HI(net1015));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][12]$_DFFE_PP__1016  (.L_HI(net1016));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][13]$_DFFE_PP__1017  (.L_HI(net1017));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][14]$_DFFE_PP__1018  (.L_HI(net1018));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][15]$_DFFE_PP__1019  (.L_HI(net1019));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][16]$_DFFE_PP__1020  (.L_HI(net1020));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][17]$_DFFE_PP__1021  (.L_HI(net1021));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][18]$_DFFE_PP__1022  (.L_HI(net1022));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][19]$_DFFE_PP__1023  (.L_HI(net1023));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][1]$_DFFE_PP__1024  (.L_HI(net1024));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][20]$_DFFE_PP__1025  (.L_HI(net1025));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][21]$_DFFE_PP__1026  (.L_HI(net1026));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][22]$_DFFE_PP__1027  (.L_HI(net1027));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][23]$_DFFE_PP__1028  (.L_HI(net1028));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][24]$_DFFE_PP__1029  (.L_HI(net1029));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][25]$_DFFE_PP__1030  (.L_HI(net1030));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][26]$_DFFE_PP__1031  (.L_HI(net1031));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][27]$_DFFE_PP__1032  (.L_HI(net1032));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][28]$_DFFE_PP__1033  (.L_HI(net1033));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][29]$_DFFE_PP__1034  (.L_HI(net1034));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][2]$_DFFE_PP__1035  (.L_HI(net1035));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][30]$_DFFE_PP__1036  (.L_HI(net1036));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][31]$_DFFE_PP__1037  (.L_HI(net1037));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][3]$_DFFE_PP__1038  (.L_HI(net1038));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][4]$_DFFE_PP__1039  (.L_HI(net1039));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][5]$_DFFE_PP__1040  (.L_HI(net1040));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][6]$_DFFE_PP__1041  (.L_HI(net1041));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][7]$_DFFE_PP__1042  (.L_HI(net1042));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][8]$_DFFE_PP__1043  (.L_HI(net1043));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[22][9]$_DFFE_PP__1044  (.L_HI(net1044));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][0]$_DFFE_PP__1045  (.L_HI(net1045));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][10]$_DFFE_PP__1046  (.L_HI(net1046));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][11]$_DFFE_PP__1047  (.L_HI(net1047));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][12]$_DFFE_PP__1048  (.L_HI(net1048));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][13]$_DFFE_PP__1049  (.L_HI(net1049));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][14]$_DFFE_PP__1050  (.L_HI(net1050));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][15]$_DFFE_PP__1051  (.L_HI(net1051));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][16]$_DFFE_PP__1052  (.L_HI(net1052));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][17]$_DFFE_PP__1053  (.L_HI(net1053));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][18]$_DFFE_PP__1054  (.L_HI(net1054));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][19]$_DFFE_PP__1055  (.L_HI(net1055));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][1]$_DFFE_PP__1056  (.L_HI(net1056));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][20]$_DFFE_PP__1057  (.L_HI(net1057));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][21]$_DFFE_PP__1058  (.L_HI(net1058));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][22]$_DFFE_PP__1059  (.L_HI(net1059));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][23]$_DFFE_PP__1060  (.L_HI(net1060));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][24]$_DFFE_PP__1061  (.L_HI(net1061));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][25]$_DFFE_PP__1062  (.L_HI(net1062));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][26]$_DFFE_PP__1063  (.L_HI(net1063));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][27]$_DFFE_PP__1064  (.L_HI(net1064));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][28]$_DFFE_PP__1065  (.L_HI(net1065));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][29]$_DFFE_PP__1066  (.L_HI(net1066));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][2]$_DFFE_PP__1067  (.L_HI(net1067));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][30]$_DFFE_PP__1068  (.L_HI(net1068));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][31]$_DFFE_PP__1069  (.L_HI(net1069));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][3]$_DFFE_PP__1070  (.L_HI(net1070));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][4]$_DFFE_PP__1071  (.L_HI(net1071));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][5]$_DFFE_PP__1072  (.L_HI(net1072));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][6]$_DFFE_PP__1073  (.L_HI(net1073));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][7]$_DFFE_PP__1074  (.L_HI(net1074));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][8]$_DFFE_PP__1075  (.L_HI(net1075));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[23][9]$_DFFE_PP__1076  (.L_HI(net1076));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][0]$_DFFE_PP__1077  (.L_HI(net1077));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][10]$_DFFE_PP__1078  (.L_HI(net1078));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][11]$_DFFE_PP__1079  (.L_HI(net1079));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][12]$_DFFE_PP__1080  (.L_HI(net1080));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][13]$_DFFE_PP__1081  (.L_HI(net1081));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][14]$_DFFE_PP__1082  (.L_HI(net1082));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][15]$_DFFE_PP__1083  (.L_HI(net1083));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][16]$_DFFE_PP__1084  (.L_HI(net1084));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][17]$_DFFE_PP__1085  (.L_HI(net1085));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][18]$_DFFE_PP__1086  (.L_HI(net1086));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][19]$_DFFE_PP__1087  (.L_HI(net1087));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][1]$_DFFE_PP__1088  (.L_HI(net1088));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][20]$_DFFE_PP__1089  (.L_HI(net1089));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][21]$_DFFE_PP__1090  (.L_HI(net1090));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][22]$_DFFE_PP__1091  (.L_HI(net1091));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][23]$_DFFE_PP__1092  (.L_HI(net1092));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][24]$_DFFE_PP__1093  (.L_HI(net1093));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][25]$_DFFE_PP__1094  (.L_HI(net1094));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][26]$_DFFE_PP__1095  (.L_HI(net1095));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][27]$_DFFE_PP__1096  (.L_HI(net1096));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][28]$_DFFE_PP__1097  (.L_HI(net1097));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][29]$_DFFE_PP__1098  (.L_HI(net1098));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][2]$_DFFE_PP__1099  (.L_HI(net1099));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][30]$_DFFE_PP__1100  (.L_HI(net1100));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][31]$_DFFE_PP__1101  (.L_HI(net1101));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][3]$_DFFE_PP__1102  (.L_HI(net1102));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][4]$_DFFE_PP__1103  (.L_HI(net1103));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][5]$_DFFE_PP__1104  (.L_HI(net1104));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][6]$_DFFE_PP__1105  (.L_HI(net1105));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][7]$_DFFE_PP__1106  (.L_HI(net1106));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][8]$_DFFE_PP__1107  (.L_HI(net1107));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[24][9]$_DFFE_PP__1108  (.L_HI(net1108));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][0]$_DFFE_PP__1109  (.L_HI(net1109));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][10]$_DFFE_PP__1110  (.L_HI(net1110));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][11]$_DFFE_PP__1111  (.L_HI(net1111));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][12]$_DFFE_PP__1112  (.L_HI(net1112));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][13]$_DFFE_PP__1113  (.L_HI(net1113));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][14]$_DFFE_PP__1114  (.L_HI(net1114));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][15]$_DFFE_PP__1115  (.L_HI(net1115));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][16]$_DFFE_PP__1116  (.L_HI(net1116));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][17]$_DFFE_PP__1117  (.L_HI(net1117));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][18]$_DFFE_PP__1118  (.L_HI(net1118));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][19]$_DFFE_PP__1119  (.L_HI(net1119));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][1]$_DFFE_PP__1120  (.L_HI(net1120));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][20]$_DFFE_PP__1121  (.L_HI(net1121));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][21]$_DFFE_PP__1122  (.L_HI(net1122));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][22]$_DFFE_PP__1123  (.L_HI(net1123));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][23]$_DFFE_PP__1124  (.L_HI(net1124));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][24]$_DFFE_PP__1125  (.L_HI(net1125));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][25]$_DFFE_PP__1126  (.L_HI(net1126));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][26]$_DFFE_PP__1127  (.L_HI(net1127));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][27]$_DFFE_PP__1128  (.L_HI(net1128));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][28]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][29]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][2]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][30]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][31]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][3]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][4]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][5]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][6]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][7]$_DFFE_PP__1138  (.L_HI(net1138));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][8]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[25][9]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][0]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][10]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][11]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][12]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][13]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][14]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][15]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][16]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][17]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][18]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][19]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][1]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][20]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][21]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][22]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][23]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][24]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][25]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][26]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][27]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][28]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][29]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][2]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][30]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][31]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][3]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][4]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][5]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][6]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][7]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][8]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[26][9]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][0]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][10]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][11]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][12]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][13]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][14]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][15]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][16]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][17]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][18]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][19]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][1]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][20]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][21]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][22]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][23]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][24]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][25]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][26]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][27]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][28]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][29]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][2]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][30]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][31]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][3]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][4]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][5]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][6]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][7]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][8]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[27][9]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][0]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][10]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][11]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][12]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][13]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][14]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][15]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][16]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][17]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][18]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][19]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][1]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][20]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][21]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][22]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][23]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][24]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][25]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][26]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][27]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][28]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][29]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][2]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][30]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][31]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][3]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][4]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][5]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][6]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][7]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][8]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[28][9]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][0]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][10]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][11]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][12]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][13]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][14]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][15]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][16]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][17]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][18]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][19]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][1]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][20]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][21]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][22]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][23]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][24]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][25]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][26]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][27]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][28]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][29]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][2]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][30]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][31]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][3]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][4]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][5]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][6]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][7]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][8]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[29][9]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][0]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][10]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][11]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][12]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][13]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][14]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][15]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][16]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][17]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][18]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][19]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][1]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][20]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][21]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][22]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][23]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][24]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][25]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][26]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][27]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][28]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][29]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][2]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][30]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][31]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][3]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][4]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][5]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][6]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][7]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][8]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[2][9]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][0]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][10]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][11]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][12]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][13]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][14]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][15]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][16]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][17]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][18]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][19]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][1]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][20]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][21]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][22]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][23]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][24]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][25]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][26]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][27]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][28]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][29]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][2]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][30]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][31]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][3]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][4]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][5]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][6]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][7]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][8]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[30][9]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][0]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][10]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][11]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][12]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][13]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][14]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][15]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][16]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][17]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][18]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][19]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][1]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][20]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][21]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][22]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][23]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][24]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][25]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][26]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][27]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][28]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][29]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][2]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][30]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][31]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][3]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][4]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][5]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][6]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][7]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][8]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[31][9]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][0]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][10]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][11]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][12]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][13]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][14]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][15]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][16]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][17]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][18]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][19]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][1]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][20]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][21]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][22]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][23]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][24]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][25]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][26]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][27]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][28]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][29]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][2]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][30]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][31]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][3]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][4]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][5]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][6]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][7]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][8]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[3][9]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][0]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][10]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][11]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][12]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][13]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][14]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][15]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][16]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][17]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][18]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][19]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][1]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][20]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][21]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][22]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][23]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][24]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][25]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][26]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][27]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][28]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][29]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][2]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][30]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][31]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][3]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][4]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][5]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][6]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][7]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][8]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[4][9]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][0]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][10]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][11]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][12]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][13]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][14]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][15]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][16]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][17]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][18]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][19]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][1]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][20]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][21]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][22]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][23]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][24]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][25]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][26]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][27]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][28]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][29]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][2]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][30]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][31]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][3]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][4]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][5]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][6]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][7]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][8]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[5][9]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][0]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][10]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][11]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][12]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][13]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][14]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][15]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][16]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][17]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][18]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][19]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][1]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][20]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][21]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][22]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][23]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][24]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][25]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][26]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][27]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][28]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][29]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][2]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][30]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][31]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][3]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][4]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][5]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][6]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][7]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][8]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[6][9]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][0]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][10]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][11]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][12]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][13]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][14]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][15]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][16]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][17]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][18]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][19]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][1]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][20]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][21]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][22]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][23]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][24]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][25]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][26]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][27]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][28]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][29]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][2]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][30]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][31]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][3]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][4]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][5]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][6]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][7]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][8]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[7][9]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][0]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][10]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][11]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][12]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][13]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][14]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][15]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][16]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][17]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][18]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][19]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][1]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][20]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][21]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][22]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][23]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][24]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][25]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][26]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][27]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][28]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][29]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][2]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][30]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][31]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][3]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][4]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][5]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][6]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][7]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][8]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[8][9]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][0]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][10]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][11]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][12]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][13]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][14]$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][15]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][16]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][17]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][18]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][19]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][1]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][20]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][21]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][22]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][23]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][24]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][25]$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][26]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][27]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][28]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][29]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][2]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][30]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][31]$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][3]$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][4]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][5]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][6]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][7]$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][8]$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.cpuregs[9][9]$_DFFE_PP__1588  (.L_HI(net1588));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[0]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[10]$_SDFFCE_PN0P__1590  (.L_HI(net1590));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[11]$_SDFFCE_PN0P__1591  (.L_HI(net1591));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[12]$_SDFFCE_PN0P__1592  (.L_HI(net1592));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[13]$_SDFFCE_PN0P__1593  (.L_HI(net1593));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[14]$_SDFFCE_PN0P__1594  (.L_HI(net1594));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[15]$_SDFFCE_PN0P__1595  (.L_HI(net1595));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[16]$_SDFFCE_PN0P__1596  (.L_HI(net1596));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[17]$_SDFFCE_PN0P__1597  (.L_HI(net1597));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[18]$_SDFFCE_PN0P__1598  (.L_HI(net1598));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[19]$_SDFFCE_PN0P__1599  (.L_HI(net1599));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[1]$_SDFFCE_PN0P__1600  (.L_HI(net1600));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[20]$_SDFFCE_PN0P__1601  (.L_HI(net1601));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[21]$_SDFFCE_PN0P__1602  (.L_HI(net1602));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[22]$_SDFFCE_PN0P__1603  (.L_HI(net1603));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[23]$_SDFFCE_PN0P__1604  (.L_HI(net1604));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[24]$_SDFFCE_PN0P__1605  (.L_HI(net1605));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[25]$_SDFFCE_PN0P__1606  (.L_HI(net1606));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[26]$_SDFFCE_PN0P__1607  (.L_HI(net1607));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[27]$_SDFFCE_PN0P__1608  (.L_HI(net1608));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[28]$_SDFFCE_PN0P__1609  (.L_HI(net1609));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[29]$_SDFFCE_PN0P__1610  (.L_HI(net1610));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[2]$_SDFFCE_PN0P__1611  (.L_HI(net1611));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[30]$_SDFFCE_PN0P__1612  (.L_HI(net1612));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[31]$_SDFFCE_PN0P__1613  (.L_HI(net1613));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[3]$_SDFFCE_PN0P__1614  (.L_HI(net1614));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[4]$_SDFFCE_PN0P__1615  (.L_HI(net1615));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[5]$_SDFFCE_PN0P__1616  (.L_HI(net1616));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[6]$_SDFFCE_PN0P__1617  (.L_HI(net1617));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[7]$_SDFFCE_PN0P__1618  (.L_HI(net1618));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[8]$_SDFFCE_PN0P__1619  (.L_HI(net1619));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm[9]$_SDFFCE_PN0P__1620  (.L_HI(net1620));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[10]$_DFFE_PN__1621  (.L_HI(net1621));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[11]$_DFFE_PN__1622  (.L_HI(net1622));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[12]$_DFFE_PN__1623  (.L_HI(net1623));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[13]$_DFFE_PN__1624  (.L_HI(net1624));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[14]$_DFFE_PN__1625  (.L_HI(net1625));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[15]$_DFFE_PN__1626  (.L_HI(net1626));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[16]$_DFFE_PN__1627  (.L_HI(net1627));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[17]$_DFFE_PN__1628  (.L_HI(net1628));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[18]$_DFFE_PN__1629  (.L_HI(net1629));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[19]$_DFFE_PN__1630  (.L_HI(net1630));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[1]$_DFFE_PN__1631  (.L_HI(net1631));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[20]$_DFFE_PN__1632  (.L_HI(net1632));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[2]$_DFFE_PN__1633  (.L_HI(net1633));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[3]$_DFFE_PN__1634  (.L_HI(net1634));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[4]$_DFFE_PN__1635  (.L_HI(net1635));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[5]$_DFFE_PN__1636  (.L_HI(net1636));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[6]$_DFFE_PN__1637  (.L_HI(net1637));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[7]$_DFFE_PN__1638  (.L_HI(net1638));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[8]$_DFFE_PN__1639  (.L_HI(net1639));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_imm_j[9]$_DFFE_PN__1640  (.L_HI(net1640));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_rd[0]$_DFFE_PN__1641  (.L_HI(net1641));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_rd[1]$_DFFE_PN__1642  (.L_HI(net1642));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_rd[2]$_DFFE_PN__1643  (.L_HI(net1643));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_rd[3]$_DFFE_PN__1644  (.L_HI(net1644));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoded_rd[4]$_DFFE_PN__1645  (.L_HI(net1645));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoder_pseudo_trigger$_SDFF_PN0__1646  (.L_HI(net1646));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.decoder_trigger$_DFF_P__1647  (.L_HI(net1647));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_add$_SDFFE_PN0P__1648  (.L_HI(net1648));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_addi$_SDFFE_PN0P__1649  (.L_HI(net1649));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_and$_SDFFE_PN0P__1650  (.L_HI(net1650));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_andi$_SDFFE_PN0P__1651  (.L_HI(net1651));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_auipc$_DFFE_PN__1652  (.L_HI(net1652));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_beq$_SDFFE_PN0P__1653  (.L_HI(net1653));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_bge$_SDFFE_PN0P__1654  (.L_HI(net1654));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_bgeu$_SDFFE_PN0P__1655  (.L_HI(net1655));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_blt$_SDFFE_PN0P__1656  (.L_HI(net1656));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_bltu$_SDFFE_PN0P__1657  (.L_HI(net1657));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_bne$_SDFFE_PN0P__1658  (.L_HI(net1658));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_fence$_SDFFE_PN0P__1659  (.L_HI(net1659));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_jal$_DFFE_PN__1660  (.L_HI(net1660));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_jalr$_DFFE_PN__1661  (.L_HI(net1661));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_lb$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_lbu$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_lh$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_lhu$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_lui$_DFFE_PN__1666  (.L_HI(net1666));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_lw$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_or$_SDFFE_PN0P__1668  (.L_HI(net1668));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_ori$_SDFFE_PN0P__1669  (.L_HI(net1669));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_rdcycle$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_rdcycleh$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_rdinstr$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_rdinstrh$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_sb$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_sh$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_sll$_SDFFE_PN0P__1676  (.L_HI(net1676));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_slli$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_slt$_SDFFE_PN0P__1678  (.L_HI(net1678));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_slti$_SDFFE_PN0P__1679  (.L_HI(net1679));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_sltiu$_SDFFE_PN0P__1680  (.L_HI(net1680));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_sltu$_SDFFE_PN0P__1681  (.L_HI(net1681));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_sra$_SDFFE_PN0P__1682  (.L_HI(net1682));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_srai$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_srl$_SDFFE_PN0P__1684  (.L_HI(net1684));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_srli$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_sub$_SDFFE_PN0P__1686  (.L_HI(net1686));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_sw$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_xor$_SDFFE_PN0P__1688  (.L_HI(net1688));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.instr_xori$_SDFFE_PN0P__1689  (.L_HI(net1689));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_alu_reg_imm$_DFFE_PN__1690  (.L_HI(net1690));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_alu_reg_reg$_DFFE_PN__1691  (.L_HI(net1691));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_beq_bne_blt_bge_bltu_bgeu$_SDFFE_PN0N__1692  (.L_HI(net1692));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_compare$_SDFF_PP0__1693  (.L_HI(net1693));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_jalr_addi_slti_sltiu_xori_ori_andi$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_lb_lh_lw_lbu_lhu$_DFFE_PN__1695  (.L_HI(net1695));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_lui_auipc_jal$_DFF_P__1696  (.L_HI(net1696));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_sb_sh_sw$_DFFE_PN__1697  (.L_HI(net1697));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_sll_srl_sra$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_slli_srli_srai$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_slti_blt_slt$_DFF_P__1700  (.L_HI(net1700));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.is_sltiu_bltu_sltu$_DFF_P__1701  (.L_HI(net1701));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.latched_branch$_SDFFE_PN0P__1702  (.L_HI(net1702));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.latched_is_lb$_SDFFE_PN0P__1703  (.L_HI(net1703));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.latched_is_lh$_SDFFE_PN0P__1704  (.L_HI(net1704));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.latched_rd[0]$_SDFFCE_PP0P__1705  (.L_HI(net1705));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.latched_rd[1]$_SDFFCE_PP0P__1706  (.L_HI(net1706));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.latched_rd[2]$_SDFFCE_PP0P__1707  (.L_HI(net1707));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.latched_rd[3]$_SDFFCE_PP0P__1708  (.L_HI(net1708));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.latched_rd[4]$_SDFFCE_PP0P__1709  (.L_HI(net1709));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.latched_stalu$_SDFFE_PN0P__1710  (.L_HI(net1710));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.latched_store$_SDFFE_PN0P__1711  (.L_HI(net1711));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[10]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[11]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[12]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[13]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[14]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[15]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[16]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[17]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[18]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[19]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[20]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[21]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[22]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[23]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[24]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[25]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[26]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[27]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[28]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[29]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[2]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[30]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[31]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[3]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[4]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[5]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[6]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[7]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[8]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_addr[9]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_do_prefetch$_SDFFE_PP0P__1742  (.L_HI(net1742));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_do_rdata$_SDFFE_PP1P__1743  (.L_HI(net1743));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_do_rinst$_SDFFE_PP1P__1744  (.L_HI(net1744));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_do_wdata$_SDFFE_PP1P__1745  (.L_HI(net1745));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[0]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[10]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[11]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[12]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[13]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[14]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[15]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[16]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[17]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[18]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[19]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[1]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[20]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[21]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[22]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[23]$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[24]$_DFFE_PP__1762  (.L_HI(net1762));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[25]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[26]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[27]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[28]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[29]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[2]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[30]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[31]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[3]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[4]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[5]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[6]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[7]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[8]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_rdata_q[9]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_state[0]$_SDFFCE_PN0P__1778  (.L_HI(net1778));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_state[1]$_SDFFCE_PN0P__1779  (.L_HI(net1779));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_valid$_SDFFCE_PN0P__1780  (.L_HI(net1780));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[0]$_DFFE_PP__1781  (.L_HI(net1781));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[10]$_DFFE_PP__1782  (.L_HI(net1782));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[11]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[12]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[13]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[14]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[15]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[16]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[17]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[18]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[19]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[1]$_DFFE_PP__1792  (.L_HI(net1792));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[20]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[21]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[22]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[23]$_DFFE_PP__1796  (.L_HI(net1796));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[24]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[25]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[26]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[27]$_DFFE_PP__1800  (.L_HI(net1800));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[28]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[29]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[2]$_DFFE_PP__1803  (.L_HI(net1803));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[30]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[31]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[3]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[4]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[5]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[6]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[7]$_DFFE_PP__1810  (.L_HI(net1810));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[8]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wdata[9]$_DFFE_PP__1812  (.L_HI(net1812));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wordsize[0]$_DFF_P__1813  (.L_HI(net1813));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wordsize[1]$_DFF_P__1814  (.L_HI(net1814));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wordsize[2]$_DFF_P__1815  (.L_HI(net1815));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wstrb[0]$_DFFE_PP__1816  (.L_HI(net1816));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wstrb[1]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wstrb[2]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.mem_wstrb[3]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[10]$_SDFFE_PN0P__1820  (.L_HI(net1820));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[11]$_SDFFE_PN0P__1821  (.L_HI(net1821));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[12]$_SDFFE_PN0P__1822  (.L_HI(net1822));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[13]$_SDFFE_PN0P__1823  (.L_HI(net1823));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[14]$_SDFFE_PN0P__1824  (.L_HI(net1824));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[15]$_SDFFE_PN0P__1825  (.L_HI(net1825));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[16]$_SDFFE_PN0P__1826  (.L_HI(net1826));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[17]$_SDFFE_PN0P__1827  (.L_HI(net1827));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[18]$_SDFFE_PN0P__1828  (.L_HI(net1828));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[19]$_SDFFE_PN0P__1829  (.L_HI(net1829));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[1]$_SDFFE_PN0P__1830  (.L_HI(net1830));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[20]$_SDFFE_PN0P__1831  (.L_HI(net1831));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[21]$_SDFFE_PN0P__1832  (.L_HI(net1832));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[22]$_SDFFE_PN0P__1833  (.L_HI(net1833));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[23]$_SDFFE_PN0P__1834  (.L_HI(net1834));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[24]$_SDFFE_PN0P__1835  (.L_HI(net1835));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[25]$_SDFFE_PN0P__1836  (.L_HI(net1836));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[26]$_SDFFE_PN0P__1837  (.L_HI(net1837));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[27]$_SDFFE_PN0P__1838  (.L_HI(net1838));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[28]$_SDFFE_PN0P__1839  (.L_HI(net1839));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[29]$_SDFFE_PN0P__1840  (.L_HI(net1840));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[2]$_SDFFE_PN0P__1841  (.L_HI(net1841));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[30]$_SDFFE_PN0P__1842  (.L_HI(net1842));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[31]$_SDFFE_PN0P__1843  (.L_HI(net1843));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[3]$_SDFFE_PN0P__1844  (.L_HI(net1844));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[4]$_SDFFE_PN0P__1845  (.L_HI(net1845));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[5]$_SDFFE_PN0P__1846  (.L_HI(net1846));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[6]$_SDFFE_PN0P__1847  (.L_HI(net1847));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[7]$_SDFFE_PN0P__1848  (.L_HI(net1848));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[8]$_SDFFE_PN0P__1849  (.L_HI(net1849));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_next_pc[9]$_SDFFE_PN0P__1850  (.L_HI(net1850));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[0]$_DFFE_PP__1851  (.L_HI(net1851));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[10]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[11]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[12]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[13]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[14]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[15]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[16]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[17]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[18]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[19]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[1]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[20]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[21]$_DFFE_PP__1864  (.L_HI(net1864));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[22]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[23]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[24]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[25]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[26]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[27]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[28]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[29]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[2]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[30]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[31]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[3]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[4]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[5]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[6]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[7]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[8]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op1[9]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[0]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[10]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[11]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[12]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[13]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[14]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[15]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[16]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[17]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[18]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[19]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[1]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[20]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[21]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[22]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[23]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[24]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[25]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[26]$_DFFE_PP__1901  (.L_HI(net1901));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[27]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[28]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[29]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[2]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[30]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[31]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[3]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[4]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[5]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[6]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[7]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[8]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_op2[9]$_DFFE_PP__1914  (.L_HI(net1914));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[0]$_DFF_P__1915  (.L_HI(net1915));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[10]$_DFF_P__1916  (.L_HI(net1916));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[11]$_DFF_P__1917  (.L_HI(net1917));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[12]$_DFF_P__1918  (.L_HI(net1918));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[13]$_DFF_P__1919  (.L_HI(net1919));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[14]$_DFF_P__1920  (.L_HI(net1920));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[15]$_DFF_P__1921  (.L_HI(net1921));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[16]$_DFF_P__1922  (.L_HI(net1922));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[17]$_DFF_P__1923  (.L_HI(net1923));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[18]$_DFF_P__1924  (.L_HI(net1924));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[19]$_DFF_P__1925  (.L_HI(net1925));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[1]$_DFF_P__1926  (.L_HI(net1926));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[20]$_DFF_P__1927  (.L_HI(net1927));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[21]$_DFF_P__1928  (.L_HI(net1928));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[22]$_DFF_P__1929  (.L_HI(net1929));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[23]$_DFF_P__1930  (.L_HI(net1930));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[24]$_DFF_P__1931  (.L_HI(net1931));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[25]$_DFF_P__1932  (.L_HI(net1932));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[26]$_DFF_P__1933  (.L_HI(net1933));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[27]$_DFF_P__1934  (.L_HI(net1934));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[28]$_DFF_P__1935  (.L_HI(net1935));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[29]$_DFF_P__1936  (.L_HI(net1936));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[2]$_DFF_P__1937  (.L_HI(net1937));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[30]$_DFF_P__1938  (.L_HI(net1938));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[31]$_DFF_P__1939  (.L_HI(net1939));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[3]$_DFF_P__1940  (.L_HI(net1940));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[4]$_DFF_P__1941  (.L_HI(net1941));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[5]$_DFF_P__1942  (.L_HI(net1942));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[6]$_DFF_P__1943  (.L_HI(net1943));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[7]$_DFF_P__1944  (.L_HI(net1944));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[8]$_DFF_P__1945  (.L_HI(net1945));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_out[9]$_DFF_P__1946  (.L_HI(net1946));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[10]$_SDFFE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[11]$_SDFFE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[12]$_SDFFE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[13]$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[14]$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[15]$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[16]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[17]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[18]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[19]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[1]$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[20]$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[21]$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[22]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[23]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[24]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[25]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[26]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[27]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[28]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[29]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[2]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[30]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[31]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[3]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[4]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[5]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[6]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[7]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[8]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_pc[9]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_sh[0]$_DFFE_PP__1978  (.L_HI(net1978));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_sh[1]$_DFFE_PP__1979  (.L_HI(net1979));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_sh[2]$_DFF_P__1980  (.L_HI(net1980));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_sh[3]$_DFF_P__1981  (.L_HI(net1981));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.reg_sh[4]$_DFF_P__1982  (.L_HI(net1982));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_picorv32.trap$_SDFF_PN0__1983  (.L_HI(net1983));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[0]$_DFFE_PP__1984  (.L_HI(net1984));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[10]$_DFFE_PP__1985  (.L_HI(net1985));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[11]$_DFFE_PP__1986  (.L_HI(net1986));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[12]$_DFFE_PP__1987  (.L_HI(net1987));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[13]$_DFFE_PP__1988  (.L_HI(net1988));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[14]$_DFFE_PP__1989  (.L_HI(net1989));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[15]$_DFFE_PP__1990  (.L_HI(net1990));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[16]$_DFFE_PP__1991  (.L_HI(net1991));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[17]$_DFFE_PP__1992  (.L_HI(net1992));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[18]$_DFFE_PP__1993  (.L_HI(net1993));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[19]$_DFFE_PP__1994  (.L_HI(net1994));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[1]$_DFFE_PP__1995  (.L_HI(net1995));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[20]$_DFFE_PP__1996  (.L_HI(net1996));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[21]$_DFFE_PP__1997  (.L_HI(net1997));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[22]$_DFFE_PP__1998  (.L_HI(net1998));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[23]$_DFFE_PP__1999  (.L_HI(net1999));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[2]$_DFFE_PP__2000  (.L_HI(net2000));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[3]$_DFFE_PP__2001  (.L_HI(net2001));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[4]$_DFFE_PP__2002  (.L_HI(net2002));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[5]$_DFFE_PP__2003  (.L_HI(net2003));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[6]$_DFFE_PP__2004  (.L_HI(net2004));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[7]$_DFFE_PP__2005  (.L_HI(net2005));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[8]$_DFFE_PP__2006  (.L_HI(net2006));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.buffer[9]$_DFFE_PP__2007  (.L_HI(net2007));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_clk$_SDFFE_PN0P__2008  (.L_HI(net2008));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_cont$_SDFFE_PN0P__2009  (.L_HI(net2009));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_csb$_SDFFE_PN0P__2010  (.L_HI(net2010));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_ddr$_SDFFE_PN0P__2011  (.L_HI(net2011));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[0]$_SDFFE_PN0P__2012  (.L_HI(net2012));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[1]$_SDFFE_PN0P__2013  (.L_HI(net2013));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[2]$_SDFFE_PN0P__2014  (.L_HI(net2014));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_do[3]$_SDFFE_PN0P__2015  (.L_HI(net2015));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_dummy[0]$_SDFFE_PN0P__2016  (.L_HI(net2016));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_dummy[1]$_SDFFE_PN0P__2017  (.L_HI(net2017));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_dummy[2]$_SDFFE_PN0P__2018  (.L_HI(net2018));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_dummy[3]$_SDFFE_PN1P__2019  (.L_HI(net2019));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_en$_SDFFE_PN1P__2020  (.L_HI(net2020));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[0]$_SDFFE_PN0P__2021  (.L_HI(net2021));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[1]$_SDFFE_PN0P__2022  (.L_HI(net2022));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[2]$_SDFFE_PN0P__2023  (.L_HI(net2023));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_oe[3]$_SDFFE_PN0P__2024  (.L_HI(net2024));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.config_qspi$_SDFFE_PN0P__2025  (.L_HI(net2025));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[0]$_SDFFCE_PN1P__2026  (.L_HI(net2026));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[1]$_SDFFCE_PN1P__2027  (.L_HI(net2027));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[2]$_SDFFCE_PN1P__2028  (.L_HI(net2028));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[3]$_SDFFCE_PN1P__2029  (.L_HI(net2029));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[4]$_SDFFCE_PN1P__2030  (.L_HI(net2030));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[5]$_SDFFCE_PN1P__2031  (.L_HI(net2031));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[6]$_SDFFCE_PN1P__2032  (.L_HI(net2032));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_data[7]$_SDFFCE_PN1P__2033  (.L_HI(net2033));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_ddr$_SDFF_PP0__2034  (.L_HI(net2034));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_qspi$_SDFF_PP0__2035  (.L_HI(net2035));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_rd$_SDFFE_PP0P__2036  (.L_HI(net2036));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[0]$_SDFFE_PP0P__2037  (.L_HI(net2037));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[1]$_SDFFE_PP0P__2038  (.L_HI(net2038));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_tag[2]$_SDFFE_PP0P__2039  (.L_HI(net2039));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.din_valid$_SDFF_PP0__2040  (.L_HI(net2040));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[10]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[11]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[12]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[13]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[14]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[15]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[16]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[17]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[18]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[19]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[20]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[21]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[22]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[23]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[2]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[3]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[4]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[5]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[6]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[7]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[8]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_addr[9]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_inc$_SDFFCE_PP0P__2063  (.L_HI(net2063));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_valid$_SDFFE_PP0P__2064  (.L_HI(net2064));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rd_wait$_SDFFCE_PP0P__2065  (.L_HI(net2065));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[0]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[10]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[11]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[12]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[13]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[14]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[15]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[16]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[17]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[18]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[19]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[1]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[20]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[21]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[22]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[23]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[24]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[25]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[26]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[27]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[28]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[29]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[2]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[30]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[31]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[3]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[4]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[5]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[6]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[7]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[8]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.rdata[9]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.softreset$_SDFF_PN1__2098  (.L_HI(net2098));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[0]$_DFF_P__2099  (.L_HI(net2099));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[10]$_DFF_P__2100  (.L_HI(net2100));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[11]$_DFF_P__2101  (.L_HI(net2101));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[12]$_DFF_P__2102  (.L_HI(net2102));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[1]$_DFF_P__2103  (.L_HI(net2103));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[2]$_DFF_P__2104  (.L_HI(net2104));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[3]$_DFF_P__2105  (.L_HI(net2105));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[4]$_DFF_P__2106  (.L_HI(net2106));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[5]$_DFF_P__2107  (.L_HI(net2107));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[6]$_DFF_P__2108  (.L_HI(net2108));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[7]$_DFF_P__2109  (.L_HI(net2109));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[8]$_DFF_P__2110  (.L_HI(net2110));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.state[9]$_DFF_P__2111  (.L_HI(net2111));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[0]$_SDFFE_PP0P__2112  (.L_HI(net2112));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[1]$_SDFFE_PP0P__2113  (.L_HI(net2113));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[2]$_SDFFE_PP0P__2114  (.L_HI(net2114));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.count[3]$_SDFFE_PN0P__2115  (.L_HI(net2115));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[0]$_SDFFE_PN0N__2116  (.L_HI(net2116));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[1]$_SDFFE_PN0N__2117  (.L_HI(net2117));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[2]$_SDFFE_PN0N__2118  (.L_HI(net2118));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.dummy_count[3]$_SDFFE_PN0N__2119  (.L_HI(net2119));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.fetch$_SDFF_PN1__2120  (.L_HI(net2120));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_clk$_SDFFE_PP0P__2121  (.L_HI(net2121));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.flash_csb$_SDFFE_PN1P__2122  (.L_HI(net2122));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[0]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[1]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[2]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[3]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[4]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[5]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[6]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.ibuffer[7]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.last_fetch$_SDFF_PN1__2131  (.L_HI(net2131));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[0]$_SDFFCE_PN0P__2132  (.L_HI(net2132));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[1]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[2]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[3]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[4]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[5]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[6]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.obuffer[7]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr$_SDFFE_PN0P__2140  (.L_HI(net2140));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_ddr_q$_DFF_P__2141  (.L_HI(net2141));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_dspi$_SDFFE_PN0P__2142  (.L_HI(net2142));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_qspi$_SDFFE_PN0P__2143  (.L_HI(net2143));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_rd$_SDFFE_PN0P__2144  (.L_HI(net2144));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[0]$_SDFFE_PN0P__2145  (.L_HI(net2145));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[1]$_SDFFE_PN0P__2146  (.L_HI(net2146));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag[2]$_SDFFE_PN0P__2147  (.L_HI(net2147));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag_q[0]$_DFF_P__2148  (.L_HI(net2148));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag_q[1]$_DFF_P__2149  (.L_HI(net2149));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer.xfer_tag_q[2]$_DFF_P__2150  (.L_HI(net2150));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io0_90$_DFF_N__2151  (.L_HI(net2151));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io1_90$_DFF_N__2152  (.L_HI(net2152));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io2_90$_DFF_N__2153  (.L_HI(net2153));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_io3_90$_DFF_N__2154  (.L_HI(net2154));
 sg13g2_tiehi \u_ac_controller_soc_inst.u_spi_flash_mem.xfer_resetn$_SDFF_PP0__2155  (.L_HI(net2155));
 sg13g2_buf_16 clkbuf_leaf_834_clk (.X(clknet_leaf_834_clk),
    .A(clknet_8_171_0_clk));
 sg13g2_buf_16 clkbuf_leaf_835_clk (.X(clknet_leaf_835_clk),
    .A(clknet_8_172_0_clk));
 sg13g2_buf_16 clkbuf_leaf_836_clk (.X(clknet_leaf_836_clk),
    .A(clknet_8_175_0_clk));
 sg13g2_buf_16 clkbuf_leaf_837_clk (.X(clknet_leaf_837_clk),
    .A(clknet_8_173_0_clk));
 sg13g2_buf_16 clkbuf_leaf_838_clk (.X(clknet_leaf_838_clk),
    .A(clknet_8_173_0_clk));
 sg13g2_buf_16 clkbuf_leaf_840_clk (.X(clknet_leaf_840_clk),
    .A(clknet_8_172_0_clk));
 sg13g2_buf_16 clkbuf_leaf_841_clk (.X(clknet_leaf_841_clk),
    .A(clknet_8_172_0_clk));
 sg13g2_buf_16 clkbuf_leaf_842_clk (.X(clknet_leaf_842_clk),
    .A(clknet_8_166_0_clk));
 sg13g2_buf_16 clkbuf_leaf_845_clk (.X(clknet_leaf_845_clk),
    .A(clknet_8_163_0_clk));
 sg13g2_buf_16 clkbuf_leaf_847_clk (.X(clknet_leaf_847_clk),
    .A(clknet_8_169_0_clk));
 sg13g2_buf_16 clkbuf_leaf_848_clk (.X(clknet_leaf_848_clk),
    .A(clknet_8_163_0_clk));
 sg13g2_buf_16 clkbuf_leaf_849_clk (.X(clknet_leaf_849_clk),
    .A(clknet_8_162_0_clk));
 sg13g2_buf_16 clkbuf_leaf_850_clk (.X(clknet_leaf_850_clk),
    .A(clknet_8_162_0_clk));
 sg13g2_buf_16 clkbuf_leaf_851_clk (.X(clknet_leaf_851_clk),
    .A(clknet_8_162_0_clk));
 sg13g2_buf_16 clkbuf_leaf_852_clk (.X(clknet_leaf_852_clk),
    .A(clknet_8_143_0_clk));
 sg13g2_buf_16 clkbuf_leaf_853_clk (.X(clknet_leaf_853_clk),
    .A(clknet_8_161_0_clk));
 sg13g2_buf_16 clkbuf_leaf_854_clk (.X(clknet_leaf_854_clk),
    .A(clknet_8_161_0_clk));
 sg13g2_buf_16 clkbuf_leaf_857_clk (.X(clknet_leaf_857_clk),
    .A(clknet_8_161_0_clk));
 sg13g2_buf_16 clkbuf_leaf_858_clk (.X(clknet_leaf_858_clk),
    .A(clknet_8_169_0_clk));
 sg13g2_buf_16 clkbuf_leaf_859_clk (.X(clknet_leaf_859_clk),
    .A(clknet_8_169_0_clk));
 sg13g2_buf_16 clkbuf_leaf_860_clk (.X(clknet_leaf_860_clk),
    .A(clknet_8_168_0_clk));
 sg13g2_buf_16 clkbuf_leaf_861_clk (.X(clknet_leaf_861_clk),
    .A(clknet_8_168_0_clk));
 sg13g2_buf_16 clkbuf_leaf_863_clk (.X(clknet_leaf_863_clk),
    .A(clknet_8_168_0_clk));
 sg13g2_buf_16 clkbuf_leaf_865_clk (.X(clknet_leaf_865_clk),
    .A(clknet_8_160_0_clk));
 sg13g2_buf_16 clkbuf_leaf_867_clk (.X(clknet_leaf_867_clk),
    .A(clknet_8_160_0_clk));
 sg13g2_buf_16 clkbuf_leaf_868_clk (.X(clknet_leaf_868_clk),
    .A(clknet_8_160_0_clk));
 sg13g2_buf_16 clkbuf_leaf_869_clk (.X(clknet_leaf_869_clk),
    .A(clknet_8_138_0_clk));
 sg13g2_buf_16 clkbuf_leaf_870_clk (.X(clknet_leaf_870_clk),
    .A(clknet_8_138_0_clk));
 sg13g2_buf_16 clkbuf_leaf_873_clk (.X(clknet_leaf_873_clk),
    .A(clknet_8_139_0_clk));
 sg13g2_buf_16 clkbuf_leaf_874_clk (.X(clknet_leaf_874_clk),
    .A(clknet_8_160_0_clk));
 sg13g2_buf_16 clkbuf_leaf_875_clk (.X(clknet_leaf_875_clk),
    .A(clknet_8_142_0_clk));
 sg13g2_buf_16 clkbuf_leaf_877_clk (.X(clknet_leaf_877_clk),
    .A(clknet_8_142_0_clk));
 sg13g2_buf_16 clkbuf_leaf_878_clk (.X(clknet_leaf_878_clk),
    .A(clknet_8_142_0_clk));
 sg13g2_buf_16 clkbuf_leaf_879_clk (.X(clknet_leaf_879_clk),
    .A(clknet_8_139_0_clk));
 sg13g2_buf_16 clkbuf_leaf_882_clk (.X(clknet_leaf_882_clk),
    .A(clknet_8_137_0_clk));
 sg13g2_buf_16 clkbuf_leaf_883_clk (.X(clknet_leaf_883_clk),
    .A(clknet_8_139_0_clk));
 sg13g2_buf_16 clkbuf_leaf_884_clk (.X(clknet_leaf_884_clk),
    .A(clknet_8_138_0_clk));
 sg13g2_buf_16 clkbuf_leaf_886_clk (.X(clknet_leaf_886_clk),
    .A(clknet_8_136_0_clk));
 sg13g2_buf_16 clkbuf_leaf_887_clk (.X(clknet_leaf_887_clk),
    .A(clknet_8_136_0_clk));
 sg13g2_buf_16 clkbuf_leaf_888_clk (.X(clknet_leaf_888_clk),
    .A(clknet_8_136_0_clk));
 sg13g2_buf_16 clkbuf_leaf_890_clk (.X(clknet_leaf_890_clk),
    .A(clknet_8_130_0_clk));
 sg13g2_buf_16 clkbuf_leaf_891_clk (.X(clknet_leaf_891_clk),
    .A(clknet_8_130_0_clk));
 sg13g2_buf_16 clkbuf_leaf_892_clk (.X(clknet_leaf_892_clk),
    .A(clknet_8_130_0_clk));
 sg13g2_buf_16 clkbuf_leaf_893_clk (.X(clknet_leaf_893_clk),
    .A(clknet_8_131_0_clk));
 sg13g2_buf_16 clkbuf_leaf_894_clk (.X(clknet_leaf_894_clk),
    .A(clknet_8_131_0_clk));
 sg13g2_buf_16 clkbuf_leaf_896_clk (.X(clknet_leaf_896_clk),
    .A(clknet_8_134_0_clk));
 sg13g2_buf_16 clkbuf_leaf_898_clk (.X(clknet_leaf_898_clk),
    .A(clknet_8_131_0_clk));
 sg13g2_buf_16 clkbuf_leaf_899_clk (.X(clknet_leaf_899_clk),
    .A(clknet_8_134_0_clk));
 sg13g2_buf_16 clkbuf_leaf_900_clk (.X(clknet_leaf_900_clk),
    .A(clknet_8_140_0_clk));
 sg13g2_buf_16 clkbuf_leaf_902_clk (.X(clknet_leaf_902_clk),
    .A(clknet_8_140_0_clk));
 sg13g2_buf_16 clkbuf_leaf_903_clk (.X(clknet_leaf_903_clk),
    .A(clknet_8_140_0_clk));
 sg13g2_buf_16 clkbuf_leaf_904_clk (.X(clknet_leaf_904_clk),
    .A(clknet_8_142_0_clk));
 sg13g2_buf_16 clkbuf_leaf_905_clk (.X(clknet_leaf_905_clk),
    .A(clknet_8_142_0_clk));
 sg13g2_buf_16 clkbuf_leaf_907_clk (.X(clknet_leaf_907_clk),
    .A(clknet_8_141_0_clk));
 sg13g2_buf_16 clkbuf_leaf_909_clk (.X(clknet_leaf_909_clk),
    .A(clknet_8_141_0_clk));
 sg13g2_buf_16 clkbuf_leaf_910_clk (.X(clknet_leaf_910_clk),
    .A(clknet_8_135_0_clk));
 sg13g2_buf_16 clkbuf_leaf_912_clk (.X(clknet_leaf_912_clk),
    .A(clknet_8_135_0_clk));
 sg13g2_buf_16 clkbuf_leaf_914_clk (.X(clknet_leaf_914_clk),
    .A(clknet_8_152_0_clk));
 sg13g2_buf_16 clkbuf_leaf_916_clk (.X(clknet_leaf_916_clk),
    .A(clknet_8_152_0_clk));
 sg13g2_buf_16 clkbuf_leaf_917_clk (.X(clknet_leaf_917_clk),
    .A(clknet_8_153_0_clk));
 sg13g2_buf_16 clkbuf_leaf_920_clk (.X(clknet_leaf_920_clk),
    .A(clknet_8_154_0_clk));
 sg13g2_buf_16 clkbuf_leaf_921_clk (.X(clknet_leaf_921_clk),
    .A(clknet_8_155_0_clk));
 sg13g2_buf_16 clkbuf_leaf_923_clk (.X(clknet_leaf_923_clk),
    .A(clknet_8_154_0_clk));
 sg13g2_buf_16 clkbuf_leaf_924_clk (.X(clknet_leaf_924_clk),
    .A(clknet_8_164_0_clk));
 sg13g2_buf_16 clkbuf_leaf_926_clk (.X(clknet_leaf_926_clk),
    .A(clknet_8_154_0_clk));
 sg13g2_buf_16 clkbuf_leaf_927_clk (.X(clknet_leaf_927_clk),
    .A(clknet_8_143_0_clk));
 sg13g2_buf_16 clkbuf_leaf_929_clk (.X(clknet_leaf_929_clk),
    .A(clknet_8_143_0_clk));
 sg13g2_buf_16 clkbuf_leaf_930_clk (.X(clknet_leaf_930_clk),
    .A(clknet_8_162_0_clk));
 sg13g2_buf_16 clkbuf_leaf_931_clk (.X(clknet_leaf_931_clk),
    .A(clknet_8_164_0_clk));
 sg13g2_buf_16 clkbuf_leaf_932_clk (.X(clknet_leaf_932_clk),
    .A(clknet_8_162_0_clk));
 sg13g2_buf_16 clkbuf_leaf_933_clk (.X(clknet_leaf_933_clk),
    .A(clknet_8_166_0_clk));
 sg13g2_buf_16 clkbuf_leaf_934_clk (.X(clknet_leaf_934_clk),
    .A(clknet_8_164_0_clk));
 sg13g2_buf_16 clkbuf_leaf_935_clk (.X(clknet_leaf_935_clk),
    .A(clknet_8_164_0_clk));
 sg13g2_buf_16 clkbuf_leaf_936_clk (.X(clknet_leaf_936_clk),
    .A(clknet_8_164_0_clk));
 sg13g2_buf_16 clkbuf_leaf_937_clk (.X(clknet_leaf_937_clk),
    .A(clknet_8_165_0_clk));
 sg13g2_buf_16 clkbuf_leaf_938_clk (.X(clknet_leaf_938_clk),
    .A(clknet_8_166_0_clk));
 sg13g2_buf_16 clkbuf_leaf_941_clk (.X(clknet_leaf_941_clk),
    .A(clknet_8_167_0_clk));
 sg13g2_buf_16 clkbuf_leaf_942_clk (.X(clknet_leaf_942_clk),
    .A(clknet_8_167_0_clk));
 sg13g2_buf_16 clkbuf_leaf_943_clk (.X(clknet_leaf_943_clk),
    .A(clknet_8_250_0_clk));
 sg13g2_buf_16 clkbuf_leaf_946_clk (.X(clknet_leaf_946_clk),
    .A(clknet_8_165_0_clk));
 sg13g2_buf_16 clkbuf_leaf_948_clk (.X(clknet_leaf_948_clk),
    .A(clknet_8_155_0_clk));
 sg13g2_buf_16 clkbuf_leaf_949_clk (.X(clknet_leaf_949_clk),
    .A(clknet_8_158_0_clk));
 sg13g2_buf_16 clkbuf_leaf_951_clk (.X(clknet_leaf_951_clk),
    .A(clknet_8_248_0_clk));
 sg13g2_buf_16 clkbuf_leaf_952_clk (.X(clknet_leaf_952_clk),
    .A(clknet_8_248_0_clk));
 sg13g2_buf_16 clkbuf_leaf_953_clk (.X(clknet_leaf_953_clk),
    .A(clknet_8_248_0_clk));
 sg13g2_buf_16 clkbuf_leaf_954_clk (.X(clknet_leaf_954_clk),
    .A(clknet_8_248_0_clk));
 sg13g2_buf_16 clkbuf_leaf_955_clk (.X(clknet_leaf_955_clk),
    .A(clknet_8_159_0_clk));
 sg13g2_buf_16 clkbuf_leaf_956_clk (.X(clknet_leaf_956_clk),
    .A(clknet_8_158_0_clk));
 sg13g2_buf_16 clkbuf_leaf_957_clk (.X(clknet_leaf_957_clk),
    .A(clknet_8_159_0_clk));
 sg13g2_buf_16 clkbuf_leaf_960_clk (.X(clknet_leaf_960_clk),
    .A(clknet_8_155_0_clk));
 sg13g2_buf_16 clkbuf_leaf_961_clk (.X(clknet_leaf_961_clk),
    .A(clknet_8_155_0_clk));
 sg13g2_buf_16 clkbuf_leaf_962_clk (.X(clknet_leaf_962_clk),
    .A(clknet_8_156_0_clk));
 sg13g2_buf_16 clkbuf_leaf_963_clk (.X(clknet_leaf_963_clk),
    .A(clknet_8_156_0_clk));
 sg13g2_buf_16 clkbuf_leaf_965_clk (.X(clknet_leaf_965_clk),
    .A(clknet_8_156_0_clk));
 sg13g2_buf_16 clkbuf_leaf_966_clk (.X(clknet_leaf_966_clk),
    .A(clknet_8_156_0_clk));
 sg13g2_buf_16 clkbuf_leaf_968_clk (.X(clknet_leaf_968_clk),
    .A(clknet_8_157_0_clk));
 sg13g2_buf_16 clkbuf_leaf_969_clk (.X(clknet_leaf_969_clk),
    .A(clknet_8_157_0_clk));
 sg13g2_buf_16 clkbuf_leaf_972_clk (.X(clknet_leaf_972_clk),
    .A(clknet_8_242_0_clk));
 sg13g2_buf_16 clkbuf_leaf_974_clk (.X(clknet_leaf_974_clk),
    .A(clknet_8_242_0_clk));
 sg13g2_buf_16 clkbuf_leaf_978_clk (.X(clknet_leaf_978_clk),
    .A(clknet_8_242_0_clk));
 sg13g2_buf_16 clkbuf_leaf_982_clk (.X(clknet_leaf_982_clk),
    .A(clknet_8_241_0_clk));
 sg13g2_buf_16 clkbuf_leaf_988_clk (.X(clknet_leaf_988_clk),
    .A(clknet_8_149_0_clk));
 sg13g2_buf_16 clkbuf_leaf_990_clk (.X(clknet_leaf_990_clk),
    .A(clknet_8_148_0_clk));
 sg13g2_buf_16 clkbuf_leaf_991_clk (.X(clknet_leaf_991_clk),
    .A(clknet_8_150_0_clk));
 sg13g2_buf_16 clkbuf_leaf_994_clk (.X(clknet_leaf_994_clk),
    .A(clknet_8_151_0_clk));
 sg13g2_buf_16 clkbuf_leaf_995_clk (.X(clknet_leaf_995_clk),
    .A(clknet_8_150_0_clk));
 sg13g2_buf_16 clkbuf_leaf_997_clk (.X(clknet_leaf_997_clk),
    .A(clknet_8_150_0_clk));
 sg13g2_buf_16 clkbuf_leaf_998_clk (.X(clknet_leaf_998_clk),
    .A(clknet_8_147_0_clk));
 sg13g2_buf_16 clkbuf_leaf_999_clk (.X(clknet_leaf_999_clk),
    .A(clknet_8_150_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1000_clk (.X(clknet_leaf_1000_clk),
    .A(clknet_8_153_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1003_clk (.X(clknet_leaf_1003_clk),
    .A(clknet_8_145_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1004_clk (.X(clknet_leaf_1004_clk),
    .A(clknet_8_145_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1005_clk (.X(clknet_leaf_1005_clk),
    .A(clknet_8_60_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1006_clk (.X(clknet_leaf_1006_clk),
    .A(clknet_8_60_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1007_clk (.X(clknet_leaf_1007_clk),
    .A(clknet_8_63_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1009_clk (.X(clknet_leaf_1009_clk),
    .A(clknet_8_148_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1010_clk (.X(clknet_leaf_1010_clk),
    .A(clknet_8_148_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1011_clk (.X(clknet_leaf_1011_clk),
    .A(clknet_8_148_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1012_clk (.X(clknet_leaf_1012_clk),
    .A(clknet_8_14_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1015_clk (.X(clknet_leaf_1015_clk),
    .A(clknet_8_62_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1017_clk (.X(clknet_leaf_1017_clk),
    .A(clknet_8_62_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1018_clk (.X(clknet_leaf_1018_clk),
    .A(clknet_8_60_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1019_clk (.X(clknet_leaf_1019_clk),
    .A(clknet_8_60_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1020_clk (.X(clknet_leaf_1020_clk),
    .A(clknet_8_60_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1021_clk (.X(clknet_leaf_1021_clk),
    .A(clknet_8_61_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1022_clk (.X(clknet_leaf_1022_clk),
    .A(clknet_8_58_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1023_clk (.X(clknet_leaf_1023_clk),
    .A(clknet_8_58_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1026_clk (.X(clknet_leaf_1026_clk),
    .A(clknet_8_45_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1027_clk (.X(clknet_leaf_1027_clk),
    .A(clknet_8_45_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1028_clk (.X(clknet_leaf_1028_clk),
    .A(clknet_8_47_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1031_clk (.X(clknet_leaf_1031_clk),
    .A(clknet_8_45_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1032_clk (.X(clknet_leaf_1032_clk),
    .A(clknet_8_44_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1033_clk (.X(clknet_leaf_1033_clk),
    .A(clknet_8_44_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1034_clk (.X(clknet_leaf_1034_clk),
    .A(clknet_8_46_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1035_clk (.X(clknet_leaf_1035_clk),
    .A(clknet_8_43_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1037_clk (.X(clknet_leaf_1037_clk),
    .A(clknet_8_46_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1038_clk (.X(clknet_leaf_1038_clk),
    .A(clknet_8_144_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1040_clk (.X(clknet_leaf_1040_clk),
    .A(clknet_8_46_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1041_clk (.X(clknet_leaf_1041_clk),
    .A(clknet_8_47_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1043_clk (.X(clknet_leaf_1043_clk),
    .A(clknet_8_145_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1044_clk (.X(clknet_leaf_1044_clk),
    .A(clknet_8_144_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1045_clk (.X(clknet_leaf_1045_clk),
    .A(clknet_8_144_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1046_clk (.X(clknet_leaf_1046_clk),
    .A(clknet_8_147_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1047_clk (.X(clknet_leaf_1047_clk),
    .A(clknet_8_147_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1048_clk (.X(clknet_leaf_1048_clk),
    .A(clknet_8_146_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1049_clk (.X(clknet_leaf_1049_clk),
    .A(clknet_8_146_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1051_clk (.X(clknet_leaf_1051_clk),
    .A(clknet_8_146_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1052_clk (.X(clknet_leaf_1052_clk),
    .A(clknet_8_146_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1053_clk (.X(clknet_leaf_1053_clk),
    .A(clknet_8_135_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1054_clk (.X(clknet_leaf_1054_clk),
    .A(clknet_8_133_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1055_clk (.X(clknet_leaf_1055_clk),
    .A(clknet_8_133_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1056_clk (.X(clknet_leaf_1056_clk),
    .A(clknet_8_144_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1057_clk (.X(clknet_leaf_1057_clk),
    .A(clknet_8_132_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1058_clk (.X(clknet_leaf_1058_clk),
    .A(clknet_8_133_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1060_clk (.X(clknet_leaf_1060_clk),
    .A(clknet_8_133_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1061_clk (.X(clknet_leaf_1061_clk),
    .A(clknet_8_132_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1062_clk (.X(clknet_leaf_1062_clk),
    .A(clknet_8_129_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1063_clk (.X(clknet_leaf_1063_clk),
    .A(clknet_8_132_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1065_clk (.X(clknet_leaf_1065_clk),
    .A(clknet_8_132_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1066_clk (.X(clknet_leaf_1066_clk),
    .A(clknet_8_134_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1067_clk (.X(clknet_leaf_1067_clk),
    .A(clknet_8_134_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1069_clk (.X(clknet_leaf_1069_clk),
    .A(clknet_8_131_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1070_clk (.X(clknet_leaf_1070_clk),
    .A(clknet_8_130_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1071_clk (.X(clknet_leaf_1071_clk),
    .A(clknet_8_130_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1072_clk (.X(clknet_leaf_1072_clk),
    .A(clknet_8_128_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1073_clk (.X(clknet_leaf_1073_clk),
    .A(clknet_8_128_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1074_clk (.X(clknet_leaf_1074_clk),
    .A(clknet_8_128_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1075_clk (.X(clknet_leaf_1075_clk),
    .A(clknet_8_129_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1076_clk (.X(clknet_leaf_1076_clk),
    .A(clknet_8_128_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1077_clk (.X(clknet_leaf_1077_clk),
    .A(clknet_8_128_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1078_clk (.X(clknet_leaf_1078_clk),
    .A(clknet_8_42_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1079_clk (.X(clknet_leaf_1079_clk),
    .A(clknet_8_42_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1080_clk (.X(clknet_leaf_1080_clk),
    .A(clknet_8_42_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1081_clk (.X(clknet_leaf_1081_clk),
    .A(clknet_8_129_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1083_clk (.X(clknet_leaf_1083_clk),
    .A(clknet_8_42_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1084_clk (.X(clknet_leaf_1084_clk),
    .A(clknet_8_43_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1085_clk (.X(clknet_leaf_1085_clk),
    .A(clknet_8_42_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1086_clk (.X(clknet_leaf_1086_clk),
    .A(clknet_8_41_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1087_clk (.X(clknet_leaf_1087_clk),
    .A(clknet_8_35_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1088_clk (.X(clknet_leaf_1088_clk),
    .A(clknet_8_41_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1089_clk (.X(clknet_leaf_1089_clk),
    .A(clknet_8_40_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1090_clk (.X(clknet_leaf_1090_clk),
    .A(clknet_8_40_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1091_clk (.X(clknet_leaf_1091_clk),
    .A(clknet_8_40_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1092_clk (.X(clknet_leaf_1092_clk),
    .A(clknet_8_40_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1093_clk (.X(clknet_leaf_1093_clk),
    .A(clknet_8_34_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1096_clk (.X(clknet_leaf_1096_clk),
    .A(clknet_8_34_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1097_clk (.X(clknet_leaf_1097_clk),
    .A(clknet_8_34_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1098_clk (.X(clknet_leaf_1098_clk),
    .A(clknet_8_32_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1099_clk (.X(clknet_leaf_1099_clk),
    .A(clknet_8_32_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1101_clk (.X(clknet_leaf_1101_clk),
    .A(clknet_8_35_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1104_clk (.X(clknet_leaf_1104_clk),
    .A(clknet_8_36_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1105_clk (.X(clknet_leaf_1105_clk),
    .A(clknet_8_36_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1106_clk (.X(clknet_leaf_1106_clk),
    .A(clknet_8_38_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1109_clk (.X(clknet_leaf_1109_clk),
    .A(clknet_8_38_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1110_clk (.X(clknet_leaf_1110_clk),
    .A(clknet_8_41_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1112_clk (.X(clknet_leaf_1112_clk),
    .A(clknet_8_41_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1113_clk (.X(clknet_leaf_1113_clk),
    .A(clknet_8_44_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1114_clk (.X(clknet_leaf_1114_clk),
    .A(clknet_8_44_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1116_clk (.X(clknet_leaf_1116_clk),
    .A(clknet_8_38_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1120_clk (.X(clknet_leaf_1120_clk),
    .A(clknet_8_37_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1122_clk (.X(clknet_leaf_1122_clk),
    .A(clknet_8_39_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1124_clk (.X(clknet_leaf_1124_clk),
    .A(clknet_8_39_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1125_clk (.X(clknet_leaf_1125_clk),
    .A(clknet_8_56_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1126_clk (.X(clknet_leaf_1126_clk),
    .A(clknet_8_56_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1127_clk (.X(clknet_leaf_1127_clk),
    .A(clknet_8_57_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1128_clk (.X(clknet_leaf_1128_clk),
    .A(clknet_8_57_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1129_clk (.X(clknet_leaf_1129_clk),
    .A(clknet_8_57_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1131_clk (.X(clknet_leaf_1131_clk),
    .A(clknet_8_56_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1133_clk (.X(clknet_leaf_1133_clk),
    .A(clknet_8_56_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1134_clk (.X(clknet_leaf_1134_clk),
    .A(clknet_8_50_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1135_clk (.X(clknet_leaf_1135_clk),
    .A(clknet_8_50_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1136_clk (.X(clknet_leaf_1136_clk),
    .A(clknet_8_48_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1138_clk (.X(clknet_leaf_1138_clk),
    .A(clknet_8_50_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1139_clk (.X(clknet_leaf_1139_clk),
    .A(clknet_8_50_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1140_clk (.X(clknet_leaf_1140_clk),
    .A(clknet_8_33_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1142_clk (.X(clknet_leaf_1142_clk),
    .A(clknet_8_36_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1144_clk (.X(clknet_leaf_1144_clk),
    .A(clknet_8_33_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1145_clk (.X(clknet_leaf_1145_clk),
    .A(clknet_8_33_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1146_clk (.X(clknet_leaf_1146_clk),
    .A(clknet_8_32_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1147_clk (.X(clknet_leaf_1147_clk),
    .A(clknet_8_32_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1148_clk (.X(clknet_leaf_1148_clk),
    .A(clknet_8_32_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1149_clk (.X(clknet_leaf_1149_clk),
    .A(clknet_8_52_0_clk));
 sg13g2_buf_16 clkbuf_leaf_1150_clk (.X(clknet_leaf_1150_clk),
    .A(clknet_8_52_0_clk));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_16 clkbuf_1_0_0_clk (.X(clknet_1_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_1_0_1_clk (.X(clknet_1_0_1_clk),
    .A(clknet_1_0_0_clk));
 sg13g2_buf_16 clkbuf_1_1_0_clk (.X(clknet_1_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_1_1_1_clk (.X(clknet_1_1_1_clk),
    .A(clknet_1_1_0_clk));
 sg13g2_buf_16 clkbuf_2_0_0_clk (.X(clknet_2_0_0_clk),
    .A(clknet_1_0_1_clk));
 sg13g2_buf_16 clkbuf_2_0_1_clk (.X(clknet_2_0_1_clk),
    .A(clknet_2_0_0_clk));
 sg13g2_buf_16 clkbuf_2_1_0_clk (.X(clknet_2_1_0_clk),
    .A(clknet_1_0_1_clk));
 sg13g2_buf_16 clkbuf_2_1_1_clk (.X(clknet_2_1_1_clk),
    .A(clknet_2_1_0_clk));
 sg13g2_buf_16 clkbuf_2_2_0_clk (.X(clknet_2_2_0_clk),
    .A(clknet_1_1_1_clk));
 sg13g2_buf_16 clkbuf_2_2_1_clk (.X(clknet_2_2_1_clk),
    .A(clknet_2_2_0_clk));
 sg13g2_buf_16 clkbuf_2_3_0_clk (.X(clknet_2_3_0_clk),
    .A(clknet_1_1_1_clk));
 sg13g2_buf_16 clkbuf_2_3_1_clk (.X(clknet_2_3_1_clk),
    .A(clknet_2_3_0_clk));
 sg13g2_buf_16 clkbuf_3_0_0_clk (.X(clknet_3_0_0_clk),
    .A(clknet_2_0_1_clk));
 sg13g2_buf_16 clkbuf_3_1_0_clk (.X(clknet_3_1_0_clk),
    .A(clknet_2_0_1_clk));
 sg13g2_buf_16 clkbuf_3_2_0_clk (.X(clknet_3_2_0_clk),
    .A(clknet_2_1_1_clk));
 sg13g2_buf_16 clkbuf_3_3_0_clk (.X(clknet_3_3_0_clk),
    .A(clknet_2_1_1_clk));
 sg13g2_buf_16 clkbuf_3_4_0_clk (.X(clknet_3_4_0_clk),
    .A(clknet_2_2_1_clk));
 sg13g2_buf_16 clkbuf_3_5_0_clk (.X(clknet_3_5_0_clk),
    .A(clknet_2_2_1_clk));
 sg13g2_buf_16 clkbuf_3_6_0_clk (.X(clknet_3_6_0_clk),
    .A(clknet_2_3_1_clk));
 sg13g2_buf_16 clkbuf_3_7_0_clk (.X(clknet_3_7_0_clk),
    .A(clknet_2_3_1_clk));
 sg13g2_buf_16 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_16 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_16 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_16 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_16 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_16 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_16 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_16 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_16 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_16 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_16 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_16 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_16 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_16 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_16 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_16 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_16 clkbuf_5_0_0_clk (.X(clknet_5_0_0_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_16 clkbuf_5_1_0_clk (.X(clknet_5_1_0_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_16 clkbuf_5_2_0_clk (.X(clknet_5_2_0_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_16 clkbuf_5_3_0_clk (.X(clknet_5_3_0_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_16 clkbuf_5_4_0_clk (.X(clknet_5_4_0_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_16 clkbuf_5_5_0_clk (.X(clknet_5_5_0_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_16 clkbuf_5_6_0_clk (.X(clknet_5_6_0_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_16 clkbuf_5_7_0_clk (.X(clknet_5_7_0_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_16 clkbuf_5_8_0_clk (.X(clknet_5_8_0_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_16 clkbuf_5_9_0_clk (.X(clknet_5_9_0_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_16 clkbuf_5_10_0_clk (.X(clknet_5_10_0_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_16 clkbuf_5_11_0_clk (.X(clknet_5_11_0_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_16 clkbuf_5_12_0_clk (.X(clknet_5_12_0_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_16 clkbuf_5_13_0_clk (.X(clknet_5_13_0_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_16 clkbuf_5_14_0_clk (.X(clknet_5_14_0_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_16 clkbuf_5_15_0_clk (.X(clknet_5_15_0_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_16 clkbuf_5_16_0_clk (.X(clknet_5_16_0_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_16 clkbuf_5_17_0_clk (.X(clknet_5_17_0_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_16 clkbuf_5_18_0_clk (.X(clknet_5_18_0_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_16 clkbuf_5_19_0_clk (.X(clknet_5_19_0_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_16 clkbuf_5_20_0_clk (.X(clknet_5_20_0_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_16 clkbuf_5_21_0_clk (.X(clknet_5_21_0_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_16 clkbuf_5_22_0_clk (.X(clknet_5_22_0_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_16 clkbuf_5_23_0_clk (.X(clknet_5_23_0_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_16 clkbuf_5_24_0_clk (.X(clknet_5_24_0_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_16 clkbuf_5_25_0_clk (.X(clknet_5_25_0_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_16 clkbuf_5_26_0_clk (.X(clknet_5_26_0_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_16 clkbuf_5_27_0_clk (.X(clknet_5_27_0_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_16 clkbuf_5_28_0_clk (.X(clknet_5_28_0_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_16 clkbuf_5_29_0_clk (.X(clknet_5_29_0_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_16 clkbuf_5_30_0_clk (.X(clknet_5_30_0_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_16 clkbuf_5_31_0_clk (.X(clknet_5_31_0_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_16 clkbuf_6_0_0_clk (.X(clknet_6_0_0_clk),
    .A(clknet_5_0_0_clk));
 sg13g2_buf_16 clkbuf_6_1_0_clk (.X(clknet_6_1_0_clk),
    .A(clknet_5_0_0_clk));
 sg13g2_buf_16 clkbuf_6_2_0_clk (.X(clknet_6_2_0_clk),
    .A(clknet_5_1_0_clk));
 sg13g2_buf_16 clkbuf_6_3_0_clk (.X(clknet_6_3_0_clk),
    .A(clknet_5_1_0_clk));
 sg13g2_buf_16 clkbuf_6_4_0_clk (.X(clknet_6_4_0_clk),
    .A(clknet_5_2_0_clk));
 sg13g2_buf_16 clkbuf_6_5_0_clk (.X(clknet_6_5_0_clk),
    .A(clknet_5_2_0_clk));
 sg13g2_buf_16 clkbuf_6_6_0_clk (.X(clknet_6_6_0_clk),
    .A(clknet_5_3_0_clk));
 sg13g2_buf_16 clkbuf_6_7_0_clk (.X(clknet_6_7_0_clk),
    .A(clknet_5_3_0_clk));
 sg13g2_buf_16 clkbuf_6_8_0_clk (.X(clknet_6_8_0_clk),
    .A(clknet_5_4_0_clk));
 sg13g2_buf_16 clkbuf_6_9_0_clk (.X(clknet_6_9_0_clk),
    .A(clknet_5_4_0_clk));
 sg13g2_buf_16 clkbuf_6_10_0_clk (.X(clknet_6_10_0_clk),
    .A(clknet_5_5_0_clk));
 sg13g2_buf_16 clkbuf_6_11_0_clk (.X(clknet_6_11_0_clk),
    .A(clknet_5_5_0_clk));
 sg13g2_buf_16 clkbuf_6_12_0_clk (.X(clknet_6_12_0_clk),
    .A(clknet_5_6_0_clk));
 sg13g2_buf_16 clkbuf_6_13_0_clk (.X(clknet_6_13_0_clk),
    .A(clknet_5_6_0_clk));
 sg13g2_buf_16 clkbuf_6_14_0_clk (.X(clknet_6_14_0_clk),
    .A(clknet_5_7_0_clk));
 sg13g2_buf_16 clkbuf_6_15_0_clk (.X(clknet_6_15_0_clk),
    .A(clknet_5_7_0_clk));
 sg13g2_buf_16 clkbuf_6_16_0_clk (.X(clknet_6_16_0_clk),
    .A(clknet_5_8_0_clk));
 sg13g2_buf_16 clkbuf_6_17_0_clk (.X(clknet_6_17_0_clk),
    .A(clknet_5_8_0_clk));
 sg13g2_buf_16 clkbuf_6_18_0_clk (.X(clknet_6_18_0_clk),
    .A(clknet_5_9_0_clk));
 sg13g2_buf_16 clkbuf_6_19_0_clk (.X(clknet_6_19_0_clk),
    .A(clknet_5_9_0_clk));
 sg13g2_buf_16 clkbuf_6_20_0_clk (.X(clknet_6_20_0_clk),
    .A(clknet_5_10_0_clk));
 sg13g2_buf_16 clkbuf_6_21_0_clk (.X(clknet_6_21_0_clk),
    .A(clknet_5_10_0_clk));
 sg13g2_buf_16 clkbuf_6_22_0_clk (.X(clknet_6_22_0_clk),
    .A(clknet_5_11_0_clk));
 sg13g2_buf_16 clkbuf_6_23_0_clk (.X(clknet_6_23_0_clk),
    .A(clknet_5_11_0_clk));
 sg13g2_buf_16 clkbuf_6_24_0_clk (.X(clknet_6_24_0_clk),
    .A(clknet_5_12_0_clk));
 sg13g2_buf_16 clkbuf_6_25_0_clk (.X(clknet_6_25_0_clk),
    .A(clknet_5_12_0_clk));
 sg13g2_buf_16 clkbuf_6_26_0_clk (.X(clknet_6_26_0_clk),
    .A(clknet_5_13_0_clk));
 sg13g2_buf_16 clkbuf_6_27_0_clk (.X(clknet_6_27_0_clk),
    .A(clknet_5_13_0_clk));
 sg13g2_buf_16 clkbuf_6_28_0_clk (.X(clknet_6_28_0_clk),
    .A(clknet_5_14_0_clk));
 sg13g2_buf_16 clkbuf_6_29_0_clk (.X(clknet_6_29_0_clk),
    .A(clknet_5_14_0_clk));
 sg13g2_buf_16 clkbuf_6_30_0_clk (.X(clknet_6_30_0_clk),
    .A(clknet_5_15_0_clk));
 sg13g2_buf_16 clkbuf_6_31_0_clk (.X(clknet_6_31_0_clk),
    .A(clknet_5_15_0_clk));
 sg13g2_buf_16 clkbuf_6_32_0_clk (.X(clknet_6_32_0_clk),
    .A(clknet_5_16_0_clk));
 sg13g2_buf_16 clkbuf_6_33_0_clk (.X(clknet_6_33_0_clk),
    .A(clknet_5_16_0_clk));
 sg13g2_buf_16 clkbuf_6_34_0_clk (.X(clknet_6_34_0_clk),
    .A(clknet_5_17_0_clk));
 sg13g2_buf_16 clkbuf_6_35_0_clk (.X(clknet_6_35_0_clk),
    .A(clknet_5_17_0_clk));
 sg13g2_buf_16 clkbuf_6_36_0_clk (.X(clknet_6_36_0_clk),
    .A(clknet_5_18_0_clk));
 sg13g2_buf_16 clkbuf_6_37_0_clk (.X(clknet_6_37_0_clk),
    .A(clknet_5_18_0_clk));
 sg13g2_buf_16 clkbuf_6_38_0_clk (.X(clknet_6_38_0_clk),
    .A(clknet_5_19_0_clk));
 sg13g2_buf_16 clkbuf_6_39_0_clk (.X(clknet_6_39_0_clk),
    .A(clknet_5_19_0_clk));
 sg13g2_buf_16 clkbuf_6_40_0_clk (.X(clknet_6_40_0_clk),
    .A(clknet_5_20_0_clk));
 sg13g2_buf_16 clkbuf_6_41_0_clk (.X(clknet_6_41_0_clk),
    .A(clknet_5_20_0_clk));
 sg13g2_buf_16 clkbuf_6_42_0_clk (.X(clknet_6_42_0_clk),
    .A(clknet_5_21_0_clk));
 sg13g2_buf_16 clkbuf_6_43_0_clk (.X(clknet_6_43_0_clk),
    .A(clknet_5_21_0_clk));
 sg13g2_buf_16 clkbuf_6_44_0_clk (.X(clknet_6_44_0_clk),
    .A(clknet_5_22_0_clk));
 sg13g2_buf_16 clkbuf_6_45_0_clk (.X(clknet_6_45_0_clk),
    .A(clknet_5_22_0_clk));
 sg13g2_buf_16 clkbuf_6_46_0_clk (.X(clknet_6_46_0_clk),
    .A(clknet_5_23_0_clk));
 sg13g2_buf_16 clkbuf_6_47_0_clk (.X(clknet_6_47_0_clk),
    .A(clknet_5_23_0_clk));
 sg13g2_buf_16 clkbuf_6_48_0_clk (.X(clknet_6_48_0_clk),
    .A(clknet_5_24_0_clk));
 sg13g2_buf_16 clkbuf_6_49_0_clk (.X(clknet_6_49_0_clk),
    .A(clknet_5_24_0_clk));
 sg13g2_buf_16 clkbuf_6_50_0_clk (.X(clknet_6_50_0_clk),
    .A(clknet_5_25_0_clk));
 sg13g2_buf_16 clkbuf_6_51_0_clk (.X(clknet_6_51_0_clk),
    .A(clknet_5_25_0_clk));
 sg13g2_buf_16 clkbuf_6_52_0_clk (.X(clknet_6_52_0_clk),
    .A(clknet_5_26_0_clk));
 sg13g2_buf_16 clkbuf_6_53_0_clk (.X(clknet_6_53_0_clk),
    .A(clknet_5_26_0_clk));
 sg13g2_buf_16 clkbuf_6_54_0_clk (.X(clknet_6_54_0_clk),
    .A(clknet_5_27_0_clk));
 sg13g2_buf_16 clkbuf_6_55_0_clk (.X(clknet_6_55_0_clk),
    .A(clknet_5_27_0_clk));
 sg13g2_buf_16 clkbuf_6_56_0_clk (.X(clknet_6_56_0_clk),
    .A(clknet_5_28_0_clk));
 sg13g2_buf_16 clkbuf_6_57_0_clk (.X(clknet_6_57_0_clk),
    .A(clknet_5_28_0_clk));
 sg13g2_buf_16 clkbuf_6_58_0_clk (.X(clknet_6_58_0_clk),
    .A(clknet_5_29_0_clk));
 sg13g2_buf_16 clkbuf_6_59_0_clk (.X(clknet_6_59_0_clk),
    .A(clknet_5_29_0_clk));
 sg13g2_buf_16 clkbuf_6_60_0_clk (.X(clknet_6_60_0_clk),
    .A(clknet_5_30_0_clk));
 sg13g2_buf_16 clkbuf_6_61_0_clk (.X(clknet_6_61_0_clk),
    .A(clknet_5_30_0_clk));
 sg13g2_buf_16 clkbuf_6_62_0_clk (.X(clknet_6_62_0_clk),
    .A(clknet_5_31_0_clk));
 sg13g2_buf_16 clkbuf_6_63_0_clk (.X(clknet_6_63_0_clk),
    .A(clknet_5_31_0_clk));
 sg13g2_buf_16 clkbuf_7_0_0_clk (.X(clknet_7_0_0_clk),
    .A(clknet_6_0_0_clk));
 sg13g2_buf_16 clkbuf_7_1_0_clk (.X(clknet_7_1_0_clk),
    .A(clknet_6_0_0_clk));
 sg13g2_buf_16 clkbuf_7_2_0_clk (.X(clknet_7_2_0_clk),
    .A(clknet_6_1_0_clk));
 sg13g2_buf_16 clkbuf_7_3_0_clk (.X(clknet_7_3_0_clk),
    .A(clknet_6_1_0_clk));
 sg13g2_buf_16 clkbuf_7_4_0_clk (.X(clknet_7_4_0_clk),
    .A(clknet_6_2_0_clk));
 sg13g2_buf_16 clkbuf_7_5_0_clk (.X(clknet_7_5_0_clk),
    .A(clknet_6_2_0_clk));
 sg13g2_buf_16 clkbuf_7_6_0_clk (.X(clknet_7_6_0_clk),
    .A(clknet_6_3_0_clk));
 sg13g2_buf_16 clkbuf_7_7_0_clk (.X(clknet_7_7_0_clk),
    .A(clknet_6_3_0_clk));
 sg13g2_buf_16 clkbuf_7_8_0_clk (.X(clknet_7_8_0_clk),
    .A(clknet_6_4_0_clk));
 sg13g2_buf_16 clkbuf_7_9_0_clk (.X(clknet_7_9_0_clk),
    .A(clknet_6_4_0_clk));
 sg13g2_buf_16 clkbuf_7_10_0_clk (.X(clknet_7_10_0_clk),
    .A(clknet_6_5_0_clk));
 sg13g2_buf_16 clkbuf_7_11_0_clk (.X(clknet_7_11_0_clk),
    .A(clknet_6_5_0_clk));
 sg13g2_buf_16 clkbuf_7_12_0_clk (.X(clknet_7_12_0_clk),
    .A(clknet_6_6_0_clk));
 sg13g2_buf_16 clkbuf_7_13_0_clk (.X(clknet_7_13_0_clk),
    .A(clknet_6_6_0_clk));
 sg13g2_buf_16 clkbuf_7_14_0_clk (.X(clknet_7_14_0_clk),
    .A(clknet_6_7_0_clk));
 sg13g2_buf_16 clkbuf_7_15_0_clk (.X(clknet_7_15_0_clk),
    .A(clknet_6_7_0_clk));
 sg13g2_buf_16 clkbuf_7_16_0_clk (.X(clknet_7_16_0_clk),
    .A(clknet_6_8_0_clk));
 sg13g2_buf_16 clkbuf_7_17_0_clk (.X(clknet_7_17_0_clk),
    .A(clknet_6_8_0_clk));
 sg13g2_buf_16 clkbuf_7_18_0_clk (.X(clknet_7_18_0_clk),
    .A(clknet_6_9_0_clk));
 sg13g2_buf_16 clkbuf_7_19_0_clk (.X(clknet_7_19_0_clk),
    .A(clknet_6_9_0_clk));
 sg13g2_buf_16 clkbuf_7_20_0_clk (.X(clknet_7_20_0_clk),
    .A(clknet_6_10_0_clk));
 sg13g2_buf_16 clkbuf_7_21_0_clk (.X(clknet_7_21_0_clk),
    .A(clknet_6_10_0_clk));
 sg13g2_buf_16 clkbuf_7_22_0_clk (.X(clknet_7_22_0_clk),
    .A(clknet_6_11_0_clk));
 sg13g2_buf_16 clkbuf_7_23_0_clk (.X(clknet_7_23_0_clk),
    .A(clknet_6_11_0_clk));
 sg13g2_buf_16 clkbuf_7_24_0_clk (.X(clknet_7_24_0_clk),
    .A(clknet_6_12_0_clk));
 sg13g2_buf_16 clkbuf_7_25_0_clk (.X(clknet_7_25_0_clk),
    .A(clknet_6_12_0_clk));
 sg13g2_buf_16 clkbuf_7_26_0_clk (.X(clknet_7_26_0_clk),
    .A(clknet_6_13_0_clk));
 sg13g2_buf_16 clkbuf_7_27_0_clk (.X(clknet_7_27_0_clk),
    .A(clknet_6_13_0_clk));
 sg13g2_buf_16 clkbuf_7_28_0_clk (.X(clknet_7_28_0_clk),
    .A(clknet_6_14_0_clk));
 sg13g2_buf_16 clkbuf_7_29_0_clk (.X(clknet_7_29_0_clk),
    .A(clknet_6_14_0_clk));
 sg13g2_buf_16 clkbuf_7_30_0_clk (.X(clknet_7_30_0_clk),
    .A(clknet_6_15_0_clk));
 sg13g2_buf_16 clkbuf_7_31_0_clk (.X(clknet_7_31_0_clk),
    .A(clknet_6_15_0_clk));
 sg13g2_buf_16 clkbuf_7_32_0_clk (.X(clknet_7_32_0_clk),
    .A(clknet_6_16_0_clk));
 sg13g2_buf_16 clkbuf_7_33_0_clk (.X(clknet_7_33_0_clk),
    .A(clknet_6_16_0_clk));
 sg13g2_buf_16 clkbuf_7_34_0_clk (.X(clknet_7_34_0_clk),
    .A(clknet_6_17_0_clk));
 sg13g2_buf_16 clkbuf_7_35_0_clk (.X(clknet_7_35_0_clk),
    .A(clknet_6_17_0_clk));
 sg13g2_buf_16 clkbuf_7_36_0_clk (.X(clknet_7_36_0_clk),
    .A(clknet_6_18_0_clk));
 sg13g2_buf_16 clkbuf_7_37_0_clk (.X(clknet_7_37_0_clk),
    .A(clknet_6_18_0_clk));
 sg13g2_buf_16 clkbuf_7_38_0_clk (.X(clknet_7_38_0_clk),
    .A(clknet_6_19_0_clk));
 sg13g2_buf_16 clkbuf_7_39_0_clk (.X(clknet_7_39_0_clk),
    .A(clknet_6_19_0_clk));
 sg13g2_buf_16 clkbuf_7_40_0_clk (.X(clknet_7_40_0_clk),
    .A(clknet_6_20_0_clk));
 sg13g2_buf_16 clkbuf_7_41_0_clk (.X(clknet_7_41_0_clk),
    .A(clknet_6_20_0_clk));
 sg13g2_buf_16 clkbuf_7_42_0_clk (.X(clknet_7_42_0_clk),
    .A(clknet_6_21_0_clk));
 sg13g2_buf_16 clkbuf_7_43_0_clk (.X(clknet_7_43_0_clk),
    .A(clknet_6_21_0_clk));
 sg13g2_buf_16 clkbuf_7_44_0_clk (.X(clknet_7_44_0_clk),
    .A(clknet_6_22_0_clk));
 sg13g2_buf_16 clkbuf_7_45_0_clk (.X(clknet_7_45_0_clk),
    .A(clknet_6_22_0_clk));
 sg13g2_buf_16 clkbuf_7_46_0_clk (.X(clknet_7_46_0_clk),
    .A(clknet_6_23_0_clk));
 sg13g2_buf_16 clkbuf_7_47_0_clk (.X(clknet_7_47_0_clk),
    .A(clknet_6_23_0_clk));
 sg13g2_buf_16 clkbuf_7_48_0_clk (.X(clknet_7_48_0_clk),
    .A(clknet_6_24_0_clk));
 sg13g2_buf_16 clkbuf_7_49_0_clk (.X(clknet_7_49_0_clk),
    .A(clknet_6_24_0_clk));
 sg13g2_buf_16 clkbuf_7_50_0_clk (.X(clknet_7_50_0_clk),
    .A(clknet_6_25_0_clk));
 sg13g2_buf_16 clkbuf_7_51_0_clk (.X(clknet_7_51_0_clk),
    .A(clknet_6_25_0_clk));
 sg13g2_buf_16 clkbuf_7_52_0_clk (.X(clknet_7_52_0_clk),
    .A(clknet_6_26_0_clk));
 sg13g2_buf_16 clkbuf_7_53_0_clk (.X(clknet_7_53_0_clk),
    .A(clknet_6_26_0_clk));
 sg13g2_buf_16 clkbuf_7_54_0_clk (.X(clknet_7_54_0_clk),
    .A(clknet_6_27_0_clk));
 sg13g2_buf_16 clkbuf_7_55_0_clk (.X(clknet_7_55_0_clk),
    .A(clknet_6_27_0_clk));
 sg13g2_buf_16 clkbuf_7_56_0_clk (.X(clknet_7_56_0_clk),
    .A(clknet_6_28_0_clk));
 sg13g2_buf_16 clkbuf_7_57_0_clk (.X(clknet_7_57_0_clk),
    .A(clknet_6_28_0_clk));
 sg13g2_buf_16 clkbuf_7_58_0_clk (.X(clknet_7_58_0_clk),
    .A(clknet_6_29_0_clk));
 sg13g2_buf_16 clkbuf_7_59_0_clk (.X(clknet_7_59_0_clk),
    .A(clknet_6_29_0_clk));
 sg13g2_buf_16 clkbuf_7_60_0_clk (.X(clknet_7_60_0_clk),
    .A(clknet_6_30_0_clk));
 sg13g2_buf_16 clkbuf_7_61_0_clk (.X(clknet_7_61_0_clk),
    .A(clknet_6_30_0_clk));
 sg13g2_buf_16 clkbuf_7_62_0_clk (.X(clknet_7_62_0_clk),
    .A(clknet_6_31_0_clk));
 sg13g2_buf_16 clkbuf_7_63_0_clk (.X(clknet_7_63_0_clk),
    .A(clknet_6_31_0_clk));
 sg13g2_buf_16 clkbuf_7_64_0_clk (.X(clknet_7_64_0_clk),
    .A(clknet_6_32_0_clk));
 sg13g2_buf_16 clkbuf_7_65_0_clk (.X(clknet_7_65_0_clk),
    .A(clknet_6_32_0_clk));
 sg13g2_buf_16 clkbuf_7_66_0_clk (.X(clknet_7_66_0_clk),
    .A(clknet_6_33_0_clk));
 sg13g2_buf_16 clkbuf_7_67_0_clk (.X(clknet_7_67_0_clk),
    .A(clknet_6_33_0_clk));
 sg13g2_buf_16 clkbuf_7_68_0_clk (.X(clknet_7_68_0_clk),
    .A(clknet_6_34_0_clk));
 sg13g2_buf_16 clkbuf_7_69_0_clk (.X(clknet_7_69_0_clk),
    .A(clknet_6_34_0_clk));
 sg13g2_buf_16 clkbuf_7_70_0_clk (.X(clknet_7_70_0_clk),
    .A(clknet_6_35_0_clk));
 sg13g2_buf_16 clkbuf_7_71_0_clk (.X(clknet_7_71_0_clk),
    .A(clknet_6_35_0_clk));
 sg13g2_buf_16 clkbuf_7_72_0_clk (.X(clknet_7_72_0_clk),
    .A(clknet_6_36_0_clk));
 sg13g2_buf_16 clkbuf_7_73_0_clk (.X(clknet_7_73_0_clk),
    .A(clknet_6_36_0_clk));
 sg13g2_buf_16 clkbuf_7_74_0_clk (.X(clknet_7_74_0_clk),
    .A(clknet_6_37_0_clk));
 sg13g2_buf_16 clkbuf_7_75_0_clk (.X(clknet_7_75_0_clk),
    .A(clknet_6_37_0_clk));
 sg13g2_buf_16 clkbuf_7_76_0_clk (.X(clknet_7_76_0_clk),
    .A(clknet_6_38_0_clk));
 sg13g2_buf_16 clkbuf_7_77_0_clk (.X(clknet_7_77_0_clk),
    .A(clknet_6_38_0_clk));
 sg13g2_buf_16 clkbuf_7_78_0_clk (.X(clknet_7_78_0_clk),
    .A(clknet_6_39_0_clk));
 sg13g2_buf_16 clkbuf_7_79_0_clk (.X(clknet_7_79_0_clk),
    .A(clknet_6_39_0_clk));
 sg13g2_buf_16 clkbuf_7_80_0_clk (.X(clknet_7_80_0_clk),
    .A(clknet_6_40_0_clk));
 sg13g2_buf_16 clkbuf_7_81_0_clk (.X(clknet_7_81_0_clk),
    .A(clknet_6_40_0_clk));
 sg13g2_buf_16 clkbuf_7_82_0_clk (.X(clknet_7_82_0_clk),
    .A(clknet_6_41_0_clk));
 sg13g2_buf_16 clkbuf_7_83_0_clk (.X(clknet_7_83_0_clk),
    .A(clknet_6_41_0_clk));
 sg13g2_buf_16 clkbuf_7_84_0_clk (.X(clknet_7_84_0_clk),
    .A(clknet_6_42_0_clk));
 sg13g2_buf_16 clkbuf_7_85_0_clk (.X(clknet_7_85_0_clk),
    .A(clknet_6_42_0_clk));
 sg13g2_buf_16 clkbuf_7_86_0_clk (.X(clknet_7_86_0_clk),
    .A(clknet_6_43_0_clk));
 sg13g2_buf_16 clkbuf_7_87_0_clk (.X(clknet_7_87_0_clk),
    .A(clknet_6_43_0_clk));
 sg13g2_buf_16 clkbuf_7_88_0_clk (.X(clknet_7_88_0_clk),
    .A(clknet_6_44_0_clk));
 sg13g2_buf_16 clkbuf_7_89_0_clk (.X(clknet_7_89_0_clk),
    .A(clknet_6_44_0_clk));
 sg13g2_buf_16 clkbuf_7_90_0_clk (.X(clknet_7_90_0_clk),
    .A(clknet_6_45_0_clk));
 sg13g2_buf_16 clkbuf_7_91_0_clk (.X(clknet_7_91_0_clk),
    .A(clknet_6_45_0_clk));
 sg13g2_buf_16 clkbuf_7_92_0_clk (.X(clknet_7_92_0_clk),
    .A(clknet_6_46_0_clk));
 sg13g2_buf_16 clkbuf_7_93_0_clk (.X(clknet_7_93_0_clk),
    .A(clknet_6_46_0_clk));
 sg13g2_buf_16 clkbuf_7_94_0_clk (.X(clknet_7_94_0_clk),
    .A(clknet_6_47_0_clk));
 sg13g2_buf_16 clkbuf_7_95_0_clk (.X(clknet_7_95_0_clk),
    .A(clknet_6_47_0_clk));
 sg13g2_buf_16 clkbuf_7_96_0_clk (.X(clknet_7_96_0_clk),
    .A(clknet_6_48_0_clk));
 sg13g2_buf_16 clkbuf_7_97_0_clk (.X(clknet_7_97_0_clk),
    .A(clknet_6_48_0_clk));
 sg13g2_buf_16 clkbuf_7_98_0_clk (.X(clknet_7_98_0_clk),
    .A(clknet_6_49_0_clk));
 sg13g2_buf_16 clkbuf_7_99_0_clk (.X(clknet_7_99_0_clk),
    .A(clknet_6_49_0_clk));
 sg13g2_buf_16 clkbuf_7_100_0_clk (.X(clknet_7_100_0_clk),
    .A(clknet_6_50_0_clk));
 sg13g2_buf_16 clkbuf_7_101_0_clk (.X(clknet_7_101_0_clk),
    .A(clknet_6_50_0_clk));
 sg13g2_buf_16 clkbuf_7_102_0_clk (.X(clknet_7_102_0_clk),
    .A(clknet_6_51_0_clk));
 sg13g2_buf_16 clkbuf_7_103_0_clk (.X(clknet_7_103_0_clk),
    .A(clknet_6_51_0_clk));
 sg13g2_buf_16 clkbuf_7_104_0_clk (.X(clknet_7_104_0_clk),
    .A(clknet_6_52_0_clk));
 sg13g2_buf_16 clkbuf_7_105_0_clk (.X(clknet_7_105_0_clk),
    .A(clknet_6_52_0_clk));
 sg13g2_buf_16 clkbuf_7_106_0_clk (.X(clknet_7_106_0_clk),
    .A(clknet_6_53_0_clk));
 sg13g2_buf_16 clkbuf_7_107_0_clk (.X(clknet_7_107_0_clk),
    .A(clknet_6_53_0_clk));
 sg13g2_buf_16 clkbuf_7_108_0_clk (.X(clknet_7_108_0_clk),
    .A(clknet_6_54_0_clk));
 sg13g2_buf_16 clkbuf_7_109_0_clk (.X(clknet_7_109_0_clk),
    .A(clknet_6_54_0_clk));
 sg13g2_buf_16 clkbuf_7_110_0_clk (.X(clknet_7_110_0_clk),
    .A(clknet_6_55_0_clk));
 sg13g2_buf_16 clkbuf_7_111_0_clk (.X(clknet_7_111_0_clk),
    .A(clknet_6_55_0_clk));
 sg13g2_buf_16 clkbuf_7_112_0_clk (.X(clknet_7_112_0_clk),
    .A(clknet_6_56_0_clk));
 sg13g2_buf_16 clkbuf_7_113_0_clk (.X(clknet_7_113_0_clk),
    .A(clknet_6_56_0_clk));
 sg13g2_buf_16 clkbuf_7_114_0_clk (.X(clknet_7_114_0_clk),
    .A(clknet_6_57_0_clk));
 sg13g2_buf_16 clkbuf_7_115_0_clk (.X(clknet_7_115_0_clk),
    .A(clknet_6_57_0_clk));
 sg13g2_buf_16 clkbuf_7_116_0_clk (.X(clknet_7_116_0_clk),
    .A(clknet_6_58_0_clk));
 sg13g2_buf_16 clkbuf_7_117_0_clk (.X(clknet_7_117_0_clk),
    .A(clknet_6_58_0_clk));
 sg13g2_buf_16 clkbuf_7_118_0_clk (.X(clknet_7_118_0_clk),
    .A(clknet_6_59_0_clk));
 sg13g2_buf_16 clkbuf_7_119_0_clk (.X(clknet_7_119_0_clk),
    .A(clknet_6_59_0_clk));
 sg13g2_buf_16 clkbuf_7_120_0_clk (.X(clknet_7_120_0_clk),
    .A(clknet_6_60_0_clk));
 sg13g2_buf_16 clkbuf_7_121_0_clk (.X(clknet_7_121_0_clk),
    .A(clknet_6_60_0_clk));
 sg13g2_buf_16 clkbuf_7_122_0_clk (.X(clknet_7_122_0_clk),
    .A(clknet_6_61_0_clk));
 sg13g2_buf_16 clkbuf_7_123_0_clk (.X(clknet_7_123_0_clk),
    .A(clknet_6_61_0_clk));
 sg13g2_buf_16 clkbuf_7_124_0_clk (.X(clknet_7_124_0_clk),
    .A(clknet_6_62_0_clk));
 sg13g2_buf_16 clkbuf_7_125_0_clk (.X(clknet_7_125_0_clk),
    .A(clknet_6_62_0_clk));
 sg13g2_buf_16 clkbuf_7_126_0_clk (.X(clknet_7_126_0_clk),
    .A(clknet_6_63_0_clk));
 sg13g2_buf_16 clkbuf_7_127_0_clk (.X(clknet_7_127_0_clk),
    .A(clknet_6_63_0_clk));
 sg13g2_buf_16 clkbuf_8_0_0_clk (.X(clknet_8_0_0_clk),
    .A(clknet_7_0_0_clk));
 sg13g2_buf_16 clkbuf_8_1_0_clk (.X(clknet_8_1_0_clk),
    .A(clknet_7_0_0_clk));
 sg13g2_buf_16 clkbuf_8_2_0_clk (.X(clknet_8_2_0_clk),
    .A(clknet_7_1_0_clk));
 sg13g2_buf_16 clkbuf_8_3_0_clk (.X(clknet_8_3_0_clk),
    .A(clknet_7_1_0_clk));
 sg13g2_buf_16 clkbuf_8_4_0_clk (.X(clknet_8_4_0_clk),
    .A(clknet_7_2_0_clk));
 sg13g2_buf_16 clkbuf_8_5_0_clk (.X(clknet_8_5_0_clk),
    .A(clknet_7_2_0_clk));
 sg13g2_buf_16 clkbuf_8_6_0_clk (.X(clknet_8_6_0_clk),
    .A(clknet_7_3_0_clk));
 sg13g2_buf_16 clkbuf_8_7_0_clk (.X(clknet_8_7_0_clk),
    .A(clknet_7_3_0_clk));
 sg13g2_buf_16 clkbuf_8_8_0_clk (.X(clknet_8_8_0_clk),
    .A(clknet_7_4_0_clk));
 sg13g2_buf_16 clkbuf_8_9_0_clk (.X(clknet_8_9_0_clk),
    .A(clknet_7_4_0_clk));
 sg13g2_buf_16 clkbuf_8_10_0_clk (.X(clknet_8_10_0_clk),
    .A(clknet_7_5_0_clk));
 sg13g2_buf_16 clkbuf_8_11_0_clk (.X(clknet_8_11_0_clk),
    .A(clknet_7_5_0_clk));
 sg13g2_buf_16 clkbuf_8_12_0_clk (.X(clknet_8_12_0_clk),
    .A(clknet_7_6_0_clk));
 sg13g2_buf_16 clkbuf_8_13_0_clk (.X(clknet_8_13_0_clk),
    .A(clknet_7_6_0_clk));
 sg13g2_buf_16 clkbuf_8_14_0_clk (.X(clknet_8_14_0_clk),
    .A(clknet_7_7_0_clk));
 sg13g2_buf_16 clkbuf_8_15_0_clk (.X(clknet_8_15_0_clk),
    .A(clknet_7_7_0_clk));
 sg13g2_buf_16 clkbuf_8_16_0_clk (.X(clknet_8_16_0_clk),
    .A(clknet_7_8_0_clk));
 sg13g2_buf_16 clkbuf_8_17_0_clk (.X(clknet_8_17_0_clk),
    .A(clknet_7_8_0_clk));
 sg13g2_buf_16 clkbuf_8_18_0_clk (.X(clknet_8_18_0_clk),
    .A(clknet_7_9_0_clk));
 sg13g2_buf_16 clkbuf_8_19_0_clk (.X(clknet_8_19_0_clk),
    .A(clknet_7_9_0_clk));
 sg13g2_buf_16 clkbuf_8_20_0_clk (.X(clknet_8_20_0_clk),
    .A(clknet_7_10_0_clk));
 sg13g2_buf_16 clkbuf_8_21_0_clk (.X(clknet_8_21_0_clk),
    .A(clknet_7_10_0_clk));
 sg13g2_buf_16 clkbuf_8_22_0_clk (.X(clknet_8_22_0_clk),
    .A(clknet_7_11_0_clk));
 sg13g2_buf_16 clkbuf_8_23_0_clk (.X(clknet_8_23_0_clk),
    .A(clknet_7_11_0_clk));
 sg13g2_buf_16 clkbuf_8_24_0_clk (.X(clknet_8_24_0_clk),
    .A(clknet_7_12_0_clk));
 sg13g2_buf_16 clkbuf_8_25_0_clk (.X(clknet_8_25_0_clk),
    .A(clknet_7_12_0_clk));
 sg13g2_buf_16 clkbuf_8_26_0_clk (.X(clknet_8_26_0_clk),
    .A(clknet_7_13_0_clk));
 sg13g2_buf_16 clkbuf_8_27_0_clk (.X(clknet_8_27_0_clk),
    .A(clknet_7_13_0_clk));
 sg13g2_buf_16 clkbuf_8_28_0_clk (.X(clknet_8_28_0_clk),
    .A(clknet_7_14_0_clk));
 sg13g2_buf_16 clkbuf_8_29_0_clk (.X(clknet_8_29_0_clk),
    .A(clknet_7_14_0_clk));
 sg13g2_buf_16 clkbuf_8_30_0_clk (.X(clknet_8_30_0_clk),
    .A(clknet_7_15_0_clk));
 sg13g2_buf_16 clkbuf_8_31_0_clk (.X(clknet_8_31_0_clk),
    .A(clknet_7_15_0_clk));
 sg13g2_buf_16 clkbuf_8_32_0_clk (.X(clknet_8_32_0_clk),
    .A(clknet_7_16_0_clk));
 sg13g2_buf_16 clkbuf_8_33_0_clk (.X(clknet_8_33_0_clk),
    .A(clknet_7_16_0_clk));
 sg13g2_buf_16 clkbuf_8_34_0_clk (.X(clknet_8_34_0_clk),
    .A(clknet_7_17_0_clk));
 sg13g2_buf_16 clkbuf_8_35_0_clk (.X(clknet_8_35_0_clk),
    .A(clknet_7_17_0_clk));
 sg13g2_buf_16 clkbuf_8_36_0_clk (.X(clknet_8_36_0_clk),
    .A(clknet_7_18_0_clk));
 sg13g2_buf_16 clkbuf_8_37_0_clk (.X(clknet_8_37_0_clk),
    .A(clknet_7_18_0_clk));
 sg13g2_buf_16 clkbuf_8_38_0_clk (.X(clknet_8_38_0_clk),
    .A(clknet_7_19_0_clk));
 sg13g2_buf_16 clkbuf_8_39_0_clk (.X(clknet_8_39_0_clk),
    .A(clknet_7_19_0_clk));
 sg13g2_buf_16 clkbuf_8_40_0_clk (.X(clknet_8_40_0_clk),
    .A(clknet_7_20_0_clk));
 sg13g2_buf_16 clkbuf_8_41_0_clk (.X(clknet_8_41_0_clk),
    .A(clknet_7_20_0_clk));
 sg13g2_buf_16 clkbuf_8_42_0_clk (.X(clknet_8_42_0_clk),
    .A(clknet_7_21_0_clk));
 sg13g2_buf_16 clkbuf_8_43_0_clk (.X(clknet_8_43_0_clk),
    .A(clknet_7_21_0_clk));
 sg13g2_buf_16 clkbuf_8_44_0_clk (.X(clknet_8_44_0_clk),
    .A(clknet_7_22_0_clk));
 sg13g2_buf_16 clkbuf_8_45_0_clk (.X(clknet_8_45_0_clk),
    .A(clknet_7_22_0_clk));
 sg13g2_buf_16 clkbuf_8_46_0_clk (.X(clknet_8_46_0_clk),
    .A(clknet_7_23_0_clk));
 sg13g2_buf_16 clkbuf_8_47_0_clk (.X(clknet_8_47_0_clk),
    .A(clknet_7_23_0_clk));
 sg13g2_buf_16 clkbuf_8_48_0_clk (.X(clknet_8_48_0_clk),
    .A(clknet_7_24_0_clk));
 sg13g2_buf_16 clkbuf_8_49_0_clk (.X(clknet_8_49_0_clk),
    .A(clknet_7_24_0_clk));
 sg13g2_buf_16 clkbuf_8_50_0_clk (.X(clknet_8_50_0_clk),
    .A(clknet_7_25_0_clk));
 sg13g2_buf_16 clkbuf_8_51_0_clk (.X(clknet_8_51_0_clk),
    .A(clknet_7_25_0_clk));
 sg13g2_buf_16 clkbuf_8_52_0_clk (.X(clknet_8_52_0_clk),
    .A(clknet_7_26_0_clk));
 sg13g2_buf_16 clkbuf_8_53_0_clk (.X(clknet_8_53_0_clk),
    .A(clknet_7_26_0_clk));
 sg13g2_buf_16 clkbuf_8_54_0_clk (.X(clknet_8_54_0_clk),
    .A(clknet_7_27_0_clk));
 sg13g2_buf_16 clkbuf_8_55_0_clk (.X(clknet_8_55_0_clk),
    .A(clknet_7_27_0_clk));
 sg13g2_buf_16 clkbuf_8_56_0_clk (.X(clknet_8_56_0_clk),
    .A(clknet_7_28_0_clk));
 sg13g2_buf_16 clkbuf_8_57_0_clk (.X(clknet_8_57_0_clk),
    .A(clknet_7_28_0_clk));
 sg13g2_buf_16 clkbuf_8_58_0_clk (.X(clknet_8_58_0_clk),
    .A(clknet_7_29_0_clk));
 sg13g2_buf_16 clkbuf_8_59_0_clk (.X(clknet_8_59_0_clk),
    .A(clknet_7_29_0_clk));
 sg13g2_buf_16 clkbuf_8_60_0_clk (.X(clknet_8_60_0_clk),
    .A(clknet_7_30_0_clk));
 sg13g2_buf_16 clkbuf_8_61_0_clk (.X(clknet_8_61_0_clk),
    .A(clknet_7_30_0_clk));
 sg13g2_buf_16 clkbuf_8_62_0_clk (.X(clknet_8_62_0_clk),
    .A(clknet_7_31_0_clk));
 sg13g2_buf_16 clkbuf_8_63_0_clk (.X(clknet_8_63_0_clk),
    .A(clknet_7_31_0_clk));
 sg13g2_buf_16 clkbuf_8_64_0_clk (.X(clknet_8_64_0_clk),
    .A(clknet_7_32_0_clk));
 sg13g2_buf_16 clkbuf_8_65_0_clk (.X(clknet_8_65_0_clk),
    .A(clknet_7_32_0_clk));
 sg13g2_buf_16 clkbuf_8_66_0_clk (.X(clknet_8_66_0_clk),
    .A(clknet_7_33_0_clk));
 sg13g2_buf_16 clkbuf_8_67_0_clk (.X(clknet_8_67_0_clk),
    .A(clknet_7_33_0_clk));
 sg13g2_buf_16 clkbuf_8_68_0_clk (.X(clknet_8_68_0_clk),
    .A(clknet_7_34_0_clk));
 sg13g2_buf_16 clkbuf_8_69_0_clk (.X(clknet_8_69_0_clk),
    .A(clknet_7_34_0_clk));
 sg13g2_buf_16 clkbuf_8_70_0_clk (.X(clknet_8_70_0_clk),
    .A(clknet_7_35_0_clk));
 sg13g2_buf_16 clkbuf_8_71_0_clk (.X(clknet_8_71_0_clk),
    .A(clknet_7_35_0_clk));
 sg13g2_buf_16 clkbuf_8_72_0_clk (.X(clknet_8_72_0_clk),
    .A(clknet_7_36_0_clk));
 sg13g2_buf_16 clkbuf_8_73_0_clk (.X(clknet_8_73_0_clk),
    .A(clknet_7_36_0_clk));
 sg13g2_buf_16 clkbuf_8_74_0_clk (.X(clknet_8_74_0_clk),
    .A(clknet_7_37_0_clk));
 sg13g2_buf_16 clkbuf_8_75_0_clk (.X(clknet_8_75_0_clk),
    .A(clknet_7_37_0_clk));
 sg13g2_buf_16 clkbuf_8_76_0_clk (.X(clknet_8_76_0_clk),
    .A(clknet_7_38_0_clk));
 sg13g2_buf_16 clkbuf_8_77_0_clk (.X(clknet_8_77_0_clk),
    .A(clknet_7_38_0_clk));
 sg13g2_buf_16 clkbuf_8_78_0_clk (.X(clknet_8_78_0_clk),
    .A(clknet_7_39_0_clk));
 sg13g2_buf_16 clkbuf_8_79_0_clk (.X(clknet_8_79_0_clk),
    .A(clknet_7_39_0_clk));
 sg13g2_buf_16 clkbuf_8_80_0_clk (.X(clknet_8_80_0_clk),
    .A(clknet_7_40_0_clk));
 sg13g2_buf_16 clkbuf_8_81_0_clk (.X(clknet_8_81_0_clk),
    .A(clknet_7_40_0_clk));
 sg13g2_buf_16 clkbuf_8_82_0_clk (.X(clknet_8_82_0_clk),
    .A(clknet_7_41_0_clk));
 sg13g2_buf_16 clkbuf_8_83_0_clk (.X(clknet_8_83_0_clk),
    .A(clknet_7_41_0_clk));
 sg13g2_buf_16 clkbuf_8_84_0_clk (.X(clknet_8_84_0_clk),
    .A(clknet_7_42_0_clk));
 sg13g2_buf_16 clkbuf_8_85_0_clk (.X(clknet_8_85_0_clk),
    .A(clknet_7_42_0_clk));
 sg13g2_buf_16 clkbuf_8_86_0_clk (.X(clknet_8_86_0_clk),
    .A(clknet_7_43_0_clk));
 sg13g2_buf_16 clkbuf_8_87_0_clk (.X(clknet_8_87_0_clk),
    .A(clknet_7_43_0_clk));
 sg13g2_buf_16 clkbuf_8_88_0_clk (.X(clknet_8_88_0_clk),
    .A(clknet_7_44_0_clk));
 sg13g2_buf_16 clkbuf_8_89_0_clk (.X(clknet_8_89_0_clk),
    .A(clknet_7_44_0_clk));
 sg13g2_buf_16 clkbuf_8_90_0_clk (.X(clknet_8_90_0_clk),
    .A(clknet_7_45_0_clk));
 sg13g2_buf_16 clkbuf_8_91_0_clk (.X(clknet_8_91_0_clk),
    .A(clknet_7_45_0_clk));
 sg13g2_buf_16 clkbuf_8_92_0_clk (.X(clknet_8_92_0_clk),
    .A(clknet_7_46_0_clk));
 sg13g2_buf_16 clkbuf_8_93_0_clk (.X(clknet_8_93_0_clk),
    .A(clknet_7_46_0_clk));
 sg13g2_buf_16 clkbuf_8_94_0_clk (.X(clknet_8_94_0_clk),
    .A(clknet_7_47_0_clk));
 sg13g2_buf_16 clkbuf_8_95_0_clk (.X(clknet_8_95_0_clk),
    .A(clknet_7_47_0_clk));
 sg13g2_buf_16 clkbuf_8_96_0_clk (.X(clknet_8_96_0_clk),
    .A(clknet_7_48_0_clk));
 sg13g2_buf_16 clkbuf_8_97_0_clk (.X(clknet_8_97_0_clk),
    .A(clknet_7_48_0_clk));
 sg13g2_buf_16 clkbuf_8_98_0_clk (.X(clknet_8_98_0_clk),
    .A(clknet_7_49_0_clk));
 sg13g2_buf_16 clkbuf_8_99_0_clk (.X(clknet_8_99_0_clk),
    .A(clknet_7_49_0_clk));
 sg13g2_buf_16 clkbuf_8_100_0_clk (.X(clknet_8_100_0_clk),
    .A(clknet_7_50_0_clk));
 sg13g2_buf_16 clkbuf_8_101_0_clk (.X(clknet_8_101_0_clk),
    .A(clknet_7_50_0_clk));
 sg13g2_buf_16 clkbuf_8_102_0_clk (.X(clknet_8_102_0_clk),
    .A(clknet_7_51_0_clk));
 sg13g2_buf_16 clkbuf_8_103_0_clk (.X(clknet_8_103_0_clk),
    .A(clknet_7_51_0_clk));
 sg13g2_buf_16 clkbuf_8_104_0_clk (.X(clknet_8_104_0_clk),
    .A(clknet_7_52_0_clk));
 sg13g2_buf_16 clkbuf_8_105_0_clk (.X(clknet_8_105_0_clk),
    .A(clknet_7_52_0_clk));
 sg13g2_buf_16 clkbuf_8_106_0_clk (.X(clknet_8_106_0_clk),
    .A(clknet_7_53_0_clk));
 sg13g2_buf_16 clkbuf_8_107_0_clk (.X(clknet_8_107_0_clk),
    .A(clknet_7_53_0_clk));
 sg13g2_buf_16 clkbuf_8_108_0_clk (.X(clknet_8_108_0_clk),
    .A(clknet_7_54_0_clk));
 sg13g2_buf_16 clkbuf_8_109_0_clk (.X(clknet_8_109_0_clk),
    .A(clknet_7_54_0_clk));
 sg13g2_buf_16 clkbuf_8_110_0_clk (.X(clknet_8_110_0_clk),
    .A(clknet_7_55_0_clk));
 sg13g2_buf_16 clkbuf_8_111_0_clk (.X(clknet_8_111_0_clk),
    .A(clknet_7_55_0_clk));
 sg13g2_buf_16 clkbuf_8_112_0_clk (.X(clknet_8_112_0_clk),
    .A(clknet_7_56_0_clk));
 sg13g2_buf_16 clkbuf_8_113_0_clk (.X(clknet_8_113_0_clk),
    .A(clknet_7_56_0_clk));
 sg13g2_buf_16 clkbuf_8_114_0_clk (.X(clknet_8_114_0_clk),
    .A(clknet_7_57_0_clk));
 sg13g2_buf_16 clkbuf_8_115_0_clk (.X(clknet_8_115_0_clk),
    .A(clknet_7_57_0_clk));
 sg13g2_buf_16 clkbuf_8_116_0_clk (.X(clknet_8_116_0_clk),
    .A(clknet_7_58_0_clk));
 sg13g2_buf_16 clkbuf_8_117_0_clk (.X(clknet_8_117_0_clk),
    .A(clknet_7_58_0_clk));
 sg13g2_buf_16 clkbuf_8_118_0_clk (.X(clknet_8_118_0_clk),
    .A(clknet_7_59_0_clk));
 sg13g2_buf_16 clkbuf_8_119_0_clk (.X(clknet_8_119_0_clk),
    .A(clknet_7_59_0_clk));
 sg13g2_buf_16 clkbuf_8_120_0_clk (.X(clknet_8_120_0_clk),
    .A(clknet_7_60_0_clk));
 sg13g2_buf_16 clkbuf_8_121_0_clk (.X(clknet_8_121_0_clk),
    .A(clknet_7_60_0_clk));
 sg13g2_buf_16 clkbuf_8_122_0_clk (.X(clknet_8_122_0_clk),
    .A(clknet_7_61_0_clk));
 sg13g2_buf_16 clkbuf_8_123_0_clk (.X(clknet_8_123_0_clk),
    .A(clknet_7_61_0_clk));
 sg13g2_buf_16 clkbuf_8_124_0_clk (.X(clknet_8_124_0_clk),
    .A(clknet_7_62_0_clk));
 sg13g2_buf_16 clkbuf_8_125_0_clk (.X(clknet_8_125_0_clk),
    .A(clknet_7_62_0_clk));
 sg13g2_buf_16 clkbuf_8_126_0_clk (.X(clknet_8_126_0_clk),
    .A(clknet_7_63_0_clk));
 sg13g2_buf_16 clkbuf_8_127_0_clk (.X(clknet_8_127_0_clk),
    .A(clknet_7_63_0_clk));
 sg13g2_buf_16 clkbuf_8_128_0_clk (.X(clknet_8_128_0_clk),
    .A(clknet_7_64_0_clk));
 sg13g2_buf_16 clkbuf_8_129_0_clk (.X(clknet_8_129_0_clk),
    .A(clknet_7_64_0_clk));
 sg13g2_buf_16 clkbuf_8_130_0_clk (.X(clknet_8_130_0_clk),
    .A(clknet_7_65_0_clk));
 sg13g2_buf_16 clkbuf_8_131_0_clk (.X(clknet_8_131_0_clk),
    .A(clknet_7_65_0_clk));
 sg13g2_buf_16 clkbuf_8_132_0_clk (.X(clknet_8_132_0_clk),
    .A(clknet_7_66_0_clk));
 sg13g2_buf_16 clkbuf_8_133_0_clk (.X(clknet_8_133_0_clk),
    .A(clknet_7_66_0_clk));
 sg13g2_buf_16 clkbuf_8_134_0_clk (.X(clknet_8_134_0_clk),
    .A(clknet_7_67_0_clk));
 sg13g2_buf_16 clkbuf_8_135_0_clk (.X(clknet_8_135_0_clk),
    .A(clknet_7_67_0_clk));
 sg13g2_buf_16 clkbuf_8_136_0_clk (.X(clknet_8_136_0_clk),
    .A(clknet_7_68_0_clk));
 sg13g2_buf_16 clkbuf_8_137_0_clk (.X(clknet_8_137_0_clk),
    .A(clknet_7_68_0_clk));
 sg13g2_buf_16 clkbuf_8_138_0_clk (.X(clknet_8_138_0_clk),
    .A(clknet_7_69_0_clk));
 sg13g2_buf_16 clkbuf_8_139_0_clk (.X(clknet_8_139_0_clk),
    .A(clknet_7_69_0_clk));
 sg13g2_buf_16 clkbuf_8_140_0_clk (.X(clknet_8_140_0_clk),
    .A(clknet_7_70_0_clk));
 sg13g2_buf_16 clkbuf_8_141_0_clk (.X(clknet_8_141_0_clk),
    .A(clknet_7_70_0_clk));
 sg13g2_buf_16 clkbuf_8_142_0_clk (.X(clknet_8_142_0_clk),
    .A(clknet_7_71_0_clk));
 sg13g2_buf_16 clkbuf_8_143_0_clk (.X(clknet_8_143_0_clk),
    .A(clknet_7_71_0_clk));
 sg13g2_buf_16 clkbuf_8_144_0_clk (.X(clknet_8_144_0_clk),
    .A(clknet_7_72_0_clk));
 sg13g2_buf_16 clkbuf_8_145_0_clk (.X(clknet_8_145_0_clk),
    .A(clknet_7_72_0_clk));
 sg13g2_buf_16 clkbuf_8_146_0_clk (.X(clknet_8_146_0_clk),
    .A(clknet_7_73_0_clk));
 sg13g2_buf_16 clkbuf_8_147_0_clk (.X(clknet_8_147_0_clk),
    .A(clknet_7_73_0_clk));
 sg13g2_buf_16 clkbuf_8_148_0_clk (.X(clknet_8_148_0_clk),
    .A(clknet_7_74_0_clk));
 sg13g2_buf_16 clkbuf_8_149_0_clk (.X(clknet_8_149_0_clk),
    .A(clknet_7_74_0_clk));
 sg13g2_buf_16 clkbuf_8_150_0_clk (.X(clknet_8_150_0_clk),
    .A(clknet_7_75_0_clk));
 sg13g2_buf_16 clkbuf_8_151_0_clk (.X(clknet_8_151_0_clk),
    .A(clknet_7_75_0_clk));
 sg13g2_buf_16 clkbuf_8_152_0_clk (.X(clknet_8_152_0_clk),
    .A(clknet_7_76_0_clk));
 sg13g2_buf_16 clkbuf_8_153_0_clk (.X(clknet_8_153_0_clk),
    .A(clknet_7_76_0_clk));
 sg13g2_buf_16 clkbuf_8_154_0_clk (.X(clknet_8_154_0_clk),
    .A(clknet_7_77_0_clk));
 sg13g2_buf_16 clkbuf_8_155_0_clk (.X(clknet_8_155_0_clk),
    .A(clknet_7_77_0_clk));
 sg13g2_buf_16 clkbuf_8_156_0_clk (.X(clknet_8_156_0_clk),
    .A(clknet_7_78_0_clk));
 sg13g2_buf_16 clkbuf_8_157_0_clk (.X(clknet_8_157_0_clk),
    .A(clknet_7_78_0_clk));
 sg13g2_buf_16 clkbuf_8_158_0_clk (.X(clknet_8_158_0_clk),
    .A(clknet_7_79_0_clk));
 sg13g2_buf_16 clkbuf_8_159_0_clk (.X(clknet_8_159_0_clk),
    .A(clknet_7_79_0_clk));
 sg13g2_buf_16 clkbuf_8_160_0_clk (.X(clknet_8_160_0_clk),
    .A(clknet_7_80_0_clk));
 sg13g2_buf_16 clkbuf_8_161_0_clk (.X(clknet_8_161_0_clk),
    .A(clknet_7_80_0_clk));
 sg13g2_buf_16 clkbuf_8_162_0_clk (.X(clknet_8_162_0_clk),
    .A(clknet_7_81_0_clk));
 sg13g2_buf_16 clkbuf_8_163_0_clk (.X(clknet_8_163_0_clk),
    .A(clknet_7_81_0_clk));
 sg13g2_buf_16 clkbuf_8_164_0_clk (.X(clknet_8_164_0_clk),
    .A(clknet_7_82_0_clk));
 sg13g2_buf_16 clkbuf_8_165_0_clk (.X(clknet_8_165_0_clk),
    .A(clknet_7_82_0_clk));
 sg13g2_buf_16 clkbuf_8_166_0_clk (.X(clknet_8_166_0_clk),
    .A(clknet_7_83_0_clk));
 sg13g2_buf_16 clkbuf_8_167_0_clk (.X(clknet_8_167_0_clk),
    .A(clknet_7_83_0_clk));
 sg13g2_buf_16 clkbuf_8_168_0_clk (.X(clknet_8_168_0_clk),
    .A(clknet_7_84_0_clk));
 sg13g2_buf_16 clkbuf_8_169_0_clk (.X(clknet_8_169_0_clk),
    .A(clknet_7_84_0_clk));
 sg13g2_buf_16 clkbuf_8_170_0_clk (.X(clknet_8_170_0_clk),
    .A(clknet_7_85_0_clk));
 sg13g2_buf_16 clkbuf_8_171_0_clk (.X(clknet_8_171_0_clk),
    .A(clknet_7_85_0_clk));
 sg13g2_buf_16 clkbuf_8_172_0_clk (.X(clknet_8_172_0_clk),
    .A(clknet_7_86_0_clk));
 sg13g2_buf_16 clkbuf_8_173_0_clk (.X(clknet_8_173_0_clk),
    .A(clknet_7_86_0_clk));
 sg13g2_buf_16 clkbuf_8_174_0_clk (.X(clknet_8_174_0_clk),
    .A(clknet_7_87_0_clk));
 sg13g2_buf_16 clkbuf_8_175_0_clk (.X(clknet_8_175_0_clk),
    .A(clknet_7_87_0_clk));
 sg13g2_buf_16 clkbuf_8_176_0_clk (.X(clknet_8_176_0_clk),
    .A(clknet_7_88_0_clk));
 sg13g2_buf_16 clkbuf_8_177_0_clk (.X(clknet_8_177_0_clk),
    .A(clknet_7_88_0_clk));
 sg13g2_buf_16 clkbuf_8_178_0_clk (.X(clknet_8_178_0_clk),
    .A(clknet_7_89_0_clk));
 sg13g2_buf_16 clkbuf_8_179_0_clk (.X(clknet_8_179_0_clk),
    .A(clknet_7_89_0_clk));
 sg13g2_buf_16 clkbuf_8_180_0_clk (.X(clknet_8_180_0_clk),
    .A(clknet_7_90_0_clk));
 sg13g2_buf_16 clkbuf_8_181_0_clk (.X(clknet_8_181_0_clk),
    .A(clknet_7_90_0_clk));
 sg13g2_buf_16 clkbuf_8_182_0_clk (.X(clknet_8_182_0_clk),
    .A(clknet_7_91_0_clk));
 sg13g2_buf_16 clkbuf_8_183_0_clk (.X(clknet_8_183_0_clk),
    .A(clknet_7_91_0_clk));
 sg13g2_buf_16 clkbuf_8_184_0_clk (.X(clknet_8_184_0_clk),
    .A(clknet_7_92_0_clk));
 sg13g2_buf_16 clkbuf_8_185_0_clk (.X(clknet_8_185_0_clk),
    .A(clknet_7_92_0_clk));
 sg13g2_buf_16 clkbuf_8_186_0_clk (.X(clknet_8_186_0_clk),
    .A(clknet_7_93_0_clk));
 sg13g2_buf_16 clkbuf_8_187_0_clk (.X(clknet_8_187_0_clk),
    .A(clknet_7_93_0_clk));
 sg13g2_buf_16 clkbuf_8_188_0_clk (.X(clknet_8_188_0_clk),
    .A(clknet_7_94_0_clk));
 sg13g2_buf_16 clkbuf_8_189_0_clk (.X(clknet_8_189_0_clk),
    .A(clknet_7_94_0_clk));
 sg13g2_buf_16 clkbuf_8_190_0_clk (.X(clknet_8_190_0_clk),
    .A(clknet_7_95_0_clk));
 sg13g2_buf_16 clkbuf_8_191_0_clk (.X(clknet_8_191_0_clk),
    .A(clknet_7_95_0_clk));
 sg13g2_buf_16 clkbuf_8_192_0_clk (.X(clknet_8_192_0_clk),
    .A(clknet_7_96_0_clk));
 sg13g2_buf_16 clkbuf_8_193_0_clk (.X(clknet_8_193_0_clk),
    .A(clknet_7_96_0_clk));
 sg13g2_buf_16 clkbuf_8_194_0_clk (.X(clknet_8_194_0_clk),
    .A(clknet_7_97_0_clk));
 sg13g2_buf_16 clkbuf_8_195_0_clk (.X(clknet_8_195_0_clk),
    .A(clknet_7_97_0_clk));
 sg13g2_buf_16 clkbuf_8_196_0_clk (.X(clknet_8_196_0_clk),
    .A(clknet_7_98_0_clk));
 sg13g2_buf_16 clkbuf_8_197_0_clk (.X(clknet_8_197_0_clk),
    .A(clknet_7_98_0_clk));
 sg13g2_buf_16 clkbuf_8_198_0_clk (.X(clknet_8_198_0_clk),
    .A(clknet_7_99_0_clk));
 sg13g2_buf_16 clkbuf_8_199_0_clk (.X(clknet_8_199_0_clk),
    .A(clknet_7_99_0_clk));
 sg13g2_buf_16 clkbuf_8_200_0_clk (.X(clknet_8_200_0_clk),
    .A(clknet_7_100_0_clk));
 sg13g2_buf_16 clkbuf_8_201_0_clk (.X(clknet_8_201_0_clk),
    .A(clknet_7_100_0_clk));
 sg13g2_buf_16 clkbuf_8_202_0_clk (.X(clknet_8_202_0_clk),
    .A(clknet_7_101_0_clk));
 sg13g2_buf_16 clkbuf_8_203_0_clk (.X(clknet_8_203_0_clk),
    .A(clknet_7_101_0_clk));
 sg13g2_buf_16 clkbuf_8_204_0_clk (.X(clknet_8_204_0_clk),
    .A(clknet_7_102_0_clk));
 sg13g2_buf_16 clkbuf_8_205_0_clk (.X(clknet_8_205_0_clk),
    .A(clknet_7_102_0_clk));
 sg13g2_buf_16 clkbuf_8_206_0_clk (.X(clknet_8_206_0_clk),
    .A(clknet_7_103_0_clk));
 sg13g2_buf_16 clkbuf_8_207_0_clk (.X(clknet_8_207_0_clk),
    .A(clknet_7_103_0_clk));
 sg13g2_buf_16 clkbuf_8_208_0_clk (.X(clknet_8_208_0_clk),
    .A(clknet_7_104_0_clk));
 sg13g2_buf_16 clkbuf_8_209_0_clk (.X(clknet_8_209_0_clk),
    .A(clknet_7_104_0_clk));
 sg13g2_buf_16 clkbuf_8_210_0_clk (.X(clknet_8_210_0_clk),
    .A(clknet_7_105_0_clk));
 sg13g2_buf_16 clkbuf_8_211_0_clk (.X(clknet_8_211_0_clk),
    .A(clknet_7_105_0_clk));
 sg13g2_buf_16 clkbuf_8_212_0_clk (.X(clknet_8_212_0_clk),
    .A(clknet_7_106_0_clk));
 sg13g2_buf_16 clkbuf_8_213_0_clk (.X(clknet_8_213_0_clk),
    .A(clknet_7_106_0_clk));
 sg13g2_buf_16 clkbuf_8_214_0_clk (.X(clknet_8_214_0_clk),
    .A(clknet_7_107_0_clk));
 sg13g2_buf_16 clkbuf_8_215_0_clk (.X(clknet_8_215_0_clk),
    .A(clknet_7_107_0_clk));
 sg13g2_buf_16 clkbuf_8_216_0_clk (.X(clknet_8_216_0_clk),
    .A(clknet_7_108_0_clk));
 sg13g2_buf_16 clkbuf_8_217_0_clk (.X(clknet_8_217_0_clk),
    .A(clknet_7_108_0_clk));
 sg13g2_buf_16 clkbuf_8_218_0_clk (.X(clknet_8_218_0_clk),
    .A(clknet_7_109_0_clk));
 sg13g2_buf_16 clkbuf_8_219_0_clk (.X(clknet_8_219_0_clk),
    .A(clknet_7_109_0_clk));
 sg13g2_buf_16 clkbuf_8_220_0_clk (.X(clknet_8_220_0_clk),
    .A(clknet_7_110_0_clk));
 sg13g2_buf_16 clkbuf_8_221_0_clk (.X(clknet_8_221_0_clk),
    .A(clknet_7_110_0_clk));
 sg13g2_buf_16 clkbuf_8_222_0_clk (.X(clknet_8_222_0_clk),
    .A(clknet_7_111_0_clk));
 sg13g2_buf_16 clkbuf_8_223_0_clk (.X(clknet_8_223_0_clk),
    .A(clknet_7_111_0_clk));
 sg13g2_buf_16 clkbuf_8_224_0_clk (.X(clknet_8_224_0_clk),
    .A(clknet_7_112_0_clk));
 sg13g2_buf_16 clkbuf_8_225_0_clk (.X(clknet_8_225_0_clk),
    .A(clknet_7_112_0_clk));
 sg13g2_buf_16 clkbuf_8_226_0_clk (.X(clknet_8_226_0_clk),
    .A(clknet_7_113_0_clk));
 sg13g2_buf_16 clkbuf_8_227_0_clk (.X(clknet_8_227_0_clk),
    .A(clknet_7_113_0_clk));
 sg13g2_buf_16 clkbuf_8_228_0_clk (.X(clknet_8_228_0_clk),
    .A(clknet_7_114_0_clk));
 sg13g2_buf_16 clkbuf_8_229_0_clk (.X(clknet_8_229_0_clk),
    .A(clknet_7_114_0_clk));
 sg13g2_buf_16 clkbuf_8_230_0_clk (.X(clknet_8_230_0_clk),
    .A(clknet_7_115_0_clk));
 sg13g2_buf_16 clkbuf_8_231_0_clk (.X(clknet_8_231_0_clk),
    .A(clknet_7_115_0_clk));
 sg13g2_buf_16 clkbuf_8_232_0_clk (.X(clknet_8_232_0_clk),
    .A(clknet_7_116_0_clk));
 sg13g2_buf_16 clkbuf_8_233_0_clk (.X(clknet_8_233_0_clk),
    .A(clknet_7_116_0_clk));
 sg13g2_buf_16 clkbuf_8_234_0_clk (.X(clknet_8_234_0_clk),
    .A(clknet_7_117_0_clk));
 sg13g2_buf_16 clkbuf_8_235_0_clk (.X(clknet_8_235_0_clk),
    .A(clknet_7_117_0_clk));
 sg13g2_buf_16 clkbuf_8_236_0_clk (.X(clknet_8_236_0_clk),
    .A(clknet_7_118_0_clk));
 sg13g2_buf_16 clkbuf_8_237_0_clk (.X(clknet_8_237_0_clk),
    .A(clknet_7_118_0_clk));
 sg13g2_buf_16 clkbuf_8_238_0_clk (.X(clknet_8_238_0_clk),
    .A(clknet_7_119_0_clk));
 sg13g2_buf_16 clkbuf_8_239_0_clk (.X(clknet_8_239_0_clk),
    .A(clknet_7_119_0_clk));
 sg13g2_buf_16 clkbuf_8_240_0_clk (.X(clknet_8_240_0_clk),
    .A(clknet_7_120_0_clk));
 sg13g2_buf_16 clkbuf_8_241_0_clk (.X(clknet_8_241_0_clk),
    .A(clknet_7_120_0_clk));
 sg13g2_buf_16 clkbuf_8_242_0_clk (.X(clknet_8_242_0_clk),
    .A(clknet_7_121_0_clk));
 sg13g2_buf_16 clkbuf_8_243_0_clk (.X(clknet_8_243_0_clk),
    .A(clknet_7_121_0_clk));
 sg13g2_buf_16 clkbuf_8_244_0_clk (.X(clknet_8_244_0_clk),
    .A(clknet_7_122_0_clk));
 sg13g2_buf_16 clkbuf_8_245_0_clk (.X(clknet_8_245_0_clk),
    .A(clknet_7_122_0_clk));
 sg13g2_buf_16 clkbuf_8_246_0_clk (.X(clknet_8_246_0_clk),
    .A(clknet_7_123_0_clk));
 sg13g2_buf_16 clkbuf_8_247_0_clk (.X(clknet_8_247_0_clk),
    .A(clknet_7_123_0_clk));
 sg13g2_buf_16 clkbuf_8_248_0_clk (.X(clknet_8_248_0_clk),
    .A(clknet_7_124_0_clk));
 sg13g2_buf_16 clkbuf_8_249_0_clk (.X(clknet_8_249_0_clk),
    .A(clknet_7_124_0_clk));
 sg13g2_buf_16 clkbuf_8_250_0_clk (.X(clknet_8_250_0_clk),
    .A(clknet_7_125_0_clk));
 sg13g2_buf_16 clkbuf_8_251_0_clk (.X(clknet_8_251_0_clk),
    .A(clknet_7_125_0_clk));
 sg13g2_buf_16 clkbuf_8_252_0_clk (.X(clknet_8_252_0_clk),
    .A(clknet_7_126_0_clk));
 sg13g2_buf_16 clkbuf_8_253_0_clk (.X(clknet_8_253_0_clk),
    .A(clknet_7_126_0_clk));
 sg13g2_buf_16 clkbuf_8_254_0_clk (.X(clknet_8_254_0_clk),
    .A(clknet_7_127_0_clk));
 sg13g2_buf_16 clkbuf_8_255_0_clk (.X(clknet_8_255_0_clk),
    .A(clknet_7_127_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_8_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_8_3_0_clk));
 sg13g2_buf_16 clkload2 (.A(clknet_8_5_0_clk));
 sg13g2_buf_16 clkload3 (.A(clknet_8_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_8_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_8_11_0_clk));
 sg13g2_inv_8 clkload6 (.A(clknet_8_13_0_clk));
 sg13g2_buf_16 clkload7 (.A(clknet_8_15_0_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_8_16_0_clk));
 sg13g2_buf_16 clkload9 (.A(clknet_8_19_0_clk));
 sg13g2_buf_16 clkload10 (.A(clknet_8_21_0_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_8_22_0_clk));
 sg13g2_inv_8 clkload12 (.A(clknet_8_25_0_clk));
 sg13g2_inv_8 clkload13 (.A(clknet_8_27_0_clk));
 sg13g2_inv_8 clkload14 (.A(clknet_8_28_0_clk));
 sg13g2_buf_16 clkload15 (.A(clknet_8_31_0_clk));
 sg13g2_inv_8 clkload16 (.A(clknet_8_33_0_clk));
 sg13g2_buf_16 clkload17 (.A(clknet_8_35_0_clk));
 sg13g2_inv_8 clkload18 (.A(clknet_8_37_0_clk));
 sg13g2_buf_16 clkload19 (.A(clknet_8_39_0_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_8_41_0_clk));
 sg13g2_inv_16 clkload21 (.A(clknet_8_43_0_clk));
 sg13g2_buf_16 clkload22 (.A(clknet_8_45_0_clk));
 sg13g2_buf_16 clkload23 (.A(clknet_8_47_0_clk));
 sg13g2_buf_16 clkload24 (.A(clknet_8_49_0_clk));
 sg13g2_inv_8 clkload25 (.A(clknet_8_51_0_clk));
 sg13g2_buf_16 clkload26 (.A(clknet_8_53_0_clk));
 sg13g2_inv_8 clkload27 (.A(clknet_8_55_0_clk));
 sg13g2_inv_1 clkload28 (.A(clknet_8_57_0_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_8_59_0_clk));
 sg13g2_inv_16 clkload30 (.A(clknet_8_61_0_clk));
 sg13g2_inv_8 clkload31 (.A(clknet_8_63_0_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_8_65_0_clk));
 sg13g2_inv_8 clkload33 (.A(clknet_8_66_0_clk));
 sg13g2_inv_4 clkload34 (.A(clknet_8_68_0_clk));
 sg13g2_inv_8 clkload35 (.A(clknet_8_71_0_clk));
 sg13g2_inv_8 clkload36 (.A(clknet_8_73_0_clk));
 sg13g2_buf_16 clkload37 (.A(clknet_8_75_0_clk));
 sg13g2_inv_4 clkload38 (.A(clknet_8_76_0_clk));
 sg13g2_inv_4 clkload39 (.A(clknet_8_78_0_clk));
 sg13g2_inv_16 clkload40 (.A(clknet_8_81_0_clk));
 sg13g2_inv_8 clkload41 (.A(clknet_8_83_0_clk));
 sg13g2_inv_4 clkload42 (.A(clknet_8_84_0_clk));
 sg13g2_inv_4 clkload43 (.A(clknet_8_86_0_clk));
 sg13g2_buf_16 clkload44 (.A(clknet_8_89_0_clk));
 sg13g2_buf_16 clkload45 (.A(clknet_8_91_0_clk));
 sg13g2_inv_16 clkload46 (.A(clknet_8_93_0_clk));
 sg13g2_inv_16 clkload47 (.A(clknet_8_95_0_clk));
 sg13g2_buf_16 clkload48 (.A(clknet_8_97_0_clk));
 sg13g2_inv_1 clkload49 (.A(clknet_8_99_0_clk));
 sg13g2_inv_8 clkload50 (.A(clknet_8_101_0_clk));
 sg13g2_buf_16 clkload51 (.A(clknet_8_103_0_clk));
 sg13g2_buf_16 clkload52 (.A(clknet_8_105_0_clk));
 sg13g2_inv_8 clkload53 (.A(clknet_8_106_0_clk));
 sg13g2_inv_8 clkload54 (.A(clknet_8_109_0_clk));
 sg13g2_buf_16 clkload55 (.A(clknet_8_111_0_clk));
 sg13g2_inv_8 clkload56 (.A(clknet_8_112_0_clk));
 sg13g2_buf_16 clkload57 (.A(clknet_8_115_0_clk));
 sg13g2_inv_8 clkload58 (.A(clknet_8_117_0_clk));
 sg13g2_buf_16 clkload59 (.A(clknet_8_119_0_clk));
 sg13g2_inv_1 clkload60 (.A(clknet_8_121_0_clk));
 sg13g2_inv_8 clkload61 (.A(clknet_8_123_0_clk));
 sg13g2_inv_1 clkload62 (.A(clknet_8_125_0_clk));
 sg13g2_inv_8 clkload63 (.A(clknet_8_127_0_clk));
 sg13g2_inv_8 clkload64 (.A(clknet_8_129_0_clk));
 sg13g2_buf_16 clkload65 (.A(clknet_8_131_0_clk));
 sg13g2_inv_1 clkload66 (.A(clknet_8_133_0_clk));
 sg13g2_buf_16 clkload67 (.A(clknet_8_135_0_clk));
 sg13g2_inv_8 clkload68 (.A(clknet_8_137_0_clk));
 sg13g2_inv_1 clkload69 (.A(clknet_8_139_0_clk));
 sg13g2_buf_16 clkload70 (.A(clknet_8_141_0_clk));
 sg13g2_inv_8 clkload71 (.A(clknet_8_143_0_clk));
 sg13g2_buf_16 clkload72 (.A(clknet_8_145_0_clk));
 sg13g2_buf_16 clkload73 (.A(clknet_8_147_0_clk));
 sg13g2_inv_8 clkload74 (.A(clknet_8_149_0_clk));
 sg13g2_inv_16 clkload75 (.A(clknet_8_151_0_clk));
 sg13g2_inv_1 clkload76 (.A(clknet_8_153_0_clk));
 sg13g2_inv_4 clkload77 (.A(clknet_8_154_0_clk));
 sg13g2_inv_8 clkload78 (.A(clknet_8_157_0_clk));
 sg13g2_inv_1 clkload79 (.A(clknet_8_159_0_clk));
 sg13g2_buf_16 clkload80 (.A(clknet_8_161_0_clk));
 sg13g2_inv_16 clkload81 (.A(clknet_8_163_0_clk));
 sg13g2_inv_16 clkload82 (.A(clknet_8_165_0_clk));
 sg13g2_buf_16 clkload83 (.A(clknet_8_167_0_clk));
 sg13g2_inv_1 clkload84 (.A(clknet_8_169_0_clk));
 sg13g2_buf_16 clkload85 (.A(clknet_8_171_0_clk));
 sg13g2_buf_16 clkload86 (.A(clknet_8_173_0_clk));
 sg13g2_buf_16 clkload87 (.A(clknet_8_175_0_clk));
 sg13g2_inv_4 clkload88 (.A(clknet_8_176_0_clk));
 sg13g2_inv_1 clkload89 (.A(clknet_8_179_0_clk));
 sg13g2_buf_16 clkload90 (.A(clknet_8_181_0_clk));
 sg13g2_inv_16 clkload91 (.A(clknet_8_182_0_clk));
 sg13g2_buf_16 clkload92 (.A(clknet_8_185_0_clk));
 sg13g2_buf_16 clkload93 (.A(clknet_8_187_0_clk));
 sg13g2_buf_16 clkload94 (.A(clknet_8_189_0_clk));
 sg13g2_inv_8 clkload95 (.A(clknet_8_191_0_clk));
 sg13g2_inv_16 clkload96 (.A(clknet_8_193_0_clk));
 sg13g2_buf_16 clkload97 (.A(clknet_8_195_0_clk));
 sg13g2_inv_1 clkload98 (.A(clknet_8_197_0_clk));
 sg13g2_inv_4 clkload99 (.A(clknet_8_198_0_clk));
 sg13g2_buf_16 clkload100 (.A(clknet_8_201_0_clk));
 sg13g2_inv_1 clkload101 (.A(clknet_8_203_0_clk));
 sg13g2_inv_1 clkload102 (.A(clknet_8_205_0_clk));
 sg13g2_inv_4 clkload103 (.A(clknet_8_206_0_clk));
 sg13g2_buf_16 clkload104 (.A(clknet_8_209_0_clk));
 sg13g2_inv_1 clkload105 (.A(clknet_8_211_0_clk));
 sg13g2_inv_8 clkload106 (.A(clknet_8_213_0_clk));
 sg13g2_inv_1 clkload107 (.A(clknet_8_215_0_clk));
 sg13g2_inv_4 clkload108 (.A(clknet_8_216_0_clk));
 sg13g2_buf_16 clkload109 (.A(clknet_8_219_0_clk));
 sg13g2_buf_16 clkload110 (.A(clknet_8_221_0_clk));
 sg13g2_inv_1 clkload111 (.A(clknet_8_223_0_clk));
 sg13g2_inv_1 clkload112 (.A(clknet_8_225_0_clk));
 sg13g2_inv_8 clkload113 (.A(clknet_8_227_0_clk));
 sg13g2_inv_8 clkload114 (.A(clknet_8_229_0_clk));
 sg13g2_inv_1 clkload115 (.A(clknet_8_231_0_clk));
 sg13g2_inv_4 clkload116 (.A(clknet_8_232_0_clk));
 sg13g2_buf_16 clkload117 (.A(clknet_8_235_0_clk));
 sg13g2_buf_16 clkload118 (.A(clknet_8_237_0_clk));
 sg13g2_inv_1 clkload119 (.A(clknet_8_239_0_clk));
 sg13g2_inv_4 clkload120 (.A(clknet_8_240_0_clk));
 sg13g2_inv_16 clkload121 (.A(clknet_8_243_0_clk));
 sg13g2_buf_16 clkload122 (.A(clknet_8_245_0_clk));
 sg13g2_buf_16 clkload123 (.A(clknet_8_247_0_clk));
 sg13g2_inv_16 clkload124 (.A(clknet_8_249_0_clk));
 sg13g2_inv_1 clkload125 (.A(clknet_8_251_0_clk));
 sg13g2_buf_16 clkload126 (.A(clknet_8_253_0_clk));
 sg13g2_buf_16 clkload127 (.A(clknet_8_255_0_clk));
 sg13g2_inv_1 clkload128 (.A(clknet_leaf_44_clk));
 sg13g2_inv_1 clkload129 (.A(clknet_leaf_46_clk));
 sg13g2_inv_1 clkload130 (.A(clknet_leaf_59_clk));
 sg13g2_inv_1 clkload131 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload132 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload133 (.A(clknet_leaf_30_clk));
 sg13g2_inv_1 clkload134 (.A(clknet_leaf_29_clk));
 sg13g2_inv_1 clkload135 (.A(clknet_leaf_60_clk));
 sg13g2_inv_1 clkload136 (.A(clknet_leaf_49_clk));
 sg13g2_inv_1 clkload137 (.A(clknet_leaf_51_clk));
 sg13g2_inv_1 clkload138 (.A(clknet_leaf_56_clk));
 sg13g2_inv_1 clkload139 (.A(clknet_leaf_57_clk));
 sg13g2_inv_1 clkload140 (.A(clknet_leaf_62_clk));
 sg13g2_inv_1 clkload141 (.A(clknet_leaf_65_clk));
 sg13g2_inv_1 clkload142 (.A(clknet_leaf_90_clk));
 sg13g2_inv_1 clkload143 (.A(clknet_leaf_84_clk));
 sg13g2_inv_1 clkload144 (.A(clknet_leaf_85_clk));
 sg13g2_inv_1 clkload145 (.A(clknet_leaf_76_clk));
 sg13g2_inv_1 clkload146 (.A(clknet_leaf_114_clk));
 sg13g2_inv_1 clkload147 (.A(clknet_leaf_116_clk));
 sg13g2_inv_1 clkload148 (.A(clknet_leaf_104_clk));
 sg13g2_inv_1 clkload149 (.A(clknet_leaf_108_clk));
 sg13g2_inv_1 clkload150 (.A(clknet_leaf_1012_clk));
 sg13g2_inv_1 clkload151 (.A(clknet_leaf_212_clk));
 sg13g2_inv_2 clkload152 (.A(clknet_leaf_69_clk));
 sg13g2_inv_2 clkload153 (.A(clknet_leaf_71_clk));
 sg13g2_inv_1 clkload154 (.A(clknet_leaf_72_clk));
 sg13g2_inv_2 clkload155 (.A(clknet_leaf_73_clk));
 sg13g2_inv_1 clkload156 (.A(clknet_leaf_205_clk));
 sg13g2_inv_1 clkload157 (.A(clknet_leaf_117_clk));
 sg13g2_inv_1 clkload158 (.A(clknet_leaf_120_clk));
 sg13g2_inv_2 clkload159 (.A(clknet_leaf_121_clk));
 sg13g2_inv_2 clkload160 (.A(clknet_leaf_156_clk));
 sg13g2_inv_1 clkload161 (.A(clknet_leaf_122_clk));
 sg13g2_inv_1 clkload162 (.A(clknet_leaf_158_clk));
 sg13g2_inv_1 clkload163 (.A(clknet_leaf_113_clk));
 sg13g2_inv_1 clkload164 (.A(clknet_leaf_124_clk));
 sg13g2_inv_2 clkload165 (.A(clknet_leaf_152_clk));
 sg13g2_inv_1 clkload166 (.A(clknet_leaf_153_clk));
 sg13g2_inv_1 clkload167 (.A(clknet_leaf_155_clk));
 sg13g2_inv_2 clkload168 (.A(clknet_leaf_137_clk));
 sg13g2_inv_2 clkload169 (.A(clknet_leaf_151_clk));
 sg13g2_inv_1 clkload170 (.A(clknet_leaf_1098_clk));
 sg13g2_inv_1 clkload171 (.A(clknet_leaf_1099_clk));
 sg13g2_inv_1 clkload172 (.A(clknet_leaf_1146_clk));
 sg13g2_inv_1 clkload173 (.A(clknet_leaf_1147_clk));
 sg13g2_inv_1 clkload174 (.A(clknet_leaf_1145_clk));
 sg13g2_inv_1 clkload175 (.A(clknet_leaf_1093_clk));
 sg13g2_inv_1 clkload176 (.A(clknet_leaf_1096_clk));
 sg13g2_inv_1 clkload177 (.A(clknet_leaf_1105_clk));
 sg13g2_inv_1 clkload178 (.A(clknet_leaf_1109_clk));
 sg13g2_inv_1 clkload179 (.A(clknet_leaf_1116_clk));
 sg13g2_inv_1 clkload180 (.A(clknet_leaf_1124_clk));
 sg13g2_inv_1 clkload181 (.A(clknet_leaf_1089_clk));
 sg13g2_inv_1 clkload182 (.A(clknet_leaf_1090_clk));
 sg13g2_inv_1 clkload183 (.A(clknet_leaf_1091_clk));
 sg13g2_inv_1 clkload184 (.A(clknet_leaf_1088_clk));
 sg13g2_inv_1 clkload185 (.A(clknet_leaf_1110_clk));
 sg13g2_inv_1 clkload186 (.A(clknet_leaf_1112_clk));
 sg13g2_inv_1 clkload187 (.A(clknet_leaf_1035_clk));
 sg13g2_inv_1 clkload188 (.A(clknet_leaf_1032_clk));
 sg13g2_inv_1 clkload189 (.A(clknet_leaf_1033_clk));
 sg13g2_inv_1 clkload190 (.A(clknet_leaf_1114_clk));
 sg13g2_inv_1 clkload191 (.A(clknet_leaf_1031_clk));
 sg13g2_inv_1 clkload192 (.A(clknet_leaf_1034_clk));
 sg13g2_inv_1 clkload193 (.A(clknet_leaf_1040_clk));
 sg13g2_inv_1 clkload194 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload195 (.A(clknet_leaf_1136_clk));
 sg13g2_inv_1 clkload196 (.A(clknet_leaf_6_clk));
 sg13g2_inv_1 clkload197 (.A(clknet_leaf_1134_clk));
 sg13g2_inv_1 clkload198 (.A(clknet_leaf_1138_clk));
 sg13g2_inv_1 clkload199 (.A(clknet_leaf_1139_clk));
 sg13g2_inv_1 clkload200 (.A(clknet_leaf_39_clk));
 sg13g2_inv_1 clkload201 (.A(clknet_leaf_0_clk));
 sg13g2_inv_1 clkload202 (.A(clknet_leaf_36_clk));
 sg13g2_inv_1 clkload203 (.A(clknet_leaf_37_clk));
 sg13g2_inv_1 clkload204 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload205 (.A(clknet_leaf_1127_clk));
 sg13g2_inv_1 clkload206 (.A(clknet_leaf_1128_clk));
 sg13g2_inv_1 clkload207 (.A(clknet_leaf_1129_clk));
 sg13g2_inv_1 clkload208 (.A(clknet_leaf_1006_clk));
 sg13g2_inv_1 clkload209 (.A(clknet_leaf_1018_clk));
 sg13g2_inv_1 clkload210 (.A(clknet_leaf_1019_clk));
 sg13g2_inv_1 clkload211 (.A(clknet_leaf_105_clk));
 sg13g2_inv_1 clkload212 (.A(clknet_leaf_1015_clk));
 sg13g2_inv_1 clkload213 (.A(clknet_leaf_221_clk));
 sg13g2_inv_1 clkload214 (.A(clknet_leaf_232_clk));
 sg13g2_inv_1 clkload215 (.A(clknet_leaf_233_clk));
 sg13g2_inv_2 clkload216 (.A(clknet_leaf_231_clk));
 sg13g2_inv_2 clkload217 (.A(clknet_leaf_234_clk));
 sg13g2_inv_2 clkload218 (.A(clknet_leaf_240_clk));
 sg13g2_inv_1 clkload219 (.A(clknet_leaf_226_clk));
 sg13g2_inv_1 clkload220 (.A(clknet_leaf_229_clk));
 sg13g2_inv_1 clkload221 (.A(clknet_leaf_246_clk));
 sg13g2_buf_1 clkload222 (.A(clknet_leaf_236_clk));
 sg13g2_inv_1 clkload223 (.A(clknet_leaf_238_clk));
 sg13g2_inv_1 clkload224 (.A(clknet_leaf_242_clk));
 sg13g2_inv_1 clkload225 (.A(clknet_leaf_275_clk));
 sg13g2_inv_1 clkload226 (.A(clknet_leaf_182_clk));
 sg13g2_inv_1 clkload227 (.A(clknet_leaf_184_clk));
 sg13g2_inv_1 clkload228 (.A(clknet_leaf_186_clk));
 sg13g2_inv_1 clkload229 (.A(clknet_leaf_248_clk));
 sg13g2_inv_1 clkload230 (.A(clknet_leaf_166_clk));
 sg13g2_inv_1 clkload231 (.A(clknet_leaf_255_clk));
 sg13g2_inv_1 clkload232 (.A(clknet_leaf_271_clk));
 sg13g2_inv_1 clkload233 (.A(clknet_leaf_261_clk));
 sg13g2_inv_1 clkload234 (.A(clknet_leaf_262_clk));
 sg13g2_inv_1 clkload235 (.A(clknet_leaf_266_clk));
 sg13g2_inv_1 clkload236 (.A(clknet_leaf_316_clk));
 sg13g2_inv_1 clkload237 (.A(clknet_leaf_319_clk));
 sg13g2_inv_1 clkload238 (.A(clknet_leaf_172_clk));
 sg13g2_inv_1 clkload239 (.A(clknet_leaf_417_clk));
 sg13g2_inv_1 clkload240 (.A(clknet_leaf_419_clk));
 sg13g2_inv_1 clkload241 (.A(clknet_leaf_412_clk));
 sg13g2_inv_1 clkload242 (.A(clknet_leaf_414_clk));
 sg13g2_inv_1 clkload243 (.A(clknet_leaf_322_clk));
 sg13g2_inv_1 clkload244 (.A(clknet_leaf_293_clk));
 sg13g2_inv_1 clkload245 (.A(clknet_leaf_342_clk));
 sg13g2_inv_1 clkload246 (.A(clknet_leaf_343_clk));
 sg13g2_inv_1 clkload247 (.A(clknet_leaf_344_clk));
 sg13g2_inv_1 clkload248 (.A(clknet_leaf_147_clk));
 sg13g2_inv_1 clkload249 (.A(clknet_leaf_148_clk));
 sg13g2_inv_1 clkload250 (.A(clknet_leaf_162_clk));
 sg13g2_inv_1 clkload251 (.A(clknet_leaf_144_clk));
 sg13g2_inv_1 clkload252 (.A(clknet_leaf_444_clk));
 sg13g2_inv_1 clkload253 (.A(clknet_leaf_425_clk));
 sg13g2_inv_1 clkload254 (.A(clknet_leaf_442_clk));
 sg13g2_inv_1 clkload255 (.A(clknet_leaf_443_clk));
 sg13g2_inv_1 clkload256 (.A(clknet_leaf_395_clk));
 sg13g2_inv_1 clkload257 (.A(clknet_leaf_408_clk));
 sg13g2_inv_1 clkload258 (.A(clknet_leaf_409_clk));
 sg13g2_inv_1 clkload259 (.A(clknet_leaf_411_clk));
 sg13g2_inv_1 clkload260 (.A(clknet_leaf_428_clk));
 sg13g2_inv_1 clkload261 (.A(clknet_leaf_429_clk));
 sg13g2_inv_1 clkload262 (.A(clknet_leaf_389_clk));
 sg13g2_inv_1 clkload263 (.A(clknet_leaf_435_clk));
 sg13g2_inv_1 clkload264 (.A(clknet_leaf_434_clk));
 sg13g2_inv_1 clkload265 (.A(clknet_leaf_469_clk));
 sg13g2_inv_1 clkload266 (.A(clknet_leaf_473_clk));
 sg13g2_inv_1 clkload267 (.A(clknet_leaf_376_clk));
 sg13g2_inv_1 clkload268 (.A(clknet_leaf_397_clk));
 sg13g2_inv_1 clkload269 (.A(clknet_leaf_432_clk));
 sg13g2_inv_1 clkload270 (.A(clknet_leaf_386_clk));
 sg13g2_inv_1 clkload271 (.A(clknet_leaf_388_clk));
 sg13g2_inv_1 clkload272 (.A(clknet_leaf_474_clk));
 sg13g2_inv_1 clkload273 (.A(clknet_leaf_328_clk));
 sg13g2_inv_1 clkload274 (.A(clknet_leaf_329_clk));
 sg13g2_inv_1 clkload275 (.A(clknet_leaf_336_clk));
 sg13g2_inv_1 clkload276 (.A(clknet_leaf_400_clk));
 sg13g2_inv_1 clkload277 (.A(clknet_leaf_403_clk));
 sg13g2_inv_1 clkload278 (.A(clknet_leaf_404_clk));
 sg13g2_inv_1 clkload279 (.A(clknet_leaf_330_clk));
 sg13g2_inv_1 clkload280 (.A(clknet_leaf_333_clk));
 sg13g2_inv_1 clkload281 (.A(clknet_leaf_334_clk));
 sg13g2_inv_1 clkload282 (.A(clknet_leaf_335_clk));
 sg13g2_inv_1 clkload283 (.A(clknet_leaf_340_clk));
 sg13g2_inv_1 clkload284 (.A(clknet_leaf_341_clk));
 sg13g2_inv_1 clkload285 (.A(clknet_leaf_349_clk));
 sg13g2_inv_1 clkload286 (.A(clknet_leaf_352_clk));
 sg13g2_inv_1 clkload287 (.A(clknet_leaf_353_clk));
 sg13g2_inv_1 clkload288 (.A(clknet_leaf_368_clk));
 sg13g2_inv_1 clkload289 (.A(clknet_leaf_371_clk));
 sg13g2_inv_1 clkload290 (.A(clknet_leaf_543_clk));
 sg13g2_inv_1 clkload291 (.A(clknet_leaf_356_clk));
 sg13g2_inv_1 clkload292 (.A(clknet_leaf_370_clk));
 sg13g2_inv_1 clkload293 (.A(clknet_leaf_366_clk));
 sg13g2_inv_1 clkload294 (.A(clknet_leaf_369_clk));
 sg13g2_inv_1 clkload295 (.A(clknet_leaf_891_clk));
 sg13g2_inv_1 clkload296 (.A(clknet_leaf_892_clk));
 sg13g2_inv_1 clkload297 (.A(clknet_leaf_1070_clk));
 sg13g2_inv_1 clkload298 (.A(clknet_leaf_1071_clk));
 sg13g2_inv_1 clkload299 (.A(clknet_leaf_893_clk));
 sg13g2_inv_1 clkload300 (.A(clknet_leaf_894_clk));
 sg13g2_inv_1 clkload301 (.A(clknet_leaf_898_clk));
 sg13g2_inv_1 clkload302 (.A(clknet_leaf_1054_clk));
 sg13g2_inv_1 clkload303 (.A(clknet_leaf_1058_clk));
 sg13g2_inv_1 clkload304 (.A(clknet_leaf_1060_clk));
 sg13g2_inv_1 clkload305 (.A(clknet_leaf_896_clk));
 sg13g2_inv_1 clkload306 (.A(clknet_leaf_1067_clk));
 sg13g2_inv_1 clkload307 (.A(clknet_leaf_887_clk));
 sg13g2_inv_1 clkload308 (.A(clknet_leaf_869_clk));
 sg13g2_inv_1 clkload309 (.A(clknet_leaf_875_clk));
 sg13g2_inv_1 clkload310 (.A(clknet_leaf_877_clk));
 sg13g2_inv_1 clkload311 (.A(clknet_leaf_878_clk));
 sg13g2_inv_1 clkload312 (.A(clknet_leaf_904_clk));
 sg13g2_inv_1 clkload313 (.A(clknet_leaf_927_clk));
 sg13g2_inv_1 clkload314 (.A(clknet_leaf_929_clk));
 sg13g2_inv_1 clkload315 (.A(clknet_leaf_1044_clk));
 sg13g2_inv_1 clkload316 (.A(clknet_leaf_1045_clk));
 sg13g2_inv_1 clkload317 (.A(clknet_leaf_1056_clk));
 sg13g2_inv_1 clkload318 (.A(clknet_leaf_1049_clk));
 sg13g2_inv_1 clkload319 (.A(clknet_leaf_1051_clk));
 sg13g2_inv_1 clkload320 (.A(clknet_leaf_998_clk));
 sg13g2_inv_1 clkload321 (.A(clknet_leaf_1047_clk));
 sg13g2_inv_1 clkload322 (.A(clknet_leaf_131_clk));
 sg13g2_inv_1 clkload323 (.A(clknet_leaf_995_clk));
 sg13g2_inv_1 clkload324 (.A(clknet_leaf_997_clk));
 sg13g2_inv_1 clkload325 (.A(clknet_leaf_999_clk));
 sg13g2_inv_1 clkload326 (.A(clknet_leaf_917_clk));
 sg13g2_inv_1 clkload327 (.A(clknet_leaf_923_clk));
 sg13g2_inv_1 clkload328 (.A(clknet_leaf_926_clk));
 sg13g2_inv_1 clkload329 (.A(clknet_leaf_921_clk));
 sg13g2_inv_1 clkload330 (.A(clknet_leaf_948_clk));
 sg13g2_inv_1 clkload331 (.A(clknet_leaf_960_clk));
 sg13g2_inv_1 clkload332 (.A(clknet_leaf_968_clk));
 sg13g2_inv_1 clkload333 (.A(clknet_leaf_949_clk));
 sg13g2_inv_1 clkload334 (.A(clknet_leaf_865_clk));
 sg13g2_inv_1 clkload335 (.A(clknet_leaf_867_clk));
 sg13g2_inv_1 clkload336 (.A(clknet_leaf_874_clk));
 sg13g2_inv_1 clkload337 (.A(clknet_leaf_849_clk));
 sg13g2_inv_1 clkload338 (.A(clknet_leaf_850_clk));
 sg13g2_inv_1 clkload339 (.A(clknet_leaf_930_clk));
 sg13g2_inv_1 clkload340 (.A(clknet_leaf_932_clk));
 sg13g2_inv_1 clkload341 (.A(clknet_leaf_848_clk));
 sg13g2_inv_1 clkload342 (.A(clknet_leaf_931_clk));
 sg13g2_inv_1 clkload343 (.A(clknet_leaf_935_clk));
 sg13g2_inv_1 clkload344 (.A(clknet_leaf_946_clk));
 sg13g2_inv_1 clkload345 (.A(clknet_leaf_847_clk));
 sg13g2_inv_1 clkload346 (.A(clknet_leaf_858_clk));
 sg13g2_inv_1 clkload347 (.A(clknet_leaf_834_clk));
 sg13g2_inv_1 clkload348 (.A(clknet_leaf_780_clk));
 sg13g2_inv_1 clkload349 (.A(clknet_leaf_781_clk));
 sg13g2_inv_1 clkload350 (.A(clknet_leaf_774_clk));
 sg13g2_inv_1 clkload351 (.A(clknet_leaf_797_clk));
 sg13g2_inv_1 clkload352 (.A(clknet_leaf_790_clk));
 sg13g2_inv_1 clkload353 (.A(clknet_leaf_792_clk));
 sg13g2_inv_1 clkload354 (.A(clknet_leaf_793_clk));
 sg13g2_inv_1 clkload355 (.A(clknet_leaf_787_clk));
 sg13g2_inv_1 clkload356 (.A(clknet_leaf_789_clk));
 sg13g2_inv_1 clkload357 (.A(clknet_leaf_795_clk));
 sg13g2_inv_1 clkload358 (.A(clknet_leaf_775_clk));
 sg13g2_inv_1 clkload359 (.A(clknet_leaf_776_clk));
 sg13g2_inv_1 clkload360 (.A(clknet_leaf_765_clk));
 sg13g2_inv_1 clkload361 (.A(clknet_leaf_767_clk));
 sg13g2_inv_1 clkload362 (.A(clknet_leaf_772_clk));
 sg13g2_inv_1 clkload363 (.A(clknet_leaf_794_clk));
 sg13g2_inv_1 clkload364 (.A(clknet_leaf_807_clk));
 sg13g2_inv_1 clkload365 (.A(clknet_leaf_801_clk));
 sg13g2_inv_1 clkload366 (.A(clknet_leaf_750_clk));
 sg13g2_inv_1 clkload367 (.A(clknet_leaf_461_clk));
 sg13g2_inv_1 clkload368 (.A(clknet_leaf_648_clk));
 sg13g2_inv_1 clkload369 (.A(clknet_leaf_463_clk));
 sg13g2_inv_1 clkload370 (.A(clknet_leaf_481_clk));
 sg13g2_inv_1 clkload371 (.A(clknet_leaf_482_clk));
 sg13g2_inv_1 clkload372 (.A(clknet_leaf_487_clk));
 sg13g2_inv_1 clkload373 (.A(clknet_leaf_488_clk));
 sg13g2_inv_1 clkload374 (.A(clknet_leaf_502_clk));
 sg13g2_inv_1 clkload375 (.A(clknet_leaf_498_clk));
 sg13g2_inv_1 clkload376 (.A(clknet_leaf_501_clk));
 sg13g2_inv_1 clkload377 (.A(clknet_leaf_594_clk));
 sg13g2_inv_1 clkload378 (.A(clknet_leaf_497_clk));
 sg13g2_inv_1 clkload379 (.A(clknet_leaf_625_clk));
 sg13g2_inv_1 clkload380 (.A(clknet_leaf_493_clk));
 sg13g2_inv_1 clkload381 (.A(clknet_leaf_496_clk));
 sg13g2_inv_1 clkload382 (.A(clknet_leaf_590_clk));
 sg13g2_inv_1 clkload383 (.A(clknet_leaf_622_clk));
 sg13g2_inv_1 clkload384 (.A(clknet_leaf_475_clk));
 sg13g2_inv_1 clkload385 (.A(clknet_leaf_518_clk));
 sg13g2_inv_1 clkload386 (.A(clknet_leaf_513_clk));
 sg13g2_inv_1 clkload387 (.A(clknet_leaf_540_clk));
 sg13g2_inv_1 clkload388 (.A(clknet_leaf_541_clk));
 sg13g2_inv_2 clkload389 (.A(clknet_leaf_537_clk));
 sg13g2_inv_1 clkload390 (.A(clknet_leaf_553_clk));
 sg13g2_inv_1 clkload391 (.A(clknet_leaf_555_clk));
 sg13g2_inv_1 clkload392 (.A(clknet_leaf_507_clk));
 sg13g2_inv_1 clkload393 (.A(clknet_leaf_509_clk));
 sg13g2_inv_1 clkload394 (.A(clknet_leaf_585_clk));
 sg13g2_inv_1 clkload395 (.A(clknet_leaf_587_clk));
 sg13g2_inv_2 clkload396 (.A(clknet_leaf_579_clk));
 sg13g2_inv_1 clkload397 (.A(clknet_leaf_565_clk));
 sg13g2_inv_1 clkload398 (.A(clknet_leaf_571_clk));
 sg13g2_inv_1 clkload399 (.A(clknet_leaf_556_clk));
 sg13g2_inv_1 clkload400 (.A(clknet_leaf_567_clk));
 sg13g2_inv_1 clkload401 (.A(clknet_leaf_580_clk));
 sg13g2_inv_1 clkload402 (.A(clknet_leaf_581_clk));
 sg13g2_inv_1 clkload403 (.A(clknet_leaf_689_clk));
 sg13g2_inv_1 clkload404 (.A(clknet_leaf_690_clk));
 sg13g2_inv_1 clkload405 (.A(clknet_leaf_692_clk));
 sg13g2_inv_1 clkload406 (.A(clknet_leaf_693_clk));
 sg13g2_inv_1 clkload407 (.A(clknet_leaf_714_clk));
 sg13g2_inv_1 clkload408 (.A(clknet_leaf_605_clk));
 sg13g2_inv_1 clkload409 (.A(clknet_leaf_611_clk));
 sg13g2_inv_1 clkload410 (.A(clknet_leaf_705_clk));
 sg13g2_inv_1 clkload411 (.A(clknet_leaf_708_clk));
 sg13g2_inv_1 clkload412 (.A(clknet_leaf_711_clk));
 sg13g2_inv_1 clkload413 (.A(clknet_leaf_718_clk));
 sg13g2_inv_1 clkload414 (.A(clknet_leaf_731_clk));
 sg13g2_inv_1 clkload415 (.A(clknet_leaf_613_clk));
 sg13g2_inv_1 clkload416 (.A(clknet_leaf_726_clk));
 sg13g2_inv_1 clkload417 (.A(clknet_leaf_727_clk));
 sg13g2_inv_1 clkload418 (.A(clknet_leaf_728_clk));
 sg13g2_inv_1 clkload419 (.A(clknet_leaf_652_clk));
 sg13g2_inv_1 clkload420 (.A(clknet_leaf_654_clk));
 sg13g2_inv_1 clkload421 (.A(clknet_leaf_951_clk));
 sg13g2_inv_1 clkload422 (.A(clknet_leaf_953_clk));
 sg13g2_inv_1 clkload423 (.A(clknet_leaf_954_clk));
 sg13g2_inv_1 clkload424 (.A(clknet_leaf_676_clk));
 sg13g2_inv_1 clkload425 (.A(clknet_leaf_679_clk));
 sg13g2_inv_1 clkload426 (.A(clknet_leaf_943_clk));
 sg13g2_inv_1 clkload427 (.A(clknet_leaf_681_clk));
 sg13g2_inv_1 clkload428 (.A(clknet_leaf_699_clk));
 sg13g2_inv_1 clkload429 (.A(clknet_leaf_641_clk));
 sg13g2_inv_1 clkload430 (.A(clknet_leaf_700_clk));
 sg13g2_inv_1 clkload431 (.A(clknet_leaf_701_clk));
 sg13g2_inv_1 clkload432 (.A(clknet_leaf_706_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_4 FILLER_0_455 ();
 sg13g2_fill_2 FILLER_0_459 ();
 sg13g2_decap_8 FILLER_0_470 ();
 sg13g2_decap_8 FILLER_0_477 ();
 sg13g2_fill_2 FILLER_0_484 ();
 sg13g2_decap_8 FILLER_0_491 ();
 sg13g2_fill_1 FILLER_0_498 ();
 sg13g2_decap_8 FILLER_0_503 ();
 sg13g2_decap_8 FILLER_0_510 ();
 sg13g2_decap_8 FILLER_0_517 ();
 sg13g2_fill_2 FILLER_0_524 ();
 sg13g2_fill_1 FILLER_0_526 ();
 sg13g2_decap_8 FILLER_0_531 ();
 sg13g2_decap_4 FILLER_0_538 ();
 sg13g2_fill_1 FILLER_0_542 ();
 sg13g2_decap_4 FILLER_0_552 ();
 sg13g2_fill_1 FILLER_0_556 ();
 sg13g2_decap_8 FILLER_0_561 ();
 sg13g2_decap_8 FILLER_0_568 ();
 sg13g2_decap_8 FILLER_0_575 ();
 sg13g2_decap_8 FILLER_0_582 ();
 sg13g2_decap_8 FILLER_0_589 ();
 sg13g2_fill_2 FILLER_0_596 ();
 sg13g2_decap_8 FILLER_0_603 ();
 sg13g2_decap_8 FILLER_0_610 ();
 sg13g2_fill_2 FILLER_0_617 ();
 sg13g2_fill_2 FILLER_0_629 ();
 sg13g2_decap_8 FILLER_0_635 ();
 sg13g2_decap_8 FILLER_0_642 ();
 sg13g2_decap_8 FILLER_0_649 ();
 sg13g2_fill_2 FILLER_0_656 ();
 sg13g2_decap_8 FILLER_0_662 ();
 sg13g2_decap_4 FILLER_0_669 ();
 sg13g2_fill_2 FILLER_0_673 ();
 sg13g2_decap_4 FILLER_0_680 ();
 sg13g2_fill_2 FILLER_0_684 ();
 sg13g2_decap_8 FILLER_0_690 ();
 sg13g2_decap_4 FILLER_0_697 ();
 sg13g2_fill_2 FILLER_0_701 ();
 sg13g2_decap_4 FILLER_0_708 ();
 sg13g2_fill_1 FILLER_0_712 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_4 FILLER_0_724 ();
 sg13g2_fill_1 FILLER_0_728 ();
 sg13g2_decap_4 FILLER_0_734 ();
 sg13g2_fill_1 FILLER_0_738 ();
 sg13g2_decap_8 FILLER_0_743 ();
 sg13g2_decap_8 FILLER_0_750 ();
 sg13g2_decap_8 FILLER_0_757 ();
 sg13g2_decap_8 FILLER_0_764 ();
 sg13g2_decap_8 FILLER_0_771 ();
 sg13g2_decap_8 FILLER_0_778 ();
 sg13g2_fill_1 FILLER_0_785 ();
 sg13g2_decap_8 FILLER_0_790 ();
 sg13g2_decap_8 FILLER_0_797 ();
 sg13g2_decap_8 FILLER_0_804 ();
 sg13g2_decap_8 FILLER_0_811 ();
 sg13g2_decap_4 FILLER_0_818 ();
 sg13g2_fill_2 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_828 ();
 sg13g2_decap_8 FILLER_0_835 ();
 sg13g2_decap_8 FILLER_0_842 ();
 sg13g2_decap_8 FILLER_0_849 ();
 sg13g2_decap_8 FILLER_0_856 ();
 sg13g2_decap_8 FILLER_0_863 ();
 sg13g2_decap_8 FILLER_0_870 ();
 sg13g2_decap_8 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_0_884 ();
 sg13g2_decap_4 FILLER_0_891 ();
 sg13g2_fill_2 FILLER_0_895 ();
 sg13g2_decap_4 FILLER_0_902 ();
 sg13g2_fill_1 FILLER_0_906 ();
 sg13g2_decap_8 FILLER_0_911 ();
 sg13g2_fill_1 FILLER_0_918 ();
 sg13g2_decap_8 FILLER_0_932 ();
 sg13g2_decap_8 FILLER_0_939 ();
 sg13g2_decap_8 FILLER_0_946 ();
 sg13g2_decap_8 FILLER_0_953 ();
 sg13g2_decap_8 FILLER_0_960 ();
 sg13g2_decap_8 FILLER_0_967 ();
 sg13g2_decap_8 FILLER_0_974 ();
 sg13g2_decap_8 FILLER_0_981 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_8 FILLER_0_1025 ();
 sg13g2_decap_8 FILLER_0_1032 ();
 sg13g2_decap_4 FILLER_0_1039 ();
 sg13g2_fill_1 FILLER_0_1043 ();
 sg13g2_decap_8 FILLER_0_1052 ();
 sg13g2_decap_4 FILLER_0_1059 ();
 sg13g2_decap_8 FILLER_0_1072 ();
 sg13g2_decap_8 FILLER_0_1079 ();
 sg13g2_decap_4 FILLER_0_1091 ();
 sg13g2_decap_8 FILLER_0_1099 ();
 sg13g2_decap_8 FILLER_0_1106 ();
 sg13g2_decap_8 FILLER_0_1113 ();
 sg13g2_decap_8 FILLER_0_1120 ();
 sg13g2_decap_8 FILLER_0_1127 ();
 sg13g2_decap_8 FILLER_0_1134 ();
 sg13g2_decap_8 FILLER_0_1141 ();
 sg13g2_decap_8 FILLER_0_1148 ();
 sg13g2_decap_8 FILLER_0_1155 ();
 sg13g2_decap_8 FILLER_0_1162 ();
 sg13g2_decap_8 FILLER_0_1169 ();
 sg13g2_decap_8 FILLER_0_1176 ();
 sg13g2_decap_8 FILLER_0_1183 ();
 sg13g2_decap_8 FILLER_0_1190 ();
 sg13g2_decap_8 FILLER_0_1197 ();
 sg13g2_decap_8 FILLER_0_1204 ();
 sg13g2_decap_8 FILLER_0_1211 ();
 sg13g2_decap_8 FILLER_0_1218 ();
 sg13g2_decap_8 FILLER_0_1225 ();
 sg13g2_decap_8 FILLER_0_1232 ();
 sg13g2_decap_8 FILLER_0_1239 ();
 sg13g2_decap_8 FILLER_0_1246 ();
 sg13g2_decap_8 FILLER_0_1253 ();
 sg13g2_decap_8 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_decap_8 FILLER_0_1281 ();
 sg13g2_decap_8 FILLER_0_1288 ();
 sg13g2_decap_8 FILLER_0_1295 ();
 sg13g2_fill_1 FILLER_0_1302 ();
 sg13g2_decap_8 FILLER_0_1307 ();
 sg13g2_decap_8 FILLER_0_1314 ();
 sg13g2_decap_8 FILLER_0_1321 ();
 sg13g2_decap_8 FILLER_0_1328 ();
 sg13g2_decap_8 FILLER_0_1335 ();
 sg13g2_decap_8 FILLER_0_1342 ();
 sg13g2_decap_8 FILLER_0_1349 ();
 sg13g2_decap_8 FILLER_0_1356 ();
 sg13g2_decap_8 FILLER_0_1363 ();
 sg13g2_decap_8 FILLER_0_1370 ();
 sg13g2_fill_2 FILLER_0_1377 ();
 sg13g2_fill_1 FILLER_0_1379 ();
 sg13g2_decap_8 FILLER_0_1384 ();
 sg13g2_decap_8 FILLER_0_1391 ();
 sg13g2_decap_8 FILLER_0_1398 ();
 sg13g2_decap_8 FILLER_0_1405 ();
 sg13g2_decap_8 FILLER_0_1412 ();
 sg13g2_decap_8 FILLER_0_1419 ();
 sg13g2_decap_8 FILLER_0_1426 ();
 sg13g2_decap_8 FILLER_0_1433 ();
 sg13g2_decap_8 FILLER_0_1440 ();
 sg13g2_decap_8 FILLER_0_1447 ();
 sg13g2_decap_8 FILLER_0_1454 ();
 sg13g2_decap_8 FILLER_0_1461 ();
 sg13g2_decap_8 FILLER_0_1468 ();
 sg13g2_decap_8 FILLER_0_1475 ();
 sg13g2_decap_8 FILLER_0_1482 ();
 sg13g2_decap_8 FILLER_0_1489 ();
 sg13g2_decap_8 FILLER_0_1496 ();
 sg13g2_decap_8 FILLER_0_1503 ();
 sg13g2_decap_8 FILLER_0_1510 ();
 sg13g2_decap_8 FILLER_0_1517 ();
 sg13g2_decap_8 FILLER_0_1524 ();
 sg13g2_decap_8 FILLER_0_1531 ();
 sg13g2_decap_8 FILLER_0_1538 ();
 sg13g2_decap_8 FILLER_0_1545 ();
 sg13g2_decap_8 FILLER_0_1552 ();
 sg13g2_decap_8 FILLER_0_1559 ();
 sg13g2_decap_8 FILLER_0_1566 ();
 sg13g2_decap_8 FILLER_0_1573 ();
 sg13g2_decap_8 FILLER_0_1580 ();
 sg13g2_decap_8 FILLER_0_1587 ();
 sg13g2_fill_2 FILLER_0_1594 ();
 sg13g2_fill_1 FILLER_0_1596 ();
 sg13g2_decap_8 FILLER_0_1601 ();
 sg13g2_decap_8 FILLER_0_1608 ();
 sg13g2_decap_8 FILLER_0_1615 ();
 sg13g2_fill_2 FILLER_0_1622 ();
 sg13g2_fill_1 FILLER_0_1624 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_fill_1 FILLER_1_455 ();
 sg13g2_fill_2 FILLER_1_482 ();
 sg13g2_fill_2 FILLER_1_514 ();
 sg13g2_fill_1 FILLER_1_516 ();
 sg13g2_fill_2 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_4 FILLER_1_581 ();
 sg13g2_fill_1 FILLER_1_585 ();
 sg13g2_fill_2 FILLER_1_590 ();
 sg13g2_fill_1 FILLER_1_592 ();
 sg13g2_fill_2 FILLER_1_598 ();
 sg13g2_decap_8 FILLER_1_604 ();
 sg13g2_fill_2 FILLER_1_676 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_fill_2 FILLER_1_777 ();
 sg13g2_decap_4 FILLER_1_810 ();
 sg13g2_fill_2 FILLER_1_814 ();
 sg13g2_decap_8 FILLER_1_842 ();
 sg13g2_decap_8 FILLER_1_849 ();
 sg13g2_decap_8 FILLER_1_856 ();
 sg13g2_decap_8 FILLER_1_863 ();
 sg13g2_decap_8 FILLER_1_870 ();
 sg13g2_decap_8 FILLER_1_877 ();
 sg13g2_decap_4 FILLER_1_884 ();
 sg13g2_fill_1 FILLER_1_888 ();
 sg13g2_decap_4 FILLER_1_915 ();
 sg13g2_fill_1 FILLER_1_919 ();
 sg13g2_decap_8 FILLER_1_946 ();
 sg13g2_fill_2 FILLER_1_953 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_fill_2 FILLER_1_973 ();
 sg13g2_fill_1 FILLER_1_1018 ();
 sg13g2_decap_8 FILLER_1_1023 ();
 sg13g2_decap_8 FILLER_1_1113 ();
 sg13g2_decap_8 FILLER_1_1120 ();
 sg13g2_decap_8 FILLER_1_1127 ();
 sg13g2_decap_8 FILLER_1_1134 ();
 sg13g2_decap_8 FILLER_1_1141 ();
 sg13g2_decap_8 FILLER_1_1148 ();
 sg13g2_decap_8 FILLER_1_1155 ();
 sg13g2_decap_8 FILLER_1_1162 ();
 sg13g2_decap_8 FILLER_1_1169 ();
 sg13g2_decap_8 FILLER_1_1176 ();
 sg13g2_decap_8 FILLER_1_1183 ();
 sg13g2_decap_8 FILLER_1_1190 ();
 sg13g2_decap_8 FILLER_1_1197 ();
 sg13g2_decap_8 FILLER_1_1204 ();
 sg13g2_decap_8 FILLER_1_1211 ();
 sg13g2_decap_8 FILLER_1_1218 ();
 sg13g2_decap_8 FILLER_1_1225 ();
 sg13g2_decap_8 FILLER_1_1232 ();
 sg13g2_decap_8 FILLER_1_1239 ();
 sg13g2_decap_8 FILLER_1_1246 ();
 sg13g2_decap_8 FILLER_1_1253 ();
 sg13g2_decap_8 FILLER_1_1260 ();
 sg13g2_decap_8 FILLER_1_1267 ();
 sg13g2_decap_8 FILLER_1_1274 ();
 sg13g2_decap_8 FILLER_1_1281 ();
 sg13g2_decap_4 FILLER_1_1288 ();
 sg13g2_decap_8 FILLER_1_1323 ();
 sg13g2_decap_8 FILLER_1_1330 ();
 sg13g2_decap_8 FILLER_1_1337 ();
 sg13g2_decap_8 FILLER_1_1344 ();
 sg13g2_decap_4 FILLER_1_1351 ();
 sg13g2_fill_1 FILLER_1_1355 ();
 sg13g2_decap_4 FILLER_1_1365 ();
 sg13g2_fill_1 FILLER_1_1369 ();
 sg13g2_decap_8 FILLER_1_1401 ();
 sg13g2_decap_8 FILLER_1_1408 ();
 sg13g2_decap_8 FILLER_1_1415 ();
 sg13g2_decap_8 FILLER_1_1422 ();
 sg13g2_decap_8 FILLER_1_1429 ();
 sg13g2_decap_8 FILLER_1_1436 ();
 sg13g2_decap_8 FILLER_1_1443 ();
 sg13g2_decap_8 FILLER_1_1450 ();
 sg13g2_decap_8 FILLER_1_1457 ();
 sg13g2_decap_8 FILLER_1_1464 ();
 sg13g2_decap_8 FILLER_1_1471 ();
 sg13g2_decap_8 FILLER_1_1478 ();
 sg13g2_decap_8 FILLER_1_1485 ();
 sg13g2_decap_8 FILLER_1_1492 ();
 sg13g2_decap_8 FILLER_1_1499 ();
 sg13g2_decap_8 FILLER_1_1506 ();
 sg13g2_decap_8 FILLER_1_1513 ();
 sg13g2_decap_8 FILLER_1_1520 ();
 sg13g2_decap_8 FILLER_1_1527 ();
 sg13g2_decap_8 FILLER_1_1534 ();
 sg13g2_decap_8 FILLER_1_1541 ();
 sg13g2_decap_8 FILLER_1_1548 ();
 sg13g2_decap_8 FILLER_1_1555 ();
 sg13g2_decap_8 FILLER_1_1562 ();
 sg13g2_decap_8 FILLER_1_1569 ();
 sg13g2_decap_8 FILLER_1_1576 ();
 sg13g2_fill_2 FILLER_1_1583 ();
 sg13g2_decap_8 FILLER_1_1616 ();
 sg13g2_fill_2 FILLER_1_1623 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_4 FILLER_2_448 ();
 sg13g2_fill_2 FILLER_2_477 ();
 sg13g2_fill_1 FILLER_2_479 ();
 sg13g2_fill_1 FILLER_2_498 ();
 sg13g2_decap_8 FILLER_2_559 ();
 sg13g2_decap_8 FILLER_2_566 ();
 sg13g2_fill_1 FILLER_2_573 ();
 sg13g2_fill_2 FILLER_2_633 ();
 sg13g2_fill_1 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_653 ();
 sg13g2_decap_4 FILLER_2_660 ();
 sg13g2_fill_1 FILLER_2_664 ();
 sg13g2_decap_4 FILLER_2_698 ();
 sg13g2_fill_1 FILLER_2_702 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_4 FILLER_2_721 ();
 sg13g2_fill_2 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_fill_1 FILLER_2_751 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_fill_1 FILLER_2_777 ();
 sg13g2_fill_2 FILLER_2_782 ();
 sg13g2_fill_2 FILLER_2_813 ();
 sg13g2_decap_8 FILLER_2_824 ();
 sg13g2_fill_2 FILLER_2_831 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_4 FILLER_2_858 ();
 sg13g2_fill_2 FILLER_2_862 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_4 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_899 ();
 sg13g2_decap_4 FILLER_2_906 ();
 sg13g2_fill_2 FILLER_2_915 ();
 sg13g2_fill_1 FILLER_2_917 ();
 sg13g2_decap_4 FILLER_2_944 ();
 sg13g2_decap_4 FILLER_2_1008 ();
 sg13g2_decap_8 FILLER_2_1047 ();
 sg13g2_decap_8 FILLER_2_1054 ();
 sg13g2_decap_4 FILLER_2_1061 ();
 sg13g2_fill_1 FILLER_2_1065 ();
 sg13g2_decap_8 FILLER_2_1070 ();
 sg13g2_decap_8 FILLER_2_1077 ();
 sg13g2_decap_4 FILLER_2_1084 ();
 sg13g2_fill_2 FILLER_2_1088 ();
 sg13g2_decap_8 FILLER_2_1094 ();
 sg13g2_fill_2 FILLER_2_1101 ();
 sg13g2_decap_8 FILLER_2_1116 ();
 sg13g2_decap_8 FILLER_2_1123 ();
 sg13g2_decap_8 FILLER_2_1130 ();
 sg13g2_decap_8 FILLER_2_1137 ();
 sg13g2_decap_8 FILLER_2_1144 ();
 sg13g2_decap_8 FILLER_2_1151 ();
 sg13g2_decap_8 FILLER_2_1158 ();
 sg13g2_decap_8 FILLER_2_1165 ();
 sg13g2_decap_8 FILLER_2_1172 ();
 sg13g2_decap_8 FILLER_2_1179 ();
 sg13g2_decap_8 FILLER_2_1186 ();
 sg13g2_decap_8 FILLER_2_1193 ();
 sg13g2_decap_8 FILLER_2_1200 ();
 sg13g2_decap_8 FILLER_2_1207 ();
 sg13g2_decap_8 FILLER_2_1214 ();
 sg13g2_decap_8 FILLER_2_1221 ();
 sg13g2_decap_8 FILLER_2_1228 ();
 sg13g2_decap_8 FILLER_2_1235 ();
 sg13g2_decap_8 FILLER_2_1242 ();
 sg13g2_decap_8 FILLER_2_1249 ();
 sg13g2_decap_8 FILLER_2_1256 ();
 sg13g2_decap_8 FILLER_2_1263 ();
 sg13g2_decap_8 FILLER_2_1270 ();
 sg13g2_decap_8 FILLER_2_1277 ();
 sg13g2_decap_8 FILLER_2_1284 ();
 sg13g2_decap_8 FILLER_2_1291 ();
 sg13g2_decap_8 FILLER_2_1298 ();
 sg13g2_fill_2 FILLER_2_1305 ();
 sg13g2_decap_4 FILLER_2_1312 ();
 sg13g2_fill_1 FILLER_2_1316 ();
 sg13g2_decap_8 FILLER_2_1321 ();
 sg13g2_decap_8 FILLER_2_1328 ();
 sg13g2_decap_8 FILLER_2_1335 ();
 sg13g2_decap_8 FILLER_2_1342 ();
 sg13g2_decap_8 FILLER_2_1349 ();
 sg13g2_decap_8 FILLER_2_1356 ();
 sg13g2_decap_8 FILLER_2_1363 ();
 sg13g2_decap_8 FILLER_2_1370 ();
 sg13g2_decap_8 FILLER_2_1377 ();
 sg13g2_decap_8 FILLER_2_1384 ();
 sg13g2_decap_8 FILLER_2_1391 ();
 sg13g2_decap_8 FILLER_2_1398 ();
 sg13g2_decap_8 FILLER_2_1405 ();
 sg13g2_decap_8 FILLER_2_1412 ();
 sg13g2_decap_8 FILLER_2_1419 ();
 sg13g2_decap_8 FILLER_2_1426 ();
 sg13g2_decap_8 FILLER_2_1433 ();
 sg13g2_decap_8 FILLER_2_1440 ();
 sg13g2_decap_8 FILLER_2_1447 ();
 sg13g2_decap_8 FILLER_2_1454 ();
 sg13g2_decap_8 FILLER_2_1461 ();
 sg13g2_decap_8 FILLER_2_1468 ();
 sg13g2_decap_8 FILLER_2_1475 ();
 sg13g2_decap_8 FILLER_2_1482 ();
 sg13g2_decap_8 FILLER_2_1489 ();
 sg13g2_decap_8 FILLER_2_1496 ();
 sg13g2_decap_8 FILLER_2_1503 ();
 sg13g2_decap_8 FILLER_2_1510 ();
 sg13g2_decap_8 FILLER_2_1517 ();
 sg13g2_decap_8 FILLER_2_1524 ();
 sg13g2_decap_8 FILLER_2_1531 ();
 sg13g2_decap_8 FILLER_2_1538 ();
 sg13g2_decap_8 FILLER_2_1545 ();
 sg13g2_decap_8 FILLER_2_1552 ();
 sg13g2_decap_8 FILLER_2_1559 ();
 sg13g2_decap_8 FILLER_2_1566 ();
 sg13g2_decap_8 FILLER_2_1573 ();
 sg13g2_decap_8 FILLER_2_1585 ();
 sg13g2_decap_8 FILLER_2_1592 ();
 sg13g2_decap_8 FILLER_2_1599 ();
 sg13g2_decap_8 FILLER_2_1606 ();
 sg13g2_decap_8 FILLER_2_1613 ();
 sg13g2_decap_4 FILLER_2_1620 ();
 sg13g2_fill_1 FILLER_2_1624 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_4 FILLER_3_413 ();
 sg13g2_fill_2 FILLER_3_417 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_decap_4 FILLER_3_430 ();
 sg13g2_fill_1 FILLER_3_434 ();
 sg13g2_fill_1 FILLER_3_461 ();
 sg13g2_decap_8 FILLER_3_470 ();
 sg13g2_fill_1 FILLER_3_477 ();
 sg13g2_fill_2 FILLER_3_510 ();
 sg13g2_decap_8 FILLER_3_516 ();
 sg13g2_fill_2 FILLER_3_523 ();
 sg13g2_fill_2 FILLER_3_564 ();
 sg13g2_fill_1 FILLER_3_634 ();
 sg13g2_decap_8 FILLER_3_660 ();
 sg13g2_decap_8 FILLER_3_667 ();
 sg13g2_fill_2 FILLER_3_674 ();
 sg13g2_decap_4 FILLER_3_707 ();
 sg13g2_fill_1 FILLER_3_741 ();
 sg13g2_decap_4 FILLER_3_767 ();
 sg13g2_fill_1 FILLER_3_771 ();
 sg13g2_decap_8 FILLER_3_807 ();
 sg13g2_fill_2 FILLER_3_814 ();
 sg13g2_fill_1 FILLER_3_816 ();
 sg13g2_fill_1 FILLER_3_824 ();
 sg13g2_fill_1 FILLER_3_851 ();
 sg13g2_decap_4 FILLER_3_883 ();
 sg13g2_fill_2 FILLER_3_891 ();
 sg13g2_fill_1 FILLER_3_898 ();
 sg13g2_decap_8 FILLER_3_903 ();
 sg13g2_decap_4 FILLER_3_910 ();
 sg13g2_fill_1 FILLER_3_914 ();
 sg13g2_fill_2 FILLER_3_924 ();
 sg13g2_decap_8 FILLER_3_951 ();
 sg13g2_decap_8 FILLER_3_967 ();
 sg13g2_fill_1 FILLER_3_974 ();
 sg13g2_decap_4 FILLER_3_1001 ();
 sg13g2_fill_2 FILLER_3_1005 ();
 sg13g2_fill_1 FILLER_3_1012 ();
 sg13g2_decap_8 FILLER_3_1017 ();
 sg13g2_decap_4 FILLER_3_1024 ();
 sg13g2_fill_2 FILLER_3_1028 ();
 sg13g2_fill_2 FILLER_3_1055 ();
 sg13g2_fill_1 FILLER_3_1057 ();
 sg13g2_decap_8 FILLER_3_1090 ();
 sg13g2_decap_8 FILLER_3_1097 ();
 sg13g2_fill_1 FILLER_3_1104 ();
 sg13g2_fill_1 FILLER_3_1131 ();
 sg13g2_decap_8 FILLER_3_1136 ();
 sg13g2_decap_8 FILLER_3_1143 ();
 sg13g2_decap_8 FILLER_3_1150 ();
 sg13g2_decap_8 FILLER_3_1157 ();
 sg13g2_decap_8 FILLER_3_1164 ();
 sg13g2_decap_8 FILLER_3_1171 ();
 sg13g2_decap_8 FILLER_3_1178 ();
 sg13g2_decap_8 FILLER_3_1185 ();
 sg13g2_decap_8 FILLER_3_1192 ();
 sg13g2_decap_8 FILLER_3_1199 ();
 sg13g2_decap_8 FILLER_3_1206 ();
 sg13g2_decap_8 FILLER_3_1213 ();
 sg13g2_decap_8 FILLER_3_1220 ();
 sg13g2_decap_8 FILLER_3_1227 ();
 sg13g2_decap_8 FILLER_3_1234 ();
 sg13g2_decap_8 FILLER_3_1241 ();
 sg13g2_decap_8 FILLER_3_1248 ();
 sg13g2_decap_8 FILLER_3_1255 ();
 sg13g2_decap_8 FILLER_3_1262 ();
 sg13g2_decap_8 FILLER_3_1269 ();
 sg13g2_decap_8 FILLER_3_1276 ();
 sg13g2_decap_8 FILLER_3_1283 ();
 sg13g2_decap_8 FILLER_3_1290 ();
 sg13g2_decap_8 FILLER_3_1297 ();
 sg13g2_decap_4 FILLER_3_1304 ();
 sg13g2_decap_8 FILLER_3_1333 ();
 sg13g2_decap_8 FILLER_3_1340 ();
 sg13g2_decap_8 FILLER_3_1347 ();
 sg13g2_decap_8 FILLER_3_1354 ();
 sg13g2_decap_8 FILLER_3_1361 ();
 sg13g2_decap_8 FILLER_3_1368 ();
 sg13g2_decap_8 FILLER_3_1375 ();
 sg13g2_decap_8 FILLER_3_1382 ();
 sg13g2_decap_8 FILLER_3_1389 ();
 sg13g2_decap_8 FILLER_3_1396 ();
 sg13g2_decap_8 FILLER_3_1403 ();
 sg13g2_decap_8 FILLER_3_1410 ();
 sg13g2_decap_8 FILLER_3_1417 ();
 sg13g2_decap_8 FILLER_3_1424 ();
 sg13g2_decap_8 FILLER_3_1431 ();
 sg13g2_decap_8 FILLER_3_1438 ();
 sg13g2_decap_8 FILLER_3_1445 ();
 sg13g2_decap_8 FILLER_3_1452 ();
 sg13g2_decap_8 FILLER_3_1459 ();
 sg13g2_decap_8 FILLER_3_1466 ();
 sg13g2_decap_8 FILLER_3_1473 ();
 sg13g2_decap_8 FILLER_3_1480 ();
 sg13g2_decap_8 FILLER_3_1487 ();
 sg13g2_decap_8 FILLER_3_1494 ();
 sg13g2_decap_8 FILLER_3_1501 ();
 sg13g2_decap_8 FILLER_3_1508 ();
 sg13g2_decap_8 FILLER_3_1515 ();
 sg13g2_decap_8 FILLER_3_1522 ();
 sg13g2_decap_8 FILLER_3_1529 ();
 sg13g2_decap_8 FILLER_3_1536 ();
 sg13g2_decap_8 FILLER_3_1543 ();
 sg13g2_decap_8 FILLER_3_1550 ();
 sg13g2_decap_8 FILLER_3_1557 ();
 sg13g2_decap_8 FILLER_3_1564 ();
 sg13g2_decap_8 FILLER_3_1571 ();
 sg13g2_decap_8 FILLER_3_1578 ();
 sg13g2_decap_8 FILLER_3_1585 ();
 sg13g2_decap_8 FILLER_3_1592 ();
 sg13g2_decap_8 FILLER_3_1599 ();
 sg13g2_decap_8 FILLER_3_1606 ();
 sg13g2_decap_8 FILLER_3_1613 ();
 sg13g2_decap_4 FILLER_3_1620 ();
 sg13g2_fill_1 FILLER_3_1624 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_fill_1 FILLER_4_385 ();
 sg13g2_decap_4 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_410 ();
 sg13g2_decap_4 FILLER_4_438 ();
 sg13g2_fill_2 FILLER_4_442 ();
 sg13g2_fill_2 FILLER_4_448 ();
 sg13g2_fill_1 FILLER_4_450 ();
 sg13g2_decap_8 FILLER_4_524 ();
 sg13g2_decap_4 FILLER_4_531 ();
 sg13g2_fill_2 FILLER_4_586 ();
 sg13g2_fill_2 FILLER_4_635 ();
 sg13g2_fill_2 FILLER_4_684 ();
 sg13g2_decap_8 FILLER_4_771 ();
 sg13g2_decap_8 FILLER_4_778 ();
 sg13g2_fill_2 FILLER_4_785 ();
 sg13g2_fill_1 FILLER_4_787 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_fill_2 FILLER_4_805 ();
 sg13g2_fill_1 FILLER_4_807 ();
 sg13g2_fill_2 FILLER_4_843 ();
 sg13g2_fill_2 FILLER_4_879 ();
 sg13g2_decap_4 FILLER_4_911 ();
 sg13g2_fill_2 FILLER_4_920 ();
 sg13g2_fill_1 FILLER_4_922 ();
 sg13g2_fill_1 FILLER_4_932 ();
 sg13g2_decap_8 FILLER_4_937 ();
 sg13g2_decap_8 FILLER_4_944 ();
 sg13g2_fill_1 FILLER_4_951 ();
 sg13g2_decap_8 FILLER_4_978 ();
 sg13g2_decap_8 FILLER_4_985 ();
 sg13g2_decap_8 FILLER_4_992 ();
 sg13g2_decap_4 FILLER_4_999 ();
 sg13g2_fill_2 FILLER_4_1063 ();
 sg13g2_decap_8 FILLER_4_1100 ();
 sg13g2_decap_4 FILLER_4_1107 ();
 sg13g2_fill_1 FILLER_4_1111 ();
 sg13g2_decap_8 FILLER_4_1150 ();
 sg13g2_decap_8 FILLER_4_1157 ();
 sg13g2_decap_8 FILLER_4_1164 ();
 sg13g2_decap_8 FILLER_4_1171 ();
 sg13g2_decap_8 FILLER_4_1178 ();
 sg13g2_decap_8 FILLER_4_1185 ();
 sg13g2_decap_8 FILLER_4_1192 ();
 sg13g2_decap_8 FILLER_4_1199 ();
 sg13g2_decap_8 FILLER_4_1206 ();
 sg13g2_decap_8 FILLER_4_1213 ();
 sg13g2_decap_8 FILLER_4_1220 ();
 sg13g2_decap_8 FILLER_4_1227 ();
 sg13g2_decap_8 FILLER_4_1234 ();
 sg13g2_decap_8 FILLER_4_1241 ();
 sg13g2_decap_8 FILLER_4_1248 ();
 sg13g2_decap_8 FILLER_4_1255 ();
 sg13g2_decap_8 FILLER_4_1262 ();
 sg13g2_decap_8 FILLER_4_1269 ();
 sg13g2_decap_8 FILLER_4_1276 ();
 sg13g2_decap_8 FILLER_4_1283 ();
 sg13g2_decap_8 FILLER_4_1290 ();
 sg13g2_decap_8 FILLER_4_1297 ();
 sg13g2_decap_4 FILLER_4_1304 ();
 sg13g2_fill_1 FILLER_4_1308 ();
 sg13g2_decap_8 FILLER_4_1335 ();
 sg13g2_decap_8 FILLER_4_1342 ();
 sg13g2_decap_8 FILLER_4_1349 ();
 sg13g2_decap_8 FILLER_4_1356 ();
 sg13g2_decap_8 FILLER_4_1363 ();
 sg13g2_decap_8 FILLER_4_1370 ();
 sg13g2_decap_8 FILLER_4_1377 ();
 sg13g2_decap_8 FILLER_4_1384 ();
 sg13g2_decap_8 FILLER_4_1391 ();
 sg13g2_decap_8 FILLER_4_1398 ();
 sg13g2_decap_8 FILLER_4_1405 ();
 sg13g2_decap_8 FILLER_4_1412 ();
 sg13g2_decap_8 FILLER_4_1419 ();
 sg13g2_decap_8 FILLER_4_1426 ();
 sg13g2_decap_8 FILLER_4_1433 ();
 sg13g2_decap_8 FILLER_4_1440 ();
 sg13g2_decap_8 FILLER_4_1447 ();
 sg13g2_decap_8 FILLER_4_1454 ();
 sg13g2_decap_8 FILLER_4_1461 ();
 sg13g2_decap_8 FILLER_4_1468 ();
 sg13g2_decap_8 FILLER_4_1475 ();
 sg13g2_decap_8 FILLER_4_1482 ();
 sg13g2_decap_8 FILLER_4_1489 ();
 sg13g2_decap_8 FILLER_4_1496 ();
 sg13g2_decap_8 FILLER_4_1503 ();
 sg13g2_decap_8 FILLER_4_1510 ();
 sg13g2_decap_8 FILLER_4_1517 ();
 sg13g2_decap_8 FILLER_4_1524 ();
 sg13g2_decap_8 FILLER_4_1531 ();
 sg13g2_decap_8 FILLER_4_1538 ();
 sg13g2_decap_8 FILLER_4_1545 ();
 sg13g2_decap_8 FILLER_4_1552 ();
 sg13g2_decap_8 FILLER_4_1559 ();
 sg13g2_decap_8 FILLER_4_1566 ();
 sg13g2_decap_8 FILLER_4_1573 ();
 sg13g2_decap_8 FILLER_4_1580 ();
 sg13g2_decap_8 FILLER_4_1587 ();
 sg13g2_decap_8 FILLER_4_1594 ();
 sg13g2_decap_8 FILLER_4_1601 ();
 sg13g2_decap_8 FILLER_4_1608 ();
 sg13g2_decap_8 FILLER_4_1615 ();
 sg13g2_fill_2 FILLER_4_1622 ();
 sg13g2_fill_1 FILLER_4_1624 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_fill_1 FILLER_5_385 ();
 sg13g2_decap_4 FILLER_5_412 ();
 sg13g2_fill_2 FILLER_5_416 ();
 sg13g2_fill_1 FILLER_5_426 ();
 sg13g2_fill_1 FILLER_5_435 ();
 sg13g2_fill_1 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_446 ();
 sg13g2_fill_2 FILLER_5_453 ();
 sg13g2_fill_1 FILLER_5_455 ();
 sg13g2_decap_4 FILLER_5_461 ();
 sg13g2_fill_1 FILLER_5_465 ();
 sg13g2_decap_8 FILLER_5_470 ();
 sg13g2_decap_8 FILLER_5_477 ();
 sg13g2_decap_8 FILLER_5_484 ();
 sg13g2_decap_8 FILLER_5_491 ();
 sg13g2_fill_2 FILLER_5_498 ();
 sg13g2_decap_4 FILLER_5_521 ();
 sg13g2_fill_2 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_fill_2 FILLER_5_546 ();
 sg13g2_fill_1 FILLER_5_574 ();
 sg13g2_fill_2 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_632 ();
 sg13g2_decap_8 FILLER_5_639 ();
 sg13g2_decap_8 FILLER_5_646 ();
 sg13g2_decap_8 FILLER_5_653 ();
 sg13g2_fill_2 FILLER_5_660 ();
 sg13g2_fill_1 FILLER_5_662 ();
 sg13g2_fill_2 FILLER_5_684 ();
 sg13g2_fill_2 FILLER_5_717 ();
 sg13g2_decap_8 FILLER_5_723 ();
 sg13g2_decap_4 FILLER_5_730 ();
 sg13g2_fill_2 FILLER_5_734 ();
 sg13g2_decap_4 FILLER_5_757 ();
 sg13g2_fill_1 FILLER_5_761 ();
 sg13g2_fill_1 FILLER_5_771 ();
 sg13g2_decap_8 FILLER_5_776 ();
 sg13g2_fill_2 FILLER_5_783 ();
 sg13g2_fill_1 FILLER_5_785 ();
 sg13g2_fill_2 FILLER_5_807 ();
 sg13g2_fill_1 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_fill_2 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_875 ();
 sg13g2_decap_8 FILLER_5_882 ();
 sg13g2_decap_4 FILLER_5_919 ();
 sg13g2_fill_2 FILLER_5_923 ();
 sg13g2_decap_8 FILLER_5_964 ();
 sg13g2_decap_8 FILLER_5_971 ();
 sg13g2_decap_8 FILLER_5_978 ();
 sg13g2_decap_4 FILLER_5_985 ();
 sg13g2_decap_4 FILLER_5_994 ();
 sg13g2_decap_4 FILLER_5_1031 ();
 sg13g2_decap_8 FILLER_5_1039 ();
 sg13g2_fill_1 FILLER_5_1046 ();
 sg13g2_decap_4 FILLER_5_1078 ();
 sg13g2_fill_2 FILLER_5_1117 ();
 sg13g2_decap_8 FILLER_5_1144 ();
 sg13g2_decap_8 FILLER_5_1151 ();
 sg13g2_decap_8 FILLER_5_1158 ();
 sg13g2_decap_8 FILLER_5_1165 ();
 sg13g2_decap_8 FILLER_5_1172 ();
 sg13g2_decap_8 FILLER_5_1179 ();
 sg13g2_decap_8 FILLER_5_1186 ();
 sg13g2_decap_8 FILLER_5_1193 ();
 sg13g2_decap_8 FILLER_5_1200 ();
 sg13g2_decap_8 FILLER_5_1207 ();
 sg13g2_decap_8 FILLER_5_1214 ();
 sg13g2_decap_8 FILLER_5_1221 ();
 sg13g2_decap_8 FILLER_5_1228 ();
 sg13g2_decap_8 FILLER_5_1235 ();
 sg13g2_decap_8 FILLER_5_1242 ();
 sg13g2_decap_8 FILLER_5_1249 ();
 sg13g2_decap_8 FILLER_5_1256 ();
 sg13g2_decap_8 FILLER_5_1263 ();
 sg13g2_decap_8 FILLER_5_1270 ();
 sg13g2_decap_8 FILLER_5_1277 ();
 sg13g2_decap_8 FILLER_5_1284 ();
 sg13g2_decap_8 FILLER_5_1291 ();
 sg13g2_decap_8 FILLER_5_1298 ();
 sg13g2_decap_8 FILLER_5_1305 ();
 sg13g2_decap_8 FILLER_5_1312 ();
 sg13g2_decap_8 FILLER_5_1319 ();
 sg13g2_decap_8 FILLER_5_1326 ();
 sg13g2_decap_8 FILLER_5_1333 ();
 sg13g2_decap_8 FILLER_5_1340 ();
 sg13g2_decap_8 FILLER_5_1347 ();
 sg13g2_decap_8 FILLER_5_1354 ();
 sg13g2_decap_8 FILLER_5_1361 ();
 sg13g2_decap_8 FILLER_5_1368 ();
 sg13g2_decap_8 FILLER_5_1375 ();
 sg13g2_decap_8 FILLER_5_1382 ();
 sg13g2_decap_8 FILLER_5_1389 ();
 sg13g2_decap_8 FILLER_5_1396 ();
 sg13g2_decap_8 FILLER_5_1403 ();
 sg13g2_decap_8 FILLER_5_1410 ();
 sg13g2_decap_8 FILLER_5_1417 ();
 sg13g2_decap_8 FILLER_5_1424 ();
 sg13g2_decap_8 FILLER_5_1431 ();
 sg13g2_decap_8 FILLER_5_1438 ();
 sg13g2_decap_8 FILLER_5_1445 ();
 sg13g2_decap_8 FILLER_5_1452 ();
 sg13g2_decap_8 FILLER_5_1459 ();
 sg13g2_decap_8 FILLER_5_1466 ();
 sg13g2_decap_8 FILLER_5_1473 ();
 sg13g2_decap_8 FILLER_5_1480 ();
 sg13g2_decap_8 FILLER_5_1487 ();
 sg13g2_decap_8 FILLER_5_1494 ();
 sg13g2_decap_8 FILLER_5_1501 ();
 sg13g2_decap_8 FILLER_5_1508 ();
 sg13g2_decap_8 FILLER_5_1515 ();
 sg13g2_decap_8 FILLER_5_1522 ();
 sg13g2_decap_8 FILLER_5_1529 ();
 sg13g2_decap_8 FILLER_5_1536 ();
 sg13g2_decap_8 FILLER_5_1543 ();
 sg13g2_decap_8 FILLER_5_1550 ();
 sg13g2_decap_8 FILLER_5_1557 ();
 sg13g2_decap_8 FILLER_5_1564 ();
 sg13g2_decap_8 FILLER_5_1571 ();
 sg13g2_decap_8 FILLER_5_1578 ();
 sg13g2_decap_8 FILLER_5_1585 ();
 sg13g2_decap_8 FILLER_5_1592 ();
 sg13g2_decap_8 FILLER_5_1599 ();
 sg13g2_decap_8 FILLER_5_1606 ();
 sg13g2_decap_8 FILLER_5_1613 ();
 sg13g2_decap_4 FILLER_5_1620 ();
 sg13g2_fill_1 FILLER_5_1624 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_4 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_fill_2 FILLER_6_386 ();
 sg13g2_fill_1 FILLER_6_413 ();
 sg13g2_fill_2 FILLER_6_419 ();
 sg13g2_decap_8 FILLER_6_446 ();
 sg13g2_decap_8 FILLER_6_453 ();
 sg13g2_decap_8 FILLER_6_460 ();
 sg13g2_fill_2 FILLER_6_467 ();
 sg13g2_fill_1 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_491 ();
 sg13g2_decap_8 FILLER_6_498 ();
 sg13g2_decap_8 FILLER_6_505 ();
 sg13g2_fill_1 FILLER_6_512 ();
 sg13g2_decap_8 FILLER_6_555 ();
 sg13g2_decap_8 FILLER_6_562 ();
 sg13g2_fill_1 FILLER_6_569 ();
 sg13g2_decap_4 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_652 ();
 sg13g2_decap_8 FILLER_6_659 ();
 sg13g2_decap_8 FILLER_6_666 ();
 sg13g2_decap_8 FILLER_6_673 ();
 sg13g2_decap_8 FILLER_6_680 ();
 sg13g2_decap_8 FILLER_6_691 ();
 sg13g2_decap_8 FILLER_6_698 ();
 sg13g2_decap_8 FILLER_6_705 ();
 sg13g2_decap_4 FILLER_6_759 ();
 sg13g2_fill_2 FILLER_6_825 ();
 sg13g2_fill_1 FILLER_6_827 ();
 sg13g2_decap_8 FILLER_6_832 ();
 sg13g2_decap_8 FILLER_6_839 ();
 sg13g2_decap_8 FILLER_6_846 ();
 sg13g2_decap_4 FILLER_6_858 ();
 sg13g2_fill_1 FILLER_6_862 ();
 sg13g2_decap_8 FILLER_6_867 ();
 sg13g2_decap_8 FILLER_6_874 ();
 sg13g2_decap_8 FILLER_6_885 ();
 sg13g2_decap_8 FILLER_6_948 ();
 sg13g2_decap_4 FILLER_6_955 ();
 sg13g2_fill_2 FILLER_6_959 ();
 sg13g2_decap_8 FILLER_6_966 ();
 sg13g2_fill_2 FILLER_6_977 ();
 sg13g2_fill_1 FILLER_6_979 ();
 sg13g2_fill_1 FILLER_6_1010 ();
 sg13g2_decap_8 FILLER_6_1032 ();
 sg13g2_fill_2 FILLER_6_1039 ();
 sg13g2_fill_1 FILLER_6_1041 ();
 sg13g2_decap_8 FILLER_6_1046 ();
 sg13g2_decap_8 FILLER_6_1053 ();
 sg13g2_decap_8 FILLER_6_1081 ();
 sg13g2_fill_1 FILLER_6_1088 ();
 sg13g2_decap_8 FILLER_6_1135 ();
 sg13g2_decap_8 FILLER_6_1142 ();
 sg13g2_decap_8 FILLER_6_1149 ();
 sg13g2_decap_8 FILLER_6_1156 ();
 sg13g2_decap_8 FILLER_6_1163 ();
 sg13g2_decap_8 FILLER_6_1170 ();
 sg13g2_decap_8 FILLER_6_1177 ();
 sg13g2_decap_8 FILLER_6_1184 ();
 sg13g2_decap_8 FILLER_6_1191 ();
 sg13g2_decap_8 FILLER_6_1198 ();
 sg13g2_decap_8 FILLER_6_1205 ();
 sg13g2_decap_8 FILLER_6_1212 ();
 sg13g2_decap_8 FILLER_6_1219 ();
 sg13g2_decap_8 FILLER_6_1226 ();
 sg13g2_decap_8 FILLER_6_1233 ();
 sg13g2_decap_8 FILLER_6_1240 ();
 sg13g2_decap_8 FILLER_6_1247 ();
 sg13g2_decap_8 FILLER_6_1254 ();
 sg13g2_decap_8 FILLER_6_1261 ();
 sg13g2_decap_8 FILLER_6_1268 ();
 sg13g2_decap_8 FILLER_6_1275 ();
 sg13g2_decap_8 FILLER_6_1282 ();
 sg13g2_decap_8 FILLER_6_1289 ();
 sg13g2_decap_8 FILLER_6_1296 ();
 sg13g2_decap_8 FILLER_6_1303 ();
 sg13g2_decap_8 FILLER_6_1310 ();
 sg13g2_decap_8 FILLER_6_1317 ();
 sg13g2_decap_8 FILLER_6_1324 ();
 sg13g2_decap_8 FILLER_6_1331 ();
 sg13g2_decap_8 FILLER_6_1338 ();
 sg13g2_decap_8 FILLER_6_1345 ();
 sg13g2_decap_8 FILLER_6_1352 ();
 sg13g2_decap_8 FILLER_6_1359 ();
 sg13g2_decap_8 FILLER_6_1366 ();
 sg13g2_decap_8 FILLER_6_1373 ();
 sg13g2_decap_8 FILLER_6_1380 ();
 sg13g2_decap_8 FILLER_6_1387 ();
 sg13g2_decap_8 FILLER_6_1394 ();
 sg13g2_decap_8 FILLER_6_1401 ();
 sg13g2_decap_8 FILLER_6_1408 ();
 sg13g2_decap_8 FILLER_6_1415 ();
 sg13g2_decap_8 FILLER_6_1422 ();
 sg13g2_decap_8 FILLER_6_1429 ();
 sg13g2_decap_8 FILLER_6_1436 ();
 sg13g2_decap_8 FILLER_6_1443 ();
 sg13g2_decap_8 FILLER_6_1450 ();
 sg13g2_decap_8 FILLER_6_1457 ();
 sg13g2_decap_8 FILLER_6_1464 ();
 sg13g2_decap_8 FILLER_6_1471 ();
 sg13g2_decap_8 FILLER_6_1478 ();
 sg13g2_decap_8 FILLER_6_1485 ();
 sg13g2_decap_8 FILLER_6_1492 ();
 sg13g2_decap_8 FILLER_6_1499 ();
 sg13g2_decap_8 FILLER_6_1506 ();
 sg13g2_decap_8 FILLER_6_1513 ();
 sg13g2_decap_8 FILLER_6_1520 ();
 sg13g2_decap_8 FILLER_6_1527 ();
 sg13g2_decap_8 FILLER_6_1534 ();
 sg13g2_decap_8 FILLER_6_1541 ();
 sg13g2_decap_8 FILLER_6_1548 ();
 sg13g2_decap_8 FILLER_6_1555 ();
 sg13g2_decap_8 FILLER_6_1562 ();
 sg13g2_decap_8 FILLER_6_1569 ();
 sg13g2_decap_8 FILLER_6_1576 ();
 sg13g2_decap_8 FILLER_6_1583 ();
 sg13g2_decap_8 FILLER_6_1590 ();
 sg13g2_decap_8 FILLER_6_1597 ();
 sg13g2_decap_8 FILLER_6_1604 ();
 sg13g2_decap_8 FILLER_6_1611 ();
 sg13g2_decap_8 FILLER_6_1618 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_4 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_467 ();
 sg13g2_decap_8 FILLER_7_495 ();
 sg13g2_decap_8 FILLER_7_502 ();
 sg13g2_decap_8 FILLER_7_509 ();
 sg13g2_decap_8 FILLER_7_516 ();
 sg13g2_fill_2 FILLER_7_523 ();
 sg13g2_fill_1 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_530 ();
 sg13g2_decap_8 FILLER_7_537 ();
 sg13g2_decap_8 FILLER_7_544 ();
 sg13g2_decap_8 FILLER_7_551 ();
 sg13g2_decap_8 FILLER_7_558 ();
 sg13g2_decap_8 FILLER_7_565 ();
 sg13g2_decap_4 FILLER_7_572 ();
 sg13g2_decap_4 FILLER_7_580 ();
 sg13g2_decap_4 FILLER_7_587 ();
 sg13g2_fill_2 FILLER_7_591 ();
 sg13g2_decap_4 FILLER_7_601 ();
 sg13g2_fill_2 FILLER_7_605 ();
 sg13g2_decap_8 FILLER_7_611 ();
 sg13g2_decap_4 FILLER_7_618 ();
 sg13g2_decap_4 FILLER_7_643 ();
 sg13g2_fill_1 FILLER_7_647 ();
 sg13g2_decap_8 FILLER_7_669 ();
 sg13g2_decap_8 FILLER_7_676 ();
 sg13g2_decap_8 FILLER_7_683 ();
 sg13g2_fill_1 FILLER_7_690 ();
 sg13g2_decap_8 FILLER_7_695 ();
 sg13g2_decap_8 FILLER_7_702 ();
 sg13g2_fill_1 FILLER_7_709 ();
 sg13g2_decap_8 FILLER_7_744 ();
 sg13g2_decap_4 FILLER_7_751 ();
 sg13g2_decap_8 FILLER_7_759 ();
 sg13g2_fill_2 FILLER_7_766 ();
 sg13g2_fill_1 FILLER_7_768 ();
 sg13g2_fill_2 FILLER_7_772 ();
 sg13g2_decap_8 FILLER_7_778 ();
 sg13g2_decap_4 FILLER_7_785 ();
 sg13g2_fill_2 FILLER_7_846 ();
 sg13g2_decap_8 FILLER_7_857 ();
 sg13g2_fill_1 FILLER_7_864 ();
 sg13g2_decap_4 FILLER_7_900 ();
 sg13g2_decap_8 FILLER_7_908 ();
 sg13g2_decap_4 FILLER_7_915 ();
 sg13g2_fill_2 FILLER_7_961 ();
 sg13g2_fill_1 FILLER_7_963 ();
 sg13g2_decap_8 FILLER_7_1019 ();
 sg13g2_decap_8 FILLER_7_1026 ();
 sg13g2_fill_1 FILLER_7_1033 ();
 sg13g2_fill_2 FILLER_7_1060 ();
 sg13g2_decap_8 FILLER_7_1083 ();
 sg13g2_decap_8 FILLER_7_1090 ();
 sg13g2_fill_2 FILLER_7_1097 ();
 sg13g2_decap_8 FILLER_7_1103 ();
 sg13g2_fill_2 FILLER_7_1110 ();
 sg13g2_fill_1 FILLER_7_1112 ();
 sg13g2_decap_8 FILLER_7_1134 ();
 sg13g2_fill_1 FILLER_7_1141 ();
 sg13g2_decap_8 FILLER_7_1146 ();
 sg13g2_decap_8 FILLER_7_1153 ();
 sg13g2_decap_8 FILLER_7_1160 ();
 sg13g2_decap_8 FILLER_7_1167 ();
 sg13g2_decap_8 FILLER_7_1174 ();
 sg13g2_decap_8 FILLER_7_1181 ();
 sg13g2_decap_8 FILLER_7_1188 ();
 sg13g2_decap_8 FILLER_7_1195 ();
 sg13g2_decap_8 FILLER_7_1202 ();
 sg13g2_decap_8 FILLER_7_1209 ();
 sg13g2_decap_8 FILLER_7_1216 ();
 sg13g2_decap_8 FILLER_7_1223 ();
 sg13g2_decap_8 FILLER_7_1230 ();
 sg13g2_decap_8 FILLER_7_1237 ();
 sg13g2_decap_8 FILLER_7_1244 ();
 sg13g2_decap_8 FILLER_7_1251 ();
 sg13g2_decap_8 FILLER_7_1258 ();
 sg13g2_decap_8 FILLER_7_1265 ();
 sg13g2_decap_8 FILLER_7_1272 ();
 sg13g2_decap_8 FILLER_7_1279 ();
 sg13g2_decap_8 FILLER_7_1286 ();
 sg13g2_decap_8 FILLER_7_1293 ();
 sg13g2_decap_8 FILLER_7_1300 ();
 sg13g2_decap_8 FILLER_7_1307 ();
 sg13g2_decap_8 FILLER_7_1314 ();
 sg13g2_decap_8 FILLER_7_1321 ();
 sg13g2_decap_8 FILLER_7_1328 ();
 sg13g2_decap_8 FILLER_7_1335 ();
 sg13g2_decap_8 FILLER_7_1342 ();
 sg13g2_decap_8 FILLER_7_1349 ();
 sg13g2_decap_8 FILLER_7_1356 ();
 sg13g2_decap_8 FILLER_7_1363 ();
 sg13g2_decap_8 FILLER_7_1370 ();
 sg13g2_decap_8 FILLER_7_1377 ();
 sg13g2_decap_8 FILLER_7_1384 ();
 sg13g2_decap_8 FILLER_7_1391 ();
 sg13g2_decap_8 FILLER_7_1398 ();
 sg13g2_decap_8 FILLER_7_1405 ();
 sg13g2_decap_8 FILLER_7_1412 ();
 sg13g2_decap_8 FILLER_7_1419 ();
 sg13g2_decap_8 FILLER_7_1426 ();
 sg13g2_decap_8 FILLER_7_1433 ();
 sg13g2_decap_8 FILLER_7_1440 ();
 sg13g2_decap_8 FILLER_7_1447 ();
 sg13g2_decap_8 FILLER_7_1454 ();
 sg13g2_decap_8 FILLER_7_1461 ();
 sg13g2_decap_8 FILLER_7_1468 ();
 sg13g2_decap_8 FILLER_7_1475 ();
 sg13g2_decap_8 FILLER_7_1482 ();
 sg13g2_decap_8 FILLER_7_1489 ();
 sg13g2_decap_8 FILLER_7_1496 ();
 sg13g2_decap_8 FILLER_7_1503 ();
 sg13g2_decap_8 FILLER_7_1510 ();
 sg13g2_decap_8 FILLER_7_1517 ();
 sg13g2_decap_8 FILLER_7_1524 ();
 sg13g2_decap_8 FILLER_7_1531 ();
 sg13g2_decap_8 FILLER_7_1538 ();
 sg13g2_decap_8 FILLER_7_1545 ();
 sg13g2_decap_8 FILLER_7_1552 ();
 sg13g2_decap_8 FILLER_7_1559 ();
 sg13g2_decap_8 FILLER_7_1566 ();
 sg13g2_decap_8 FILLER_7_1573 ();
 sg13g2_decap_8 FILLER_7_1580 ();
 sg13g2_decap_8 FILLER_7_1587 ();
 sg13g2_decap_8 FILLER_7_1594 ();
 sg13g2_decap_8 FILLER_7_1601 ();
 sg13g2_decap_8 FILLER_7_1608 ();
 sg13g2_decap_8 FILLER_7_1615 ();
 sg13g2_fill_2 FILLER_7_1622 ();
 sg13g2_fill_1 FILLER_7_1624 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_4 FILLER_8_350 ();
 sg13g2_fill_1 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_decap_4 FILLER_8_366 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_fill_2 FILLER_8_400 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_4 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_421 ();
 sg13g2_decap_4 FILLER_8_437 ();
 sg13g2_fill_2 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_464 ();
 sg13g2_decap_8 FILLER_8_471 ();
 sg13g2_decap_8 FILLER_8_478 ();
 sg13g2_decap_8 FILLER_8_485 ();
 sg13g2_decap_8 FILLER_8_513 ();
 sg13g2_fill_2 FILLER_8_520 ();
 sg13g2_fill_1 FILLER_8_522 ();
 sg13g2_fill_1 FILLER_8_563 ();
 sg13g2_decap_8 FILLER_8_568 ();
 sg13g2_decap_8 FILLER_8_575 ();
 sg13g2_decap_8 FILLER_8_582 ();
 sg13g2_fill_1 FILLER_8_589 ();
 sg13g2_fill_2 FILLER_8_594 ();
 sg13g2_decap_8 FILLER_8_601 ();
 sg13g2_decap_8 FILLER_8_608 ();
 sg13g2_fill_2 FILLER_8_615 ();
 sg13g2_fill_1 FILLER_8_617 ();
 sg13g2_decap_8 FILLER_8_622 ();
 sg13g2_fill_2 FILLER_8_629 ();
 sg13g2_fill_1 FILLER_8_631 ();
 sg13g2_decap_8 FILLER_8_653 ();
 sg13g2_decap_8 FILLER_8_660 ();
 sg13g2_fill_2 FILLER_8_667 ();
 sg13g2_fill_1 FILLER_8_669 ();
 sg13g2_fill_2 FILLER_8_710 ();
 sg13g2_fill_1 FILLER_8_712 ();
 sg13g2_fill_1 FILLER_8_742 ();
 sg13g2_fill_1 FILLER_8_794 ();
 sg13g2_fill_2 FILLER_8_845 ();
 sg13g2_decap_8 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_8_884 ();
 sg13g2_decap_8 FILLER_8_891 ();
 sg13g2_decap_8 FILLER_8_898 ();
 sg13g2_decap_8 FILLER_8_905 ();
 sg13g2_fill_2 FILLER_8_912 ();
 sg13g2_fill_1 FILLER_8_939 ();
 sg13g2_fill_1 FILLER_8_961 ();
 sg13g2_decap_4 FILLER_8_966 ();
 sg13g2_fill_2 FILLER_8_970 ();
 sg13g2_fill_1 FILLER_8_1002 ();
 sg13g2_decap_8 FILLER_8_1028 ();
 sg13g2_fill_2 FILLER_8_1035 ();
 sg13g2_fill_1 FILLER_8_1037 ();
 sg13g2_decap_8 FILLER_8_1043 ();
 sg13g2_decap_4 FILLER_8_1050 ();
 sg13g2_fill_1 FILLER_8_1054 ();
 sg13g2_decap_8 FILLER_8_1059 ();
 sg13g2_decap_8 FILLER_8_1066 ();
 sg13g2_fill_2 FILLER_8_1073 ();
 sg13g2_fill_1 FILLER_8_1075 ();
 sg13g2_decap_8 FILLER_8_1111 ();
 sg13g2_decap_4 FILLER_8_1118 ();
 sg13g2_fill_2 FILLER_8_1131 ();
 sg13g2_fill_1 FILLER_8_1133 ();
 sg13g2_decap_8 FILLER_8_1160 ();
 sg13g2_decap_8 FILLER_8_1167 ();
 sg13g2_decap_8 FILLER_8_1174 ();
 sg13g2_decap_8 FILLER_8_1181 ();
 sg13g2_decap_8 FILLER_8_1188 ();
 sg13g2_decap_8 FILLER_8_1195 ();
 sg13g2_decap_8 FILLER_8_1202 ();
 sg13g2_decap_8 FILLER_8_1209 ();
 sg13g2_decap_8 FILLER_8_1216 ();
 sg13g2_decap_8 FILLER_8_1223 ();
 sg13g2_decap_8 FILLER_8_1230 ();
 sg13g2_decap_8 FILLER_8_1237 ();
 sg13g2_decap_8 FILLER_8_1244 ();
 sg13g2_decap_8 FILLER_8_1251 ();
 sg13g2_decap_8 FILLER_8_1258 ();
 sg13g2_decap_8 FILLER_8_1265 ();
 sg13g2_decap_8 FILLER_8_1272 ();
 sg13g2_decap_8 FILLER_8_1279 ();
 sg13g2_decap_8 FILLER_8_1286 ();
 sg13g2_decap_8 FILLER_8_1293 ();
 sg13g2_decap_8 FILLER_8_1300 ();
 sg13g2_decap_8 FILLER_8_1307 ();
 sg13g2_decap_8 FILLER_8_1314 ();
 sg13g2_decap_8 FILLER_8_1321 ();
 sg13g2_decap_8 FILLER_8_1328 ();
 sg13g2_decap_8 FILLER_8_1335 ();
 sg13g2_decap_8 FILLER_8_1342 ();
 sg13g2_decap_8 FILLER_8_1349 ();
 sg13g2_decap_8 FILLER_8_1356 ();
 sg13g2_decap_8 FILLER_8_1363 ();
 sg13g2_decap_8 FILLER_8_1370 ();
 sg13g2_decap_8 FILLER_8_1377 ();
 sg13g2_decap_8 FILLER_8_1384 ();
 sg13g2_decap_8 FILLER_8_1391 ();
 sg13g2_decap_8 FILLER_8_1398 ();
 sg13g2_decap_8 FILLER_8_1405 ();
 sg13g2_decap_8 FILLER_8_1412 ();
 sg13g2_decap_8 FILLER_8_1419 ();
 sg13g2_decap_8 FILLER_8_1426 ();
 sg13g2_decap_8 FILLER_8_1433 ();
 sg13g2_decap_8 FILLER_8_1440 ();
 sg13g2_decap_8 FILLER_8_1447 ();
 sg13g2_decap_8 FILLER_8_1454 ();
 sg13g2_decap_8 FILLER_8_1461 ();
 sg13g2_decap_8 FILLER_8_1468 ();
 sg13g2_decap_8 FILLER_8_1475 ();
 sg13g2_decap_8 FILLER_8_1482 ();
 sg13g2_decap_8 FILLER_8_1489 ();
 sg13g2_decap_8 FILLER_8_1496 ();
 sg13g2_decap_8 FILLER_8_1503 ();
 sg13g2_decap_8 FILLER_8_1510 ();
 sg13g2_decap_8 FILLER_8_1517 ();
 sg13g2_decap_8 FILLER_8_1524 ();
 sg13g2_decap_8 FILLER_8_1531 ();
 sg13g2_decap_8 FILLER_8_1538 ();
 sg13g2_decap_8 FILLER_8_1545 ();
 sg13g2_decap_8 FILLER_8_1552 ();
 sg13g2_decap_8 FILLER_8_1559 ();
 sg13g2_decap_8 FILLER_8_1566 ();
 sg13g2_decap_8 FILLER_8_1573 ();
 sg13g2_decap_8 FILLER_8_1580 ();
 sg13g2_decap_8 FILLER_8_1587 ();
 sg13g2_decap_8 FILLER_8_1594 ();
 sg13g2_decap_8 FILLER_8_1601 ();
 sg13g2_decap_8 FILLER_8_1608 ();
 sg13g2_decap_8 FILLER_8_1615 ();
 sg13g2_fill_2 FILLER_8_1622 ();
 sg13g2_fill_1 FILLER_8_1624 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_fill_2 FILLER_9_315 ();
 sg13g2_fill_1 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_337 ();
 sg13g2_decap_4 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_374 ();
 sg13g2_fill_2 FILLER_9_381 ();
 sg13g2_fill_1 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_fill_1 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_4 FILLER_9_424 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_fill_1 FILLER_9_435 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_8 FILLER_9_466 ();
 sg13g2_fill_1 FILLER_9_473 ();
 sg13g2_decap_4 FILLER_9_478 ();
 sg13g2_fill_1 FILLER_9_482 ();
 sg13g2_decap_8 FILLER_9_492 ();
 sg13g2_decap_8 FILLER_9_499 ();
 sg13g2_fill_1 FILLER_9_506 ();
 sg13g2_decap_8 FILLER_9_528 ();
 sg13g2_decap_4 FILLER_9_535 ();
 sg13g2_fill_2 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_545 ();
 sg13g2_fill_2 FILLER_9_552 ();
 sg13g2_fill_2 FILLER_9_580 ();
 sg13g2_fill_2 FILLER_9_608 ();
 sg13g2_fill_1 FILLER_9_610 ();
 sg13g2_fill_1 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_659 ();
 sg13g2_decap_4 FILLER_9_666 ();
 sg13g2_decap_8 FILLER_9_674 ();
 sg13g2_decap_8 FILLER_9_681 ();
 sg13g2_fill_2 FILLER_9_697 ();
 sg13g2_fill_2 FILLER_9_756 ();
 sg13g2_fill_1 FILLER_9_758 ();
 sg13g2_fill_1 FILLER_9_764 ();
 sg13g2_fill_1 FILLER_9_837 ();
 sg13g2_decap_4 FILLER_9_893 ();
 sg13g2_fill_2 FILLER_9_901 ();
 sg13g2_fill_1 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_913 ();
 sg13g2_decap_8 FILLER_9_920 ();
 sg13g2_decap_8 FILLER_9_927 ();
 sg13g2_decap_4 FILLER_9_934 ();
 sg13g2_decap_4 FILLER_9_972 ();
 sg13g2_fill_1 FILLER_9_976 ();
 sg13g2_fill_1 FILLER_9_1007 ();
 sg13g2_decap_8 FILLER_9_1033 ();
 sg13g2_decap_8 FILLER_9_1040 ();
 sg13g2_fill_2 FILLER_9_1047 ();
 sg13g2_fill_1 FILLER_9_1049 ();
 sg13g2_decap_8 FILLER_9_1071 ();
 sg13g2_decap_8 FILLER_9_1078 ();
 sg13g2_decap_8 FILLER_9_1085 ();
 sg13g2_fill_1 FILLER_9_1092 ();
 sg13g2_decap_8 FILLER_9_1097 ();
 sg13g2_decap_4 FILLER_9_1104 ();
 sg13g2_fill_1 FILLER_9_1108 ();
 sg13g2_decap_8 FILLER_9_1130 ();
 sg13g2_decap_8 FILLER_9_1137 ();
 sg13g2_decap_8 FILLER_9_1144 ();
 sg13g2_decap_8 FILLER_9_1151 ();
 sg13g2_decap_8 FILLER_9_1158 ();
 sg13g2_decap_8 FILLER_9_1165 ();
 sg13g2_decap_8 FILLER_9_1172 ();
 sg13g2_decap_8 FILLER_9_1179 ();
 sg13g2_decap_8 FILLER_9_1186 ();
 sg13g2_decap_8 FILLER_9_1193 ();
 sg13g2_decap_8 FILLER_9_1200 ();
 sg13g2_decap_8 FILLER_9_1207 ();
 sg13g2_decap_8 FILLER_9_1214 ();
 sg13g2_decap_8 FILLER_9_1221 ();
 sg13g2_decap_8 FILLER_9_1228 ();
 sg13g2_decap_8 FILLER_9_1235 ();
 sg13g2_decap_8 FILLER_9_1242 ();
 sg13g2_decap_8 FILLER_9_1249 ();
 sg13g2_decap_8 FILLER_9_1256 ();
 sg13g2_decap_8 FILLER_9_1263 ();
 sg13g2_decap_8 FILLER_9_1270 ();
 sg13g2_decap_8 FILLER_9_1277 ();
 sg13g2_decap_8 FILLER_9_1284 ();
 sg13g2_decap_8 FILLER_9_1291 ();
 sg13g2_decap_8 FILLER_9_1298 ();
 sg13g2_decap_8 FILLER_9_1305 ();
 sg13g2_decap_8 FILLER_9_1312 ();
 sg13g2_decap_8 FILLER_9_1319 ();
 sg13g2_decap_8 FILLER_9_1326 ();
 sg13g2_decap_8 FILLER_9_1333 ();
 sg13g2_decap_8 FILLER_9_1340 ();
 sg13g2_decap_8 FILLER_9_1347 ();
 sg13g2_decap_8 FILLER_9_1354 ();
 sg13g2_decap_8 FILLER_9_1361 ();
 sg13g2_decap_8 FILLER_9_1368 ();
 sg13g2_decap_8 FILLER_9_1375 ();
 sg13g2_decap_8 FILLER_9_1382 ();
 sg13g2_decap_8 FILLER_9_1389 ();
 sg13g2_decap_8 FILLER_9_1396 ();
 sg13g2_decap_8 FILLER_9_1403 ();
 sg13g2_decap_8 FILLER_9_1410 ();
 sg13g2_decap_8 FILLER_9_1417 ();
 sg13g2_decap_8 FILLER_9_1424 ();
 sg13g2_decap_8 FILLER_9_1431 ();
 sg13g2_decap_8 FILLER_9_1438 ();
 sg13g2_decap_8 FILLER_9_1445 ();
 sg13g2_decap_8 FILLER_9_1452 ();
 sg13g2_decap_8 FILLER_9_1459 ();
 sg13g2_decap_8 FILLER_9_1466 ();
 sg13g2_decap_8 FILLER_9_1473 ();
 sg13g2_decap_8 FILLER_9_1480 ();
 sg13g2_decap_8 FILLER_9_1487 ();
 sg13g2_decap_8 FILLER_9_1494 ();
 sg13g2_decap_8 FILLER_9_1501 ();
 sg13g2_decap_8 FILLER_9_1508 ();
 sg13g2_decap_8 FILLER_9_1515 ();
 sg13g2_decap_8 FILLER_9_1522 ();
 sg13g2_decap_8 FILLER_9_1529 ();
 sg13g2_decap_8 FILLER_9_1536 ();
 sg13g2_decap_8 FILLER_9_1543 ();
 sg13g2_decap_8 FILLER_9_1550 ();
 sg13g2_decap_8 FILLER_9_1557 ();
 sg13g2_decap_8 FILLER_9_1564 ();
 sg13g2_decap_8 FILLER_9_1571 ();
 sg13g2_decap_8 FILLER_9_1578 ();
 sg13g2_decap_8 FILLER_9_1585 ();
 sg13g2_decap_8 FILLER_9_1592 ();
 sg13g2_decap_8 FILLER_9_1599 ();
 sg13g2_decap_8 FILLER_9_1606 ();
 sg13g2_decap_8 FILLER_9_1613 ();
 sg13g2_decap_4 FILLER_9_1620 ();
 sg13g2_fill_1 FILLER_9_1624 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_4 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_4 FILLER_10_338 ();
 sg13g2_fill_2 FILLER_10_342 ();
 sg13g2_fill_2 FILLER_10_362 ();
 sg13g2_fill_1 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_fill_2 FILLER_10_424 ();
 sg13g2_fill_2 FILLER_10_435 ();
 sg13g2_fill_1 FILLER_10_498 ();
 sg13g2_decap_8 FILLER_10_507 ();
 sg13g2_decap_4 FILLER_10_514 ();
 sg13g2_decap_8 FILLER_10_522 ();
 sg13g2_fill_2 FILLER_10_529 ();
 sg13g2_decap_8 FILLER_10_535 ();
 sg13g2_decap_8 FILLER_10_542 ();
 sg13g2_decap_8 FILLER_10_549 ();
 sg13g2_fill_2 FILLER_10_556 ();
 sg13g2_decap_4 FILLER_10_567 ();
 sg13g2_fill_2 FILLER_10_575 ();
 sg13g2_fill_1 FILLER_10_577 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_fill_1 FILLER_10_630 ();
 sg13g2_fill_2 FILLER_10_635 ();
 sg13g2_fill_1 FILLER_10_637 ();
 sg13g2_fill_2 FILLER_10_659 ();
 sg13g2_fill_2 FILLER_10_687 ();
 sg13g2_fill_2 FILLER_10_836 ();
 sg13g2_fill_2 FILLER_10_864 ();
 sg13g2_fill_1 FILLER_10_866 ();
 sg13g2_fill_2 FILLER_10_888 ();
 sg13g2_fill_1 FILLER_10_921 ();
 sg13g2_decap_4 FILLER_10_926 ();
 sg13g2_fill_1 FILLER_10_930 ();
 sg13g2_fill_2 FILLER_10_1031 ();
 sg13g2_decap_4 FILLER_10_1046 ();
 sg13g2_decap_8 FILLER_10_1071 ();
 sg13g2_fill_2 FILLER_10_1078 ();
 sg13g2_fill_2 FILLER_10_1091 ();
 sg13g2_decap_8 FILLER_10_1118 ();
 sg13g2_decap_8 FILLER_10_1125 ();
 sg13g2_fill_1 FILLER_10_1137 ();
 sg13g2_decap_8 FILLER_10_1142 ();
 sg13g2_decap_8 FILLER_10_1149 ();
 sg13g2_decap_8 FILLER_10_1156 ();
 sg13g2_fill_1 FILLER_10_1163 ();
 sg13g2_decap_8 FILLER_10_1168 ();
 sg13g2_decap_8 FILLER_10_1175 ();
 sg13g2_decap_8 FILLER_10_1182 ();
 sg13g2_decap_8 FILLER_10_1189 ();
 sg13g2_decap_8 FILLER_10_1196 ();
 sg13g2_decap_8 FILLER_10_1203 ();
 sg13g2_decap_8 FILLER_10_1210 ();
 sg13g2_decap_8 FILLER_10_1217 ();
 sg13g2_decap_8 FILLER_10_1224 ();
 sg13g2_decap_8 FILLER_10_1231 ();
 sg13g2_decap_8 FILLER_10_1238 ();
 sg13g2_decap_8 FILLER_10_1245 ();
 sg13g2_decap_8 FILLER_10_1252 ();
 sg13g2_decap_8 FILLER_10_1259 ();
 sg13g2_decap_8 FILLER_10_1266 ();
 sg13g2_decap_8 FILLER_10_1273 ();
 sg13g2_decap_8 FILLER_10_1280 ();
 sg13g2_decap_8 FILLER_10_1287 ();
 sg13g2_decap_8 FILLER_10_1294 ();
 sg13g2_decap_8 FILLER_10_1301 ();
 sg13g2_decap_8 FILLER_10_1308 ();
 sg13g2_decap_8 FILLER_10_1315 ();
 sg13g2_decap_8 FILLER_10_1322 ();
 sg13g2_decap_8 FILLER_10_1329 ();
 sg13g2_decap_8 FILLER_10_1336 ();
 sg13g2_decap_8 FILLER_10_1343 ();
 sg13g2_decap_8 FILLER_10_1350 ();
 sg13g2_decap_8 FILLER_10_1357 ();
 sg13g2_decap_8 FILLER_10_1364 ();
 sg13g2_decap_8 FILLER_10_1371 ();
 sg13g2_decap_8 FILLER_10_1378 ();
 sg13g2_decap_8 FILLER_10_1385 ();
 sg13g2_decap_8 FILLER_10_1392 ();
 sg13g2_decap_8 FILLER_10_1399 ();
 sg13g2_decap_8 FILLER_10_1406 ();
 sg13g2_decap_8 FILLER_10_1413 ();
 sg13g2_decap_8 FILLER_10_1420 ();
 sg13g2_decap_8 FILLER_10_1427 ();
 sg13g2_decap_8 FILLER_10_1434 ();
 sg13g2_decap_8 FILLER_10_1441 ();
 sg13g2_decap_8 FILLER_10_1448 ();
 sg13g2_decap_8 FILLER_10_1455 ();
 sg13g2_decap_8 FILLER_10_1462 ();
 sg13g2_decap_8 FILLER_10_1469 ();
 sg13g2_decap_8 FILLER_10_1476 ();
 sg13g2_decap_8 FILLER_10_1483 ();
 sg13g2_decap_8 FILLER_10_1490 ();
 sg13g2_decap_8 FILLER_10_1497 ();
 sg13g2_decap_8 FILLER_10_1504 ();
 sg13g2_decap_8 FILLER_10_1511 ();
 sg13g2_decap_8 FILLER_10_1518 ();
 sg13g2_decap_8 FILLER_10_1525 ();
 sg13g2_decap_8 FILLER_10_1532 ();
 sg13g2_decap_8 FILLER_10_1539 ();
 sg13g2_decap_8 FILLER_10_1546 ();
 sg13g2_decap_8 FILLER_10_1553 ();
 sg13g2_decap_8 FILLER_10_1560 ();
 sg13g2_decap_8 FILLER_10_1567 ();
 sg13g2_decap_8 FILLER_10_1574 ();
 sg13g2_decap_8 FILLER_10_1581 ();
 sg13g2_decap_8 FILLER_10_1588 ();
 sg13g2_decap_8 FILLER_10_1595 ();
 sg13g2_decap_8 FILLER_10_1602 ();
 sg13g2_decap_8 FILLER_10_1609 ();
 sg13g2_decap_8 FILLER_10_1616 ();
 sg13g2_fill_2 FILLER_10_1623 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_4 FILLER_11_336 ();
 sg13g2_fill_2 FILLER_11_418 ();
 sg13g2_decap_8 FILLER_11_449 ();
 sg13g2_decap_8 FILLER_11_456 ();
 sg13g2_decap_4 FILLER_11_463 ();
 sg13g2_fill_1 FILLER_11_549 ();
 sg13g2_decap_4 FILLER_11_611 ();
 sg13g2_fill_1 FILLER_11_615 ();
 sg13g2_decap_8 FILLER_11_641 ();
 sg13g2_decap_4 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_661 ();
 sg13g2_decap_8 FILLER_11_668 ();
 sg13g2_decap_4 FILLER_11_675 ();
 sg13g2_fill_2 FILLER_11_679 ();
 sg13g2_fill_1 FILLER_11_716 ();
 sg13g2_decap_4 FILLER_11_722 ();
 sg13g2_fill_2 FILLER_11_726 ();
 sg13g2_decap_8 FILLER_11_732 ();
 sg13g2_fill_2 FILLER_11_739 ();
 sg13g2_fill_1 FILLER_11_741 ();
 sg13g2_decap_4 FILLER_11_776 ();
 sg13g2_fill_2 FILLER_11_780 ();
 sg13g2_decap_8 FILLER_11_786 ();
 sg13g2_decap_8 FILLER_11_793 ();
 sg13g2_fill_1 FILLER_11_800 ();
 sg13g2_fill_2 FILLER_11_810 ();
 sg13g2_fill_2 FILLER_11_841 ();
 sg13g2_fill_1 FILLER_11_843 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_8 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_11_865 ();
 sg13g2_decap_8 FILLER_11_872 ();
 sg13g2_decap_8 FILLER_11_879 ();
 sg13g2_decap_8 FILLER_11_886 ();
 sg13g2_decap_8 FILLER_11_893 ();
 sg13g2_fill_2 FILLER_11_900 ();
 sg13g2_fill_1 FILLER_11_902 ();
 sg13g2_decap_4 FILLER_11_911 ();
 sg13g2_fill_2 FILLER_11_956 ();
 sg13g2_fill_1 FILLER_11_958 ();
 sg13g2_fill_2 FILLER_11_990 ();
 sg13g2_fill_1 FILLER_11_1005 ();
 sg13g2_decap_8 FILLER_11_1053 ();
 sg13g2_fill_2 FILLER_11_1060 ();
 sg13g2_fill_1 FILLER_11_1062 ();
 sg13g2_fill_2 FILLER_11_1098 ();
 sg13g2_decap_4 FILLER_11_1104 ();
 sg13g2_fill_1 FILLER_11_1108 ();
 sg13g2_fill_1 FILLER_11_1130 ();
 sg13g2_decap_8 FILLER_11_1183 ();
 sg13g2_decap_8 FILLER_11_1190 ();
 sg13g2_decap_8 FILLER_11_1197 ();
 sg13g2_decap_8 FILLER_11_1204 ();
 sg13g2_decap_8 FILLER_11_1211 ();
 sg13g2_decap_8 FILLER_11_1218 ();
 sg13g2_decap_8 FILLER_11_1225 ();
 sg13g2_decap_8 FILLER_11_1232 ();
 sg13g2_decap_8 FILLER_11_1239 ();
 sg13g2_decap_8 FILLER_11_1246 ();
 sg13g2_decap_8 FILLER_11_1253 ();
 sg13g2_decap_8 FILLER_11_1260 ();
 sg13g2_decap_8 FILLER_11_1267 ();
 sg13g2_decap_8 FILLER_11_1274 ();
 sg13g2_decap_8 FILLER_11_1281 ();
 sg13g2_decap_8 FILLER_11_1288 ();
 sg13g2_decap_8 FILLER_11_1295 ();
 sg13g2_decap_8 FILLER_11_1302 ();
 sg13g2_decap_8 FILLER_11_1309 ();
 sg13g2_decap_8 FILLER_11_1316 ();
 sg13g2_decap_8 FILLER_11_1323 ();
 sg13g2_decap_8 FILLER_11_1330 ();
 sg13g2_decap_8 FILLER_11_1337 ();
 sg13g2_decap_8 FILLER_11_1344 ();
 sg13g2_decap_8 FILLER_11_1351 ();
 sg13g2_decap_8 FILLER_11_1358 ();
 sg13g2_decap_8 FILLER_11_1365 ();
 sg13g2_decap_8 FILLER_11_1372 ();
 sg13g2_decap_8 FILLER_11_1379 ();
 sg13g2_decap_8 FILLER_11_1386 ();
 sg13g2_decap_8 FILLER_11_1393 ();
 sg13g2_decap_8 FILLER_11_1400 ();
 sg13g2_decap_8 FILLER_11_1407 ();
 sg13g2_decap_8 FILLER_11_1414 ();
 sg13g2_decap_8 FILLER_11_1421 ();
 sg13g2_decap_8 FILLER_11_1428 ();
 sg13g2_decap_8 FILLER_11_1435 ();
 sg13g2_decap_8 FILLER_11_1442 ();
 sg13g2_decap_8 FILLER_11_1449 ();
 sg13g2_decap_8 FILLER_11_1456 ();
 sg13g2_decap_8 FILLER_11_1463 ();
 sg13g2_decap_8 FILLER_11_1470 ();
 sg13g2_decap_8 FILLER_11_1477 ();
 sg13g2_decap_8 FILLER_11_1484 ();
 sg13g2_decap_8 FILLER_11_1491 ();
 sg13g2_decap_8 FILLER_11_1498 ();
 sg13g2_decap_8 FILLER_11_1505 ();
 sg13g2_decap_8 FILLER_11_1512 ();
 sg13g2_decap_8 FILLER_11_1519 ();
 sg13g2_decap_8 FILLER_11_1526 ();
 sg13g2_decap_8 FILLER_11_1533 ();
 sg13g2_decap_8 FILLER_11_1540 ();
 sg13g2_decap_8 FILLER_11_1547 ();
 sg13g2_decap_8 FILLER_11_1554 ();
 sg13g2_decap_8 FILLER_11_1561 ();
 sg13g2_decap_8 FILLER_11_1568 ();
 sg13g2_decap_8 FILLER_11_1575 ();
 sg13g2_decap_8 FILLER_11_1582 ();
 sg13g2_decap_8 FILLER_11_1589 ();
 sg13g2_decap_8 FILLER_11_1596 ();
 sg13g2_decap_8 FILLER_11_1603 ();
 sg13g2_decap_8 FILLER_11_1610 ();
 sg13g2_decap_8 FILLER_11_1617 ();
 sg13g2_fill_1 FILLER_11_1624 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_4 FILLER_12_336 ();
 sg13g2_fill_2 FILLER_12_340 ();
 sg13g2_fill_2 FILLER_12_368 ();
 sg13g2_fill_1 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_12_414 ();
 sg13g2_decap_4 FILLER_12_421 ();
 sg13g2_fill_1 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_506 ();
 sg13g2_decap_8 FILLER_12_513 ();
 sg13g2_decap_8 FILLER_12_520 ();
 sg13g2_decap_8 FILLER_12_527 ();
 sg13g2_decap_8 FILLER_12_534 ();
 sg13g2_decap_8 FILLER_12_541 ();
 sg13g2_fill_2 FILLER_12_548 ();
 sg13g2_fill_1 FILLER_12_550 ();
 sg13g2_fill_2 FILLER_12_577 ();
 sg13g2_fill_1 FILLER_12_579 ();
 sg13g2_decap_4 FILLER_12_606 ();
 sg13g2_fill_1 FILLER_12_610 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_fill_2 FILLER_12_658 ();
 sg13g2_fill_2 FILLER_12_693 ();
 sg13g2_fill_1 FILLER_12_695 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_4 FILLER_12_707 ();
 sg13g2_fill_1 FILLER_12_711 ();
 sg13g2_decap_8 FILLER_12_717 ();
 sg13g2_fill_1 FILLER_12_724 ();
 sg13g2_decap_4 FILLER_12_746 ();
 sg13g2_fill_2 FILLER_12_785 ();
 sg13g2_decap_8 FILLER_12_796 ();
 sg13g2_decap_4 FILLER_12_803 ();
 sg13g2_fill_1 FILLER_12_807 ();
 sg13g2_decap_4 FILLER_12_812 ();
 sg13g2_fill_1 FILLER_12_816 ();
 sg13g2_decap_8 FILLER_12_859 ();
 sg13g2_fill_2 FILLER_12_892 ();
 sg13g2_fill_1 FILLER_12_894 ();
 sg13g2_decap_8 FILLER_12_899 ();
 sg13g2_fill_2 FILLER_12_956 ();
 sg13g2_decap_8 FILLER_12_967 ();
 sg13g2_fill_2 FILLER_12_974 ();
 sg13g2_fill_1 FILLER_12_976 ();
 sg13g2_decap_8 FILLER_12_1003 ();
 sg13g2_decap_8 FILLER_12_1010 ();
 sg13g2_decap_4 FILLER_12_1017 ();
 sg13g2_decap_8 FILLER_12_1046 ();
 sg13g2_decap_8 FILLER_12_1053 ();
 sg13g2_decap_4 FILLER_12_1060 ();
 sg13g2_fill_2 FILLER_12_1064 ();
 sg13g2_decap_8 FILLER_12_1071 ();
 sg13g2_decap_8 FILLER_12_1078 ();
 sg13g2_fill_2 FILLER_12_1085 ();
 sg13g2_decap_8 FILLER_12_1118 ();
 sg13g2_decap_4 FILLER_12_1125 ();
 sg13g2_decap_8 FILLER_12_1133 ();
 sg13g2_decap_8 FILLER_12_1140 ();
 sg13g2_decap_8 FILLER_12_1147 ();
 sg13g2_fill_2 FILLER_12_1154 ();
 sg13g2_fill_1 FILLER_12_1156 ();
 sg13g2_decap_8 FILLER_12_1186 ();
 sg13g2_fill_1 FILLER_12_1193 ();
 sg13g2_decap_8 FILLER_12_1198 ();
 sg13g2_decap_8 FILLER_12_1205 ();
 sg13g2_decap_8 FILLER_12_1212 ();
 sg13g2_decap_8 FILLER_12_1219 ();
 sg13g2_decap_8 FILLER_12_1226 ();
 sg13g2_decap_8 FILLER_12_1233 ();
 sg13g2_decap_8 FILLER_12_1240 ();
 sg13g2_decap_8 FILLER_12_1247 ();
 sg13g2_decap_8 FILLER_12_1254 ();
 sg13g2_decap_8 FILLER_12_1261 ();
 sg13g2_decap_8 FILLER_12_1268 ();
 sg13g2_decap_8 FILLER_12_1275 ();
 sg13g2_decap_8 FILLER_12_1282 ();
 sg13g2_decap_8 FILLER_12_1289 ();
 sg13g2_decap_8 FILLER_12_1296 ();
 sg13g2_decap_8 FILLER_12_1303 ();
 sg13g2_decap_8 FILLER_12_1310 ();
 sg13g2_decap_8 FILLER_12_1317 ();
 sg13g2_decap_8 FILLER_12_1324 ();
 sg13g2_decap_8 FILLER_12_1331 ();
 sg13g2_decap_8 FILLER_12_1338 ();
 sg13g2_decap_8 FILLER_12_1345 ();
 sg13g2_decap_8 FILLER_12_1352 ();
 sg13g2_decap_8 FILLER_12_1359 ();
 sg13g2_decap_8 FILLER_12_1366 ();
 sg13g2_decap_8 FILLER_12_1373 ();
 sg13g2_decap_8 FILLER_12_1380 ();
 sg13g2_decap_8 FILLER_12_1387 ();
 sg13g2_decap_8 FILLER_12_1394 ();
 sg13g2_decap_8 FILLER_12_1401 ();
 sg13g2_decap_8 FILLER_12_1408 ();
 sg13g2_decap_8 FILLER_12_1415 ();
 sg13g2_decap_8 FILLER_12_1422 ();
 sg13g2_decap_8 FILLER_12_1429 ();
 sg13g2_decap_8 FILLER_12_1436 ();
 sg13g2_decap_8 FILLER_12_1443 ();
 sg13g2_decap_8 FILLER_12_1450 ();
 sg13g2_decap_8 FILLER_12_1457 ();
 sg13g2_decap_8 FILLER_12_1464 ();
 sg13g2_decap_8 FILLER_12_1471 ();
 sg13g2_decap_8 FILLER_12_1478 ();
 sg13g2_decap_8 FILLER_12_1485 ();
 sg13g2_decap_8 FILLER_12_1492 ();
 sg13g2_decap_8 FILLER_12_1499 ();
 sg13g2_decap_8 FILLER_12_1506 ();
 sg13g2_decap_8 FILLER_12_1513 ();
 sg13g2_decap_8 FILLER_12_1520 ();
 sg13g2_decap_8 FILLER_12_1527 ();
 sg13g2_decap_8 FILLER_12_1534 ();
 sg13g2_decap_8 FILLER_12_1541 ();
 sg13g2_decap_8 FILLER_12_1548 ();
 sg13g2_decap_8 FILLER_12_1555 ();
 sg13g2_decap_8 FILLER_12_1562 ();
 sg13g2_decap_8 FILLER_12_1569 ();
 sg13g2_decap_8 FILLER_12_1576 ();
 sg13g2_decap_8 FILLER_12_1583 ();
 sg13g2_decap_8 FILLER_12_1590 ();
 sg13g2_decap_8 FILLER_12_1597 ();
 sg13g2_decap_8 FILLER_12_1604 ();
 sg13g2_decap_8 FILLER_12_1611 ();
 sg13g2_decap_8 FILLER_12_1618 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_4 FILLER_13_343 ();
 sg13g2_fill_2 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_fill_2 FILLER_13_367 ();
 sg13g2_fill_1 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_fill_2 FILLER_13_403 ();
 sg13g2_fill_1 FILLER_13_405 ();
 sg13g2_fill_1 FILLER_13_519 ();
 sg13g2_fill_1 FILLER_13_549 ();
 sg13g2_decap_8 FILLER_13_559 ();
 sg13g2_decap_4 FILLER_13_595 ();
 sg13g2_fill_2 FILLER_13_604 ();
 sg13g2_decap_8 FILLER_13_610 ();
 sg13g2_decap_8 FILLER_13_621 ();
 sg13g2_decap_8 FILLER_13_628 ();
 sg13g2_decap_8 FILLER_13_635 ();
 sg13g2_decap_8 FILLER_13_642 ();
 sg13g2_decap_8 FILLER_13_715 ();
 sg13g2_fill_2 FILLER_13_722 ();
 sg13g2_fill_1 FILLER_13_724 ();
 sg13g2_decap_8 FILLER_13_746 ();
 sg13g2_decap_8 FILLER_13_753 ();
 sg13g2_decap_8 FILLER_13_760 ();
 sg13g2_decap_8 FILLER_13_767 ();
 sg13g2_fill_1 FILLER_13_774 ();
 sg13g2_fill_2 FILLER_13_857 ();
 sg13g2_fill_1 FILLER_13_859 ();
 sg13g2_fill_2 FILLER_13_864 ();
 sg13g2_fill_1 FILLER_13_866 ();
 sg13g2_fill_1 FILLER_13_888 ();
 sg13g2_fill_1 FILLER_13_915 ();
 sg13g2_fill_1 FILLER_13_921 ();
 sg13g2_fill_2 FILLER_13_935 ();
 sg13g2_decap_8 FILLER_13_958 ();
 sg13g2_decap_8 FILLER_13_965 ();
 sg13g2_decap_8 FILLER_13_972 ();
 sg13g2_decap_8 FILLER_13_979 ();
 sg13g2_decap_8 FILLER_13_990 ();
 sg13g2_decap_8 FILLER_13_997 ();
 sg13g2_decap_4 FILLER_13_1004 ();
 sg13g2_decap_8 FILLER_13_1029 ();
 sg13g2_decap_8 FILLER_13_1036 ();
 sg13g2_decap_8 FILLER_13_1047 ();
 sg13g2_fill_2 FILLER_13_1054 ();
 sg13g2_fill_1 FILLER_13_1056 ();
 sg13g2_fill_2 FILLER_13_1066 ();
 sg13g2_fill_1 FILLER_13_1068 ();
 sg13g2_fill_2 FILLER_13_1101 ();
 sg13g2_fill_1 FILLER_13_1103 ();
 sg13g2_fill_2 FILLER_13_1134 ();
 sg13g2_decap_8 FILLER_13_1140 ();
 sg13g2_decap_8 FILLER_13_1147 ();
 sg13g2_decap_8 FILLER_13_1154 ();
 sg13g2_fill_1 FILLER_13_1174 ();
 sg13g2_decap_8 FILLER_13_1211 ();
 sg13g2_decap_8 FILLER_13_1218 ();
 sg13g2_decap_4 FILLER_13_1225 ();
 sg13g2_fill_1 FILLER_13_1229 ();
 sg13g2_decap_8 FILLER_13_1234 ();
 sg13g2_decap_8 FILLER_13_1241 ();
 sg13g2_decap_8 FILLER_13_1248 ();
 sg13g2_decap_8 FILLER_13_1255 ();
 sg13g2_decap_8 FILLER_13_1262 ();
 sg13g2_decap_8 FILLER_13_1269 ();
 sg13g2_decap_8 FILLER_13_1276 ();
 sg13g2_decap_8 FILLER_13_1283 ();
 sg13g2_decap_8 FILLER_13_1290 ();
 sg13g2_decap_8 FILLER_13_1297 ();
 sg13g2_decap_8 FILLER_13_1304 ();
 sg13g2_decap_8 FILLER_13_1311 ();
 sg13g2_decap_8 FILLER_13_1318 ();
 sg13g2_decap_8 FILLER_13_1325 ();
 sg13g2_decap_8 FILLER_13_1332 ();
 sg13g2_decap_8 FILLER_13_1339 ();
 sg13g2_decap_8 FILLER_13_1346 ();
 sg13g2_decap_8 FILLER_13_1353 ();
 sg13g2_decap_8 FILLER_13_1360 ();
 sg13g2_decap_8 FILLER_13_1367 ();
 sg13g2_decap_8 FILLER_13_1374 ();
 sg13g2_decap_8 FILLER_13_1381 ();
 sg13g2_decap_8 FILLER_13_1388 ();
 sg13g2_decap_8 FILLER_13_1395 ();
 sg13g2_decap_8 FILLER_13_1402 ();
 sg13g2_decap_8 FILLER_13_1409 ();
 sg13g2_decap_8 FILLER_13_1416 ();
 sg13g2_decap_8 FILLER_13_1423 ();
 sg13g2_decap_8 FILLER_13_1430 ();
 sg13g2_decap_8 FILLER_13_1437 ();
 sg13g2_decap_8 FILLER_13_1444 ();
 sg13g2_decap_8 FILLER_13_1451 ();
 sg13g2_decap_8 FILLER_13_1458 ();
 sg13g2_decap_8 FILLER_13_1465 ();
 sg13g2_decap_8 FILLER_13_1472 ();
 sg13g2_decap_8 FILLER_13_1479 ();
 sg13g2_decap_8 FILLER_13_1486 ();
 sg13g2_decap_8 FILLER_13_1493 ();
 sg13g2_decap_8 FILLER_13_1500 ();
 sg13g2_decap_8 FILLER_13_1507 ();
 sg13g2_decap_8 FILLER_13_1514 ();
 sg13g2_decap_8 FILLER_13_1521 ();
 sg13g2_decap_8 FILLER_13_1528 ();
 sg13g2_decap_8 FILLER_13_1535 ();
 sg13g2_decap_8 FILLER_13_1542 ();
 sg13g2_decap_8 FILLER_13_1549 ();
 sg13g2_decap_8 FILLER_13_1556 ();
 sg13g2_decap_8 FILLER_13_1563 ();
 sg13g2_decap_8 FILLER_13_1570 ();
 sg13g2_decap_8 FILLER_13_1577 ();
 sg13g2_decap_8 FILLER_13_1584 ();
 sg13g2_decap_8 FILLER_13_1591 ();
 sg13g2_decap_8 FILLER_13_1598 ();
 sg13g2_decap_8 FILLER_13_1605 ();
 sg13g2_decap_8 FILLER_13_1612 ();
 sg13g2_decap_4 FILLER_13_1619 ();
 sg13g2_fill_2 FILLER_13_1623 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_fill_2 FILLER_14_364 ();
 sg13g2_fill_1 FILLER_14_375 ();
 sg13g2_fill_2 FILLER_14_380 ();
 sg13g2_fill_2 FILLER_14_392 ();
 sg13g2_fill_1 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_446 ();
 sg13g2_decap_4 FILLER_14_453 ();
 sg13g2_fill_2 FILLER_14_457 ();
 sg13g2_fill_2 FILLER_14_480 ();
 sg13g2_fill_1 FILLER_14_482 ();
 sg13g2_fill_2 FILLER_14_504 ();
 sg13g2_fill_1 FILLER_14_506 ();
 sg13g2_fill_2 FILLER_14_533 ();
 sg13g2_decap_8 FILLER_14_561 ();
 sg13g2_fill_1 FILLER_14_568 ();
 sg13g2_fill_1 FILLER_14_594 ();
 sg13g2_fill_2 FILLER_14_661 ();
 sg13g2_fill_1 FILLER_14_663 ();
 sg13g2_decap_8 FILLER_14_668 ();
 sg13g2_decap_8 FILLER_14_675 ();
 sg13g2_decap_8 FILLER_14_682 ();
 sg13g2_decap_8 FILLER_14_689 ();
 sg13g2_decap_8 FILLER_14_696 ();
 sg13g2_decap_8 FILLER_14_703 ();
 sg13g2_decap_8 FILLER_14_719 ();
 sg13g2_decap_8 FILLER_14_726 ();
 sg13g2_decap_8 FILLER_14_733 ();
 sg13g2_decap_4 FILLER_14_740 ();
 sg13g2_fill_2 FILLER_14_744 ();
 sg13g2_decap_4 FILLER_14_767 ();
 sg13g2_fill_1 FILLER_14_771 ();
 sg13g2_decap_8 FILLER_14_797 ();
 sg13g2_decap_8 FILLER_14_804 ();
 sg13g2_fill_2 FILLER_14_811 ();
 sg13g2_decap_8 FILLER_14_869 ();
 sg13g2_decap_8 FILLER_14_876 ();
 sg13g2_decap_4 FILLER_14_883 ();
 sg13g2_fill_2 FILLER_14_887 ();
 sg13g2_decap_8 FILLER_14_893 ();
 sg13g2_decap_8 FILLER_14_900 ();
 sg13g2_decap_8 FILLER_14_907 ();
 sg13g2_fill_2 FILLER_14_914 ();
 sg13g2_fill_1 FILLER_14_916 ();
 sg13g2_decap_4 FILLER_14_943 ();
 sg13g2_fill_1 FILLER_14_947 ();
 sg13g2_decap_8 FILLER_14_973 ();
 sg13g2_fill_1 FILLER_14_980 ();
 sg13g2_decap_4 FILLER_14_986 ();
 sg13g2_fill_1 FILLER_14_995 ();
 sg13g2_decap_8 FILLER_14_1004 ();
 sg13g2_decap_8 FILLER_14_1011 ();
 sg13g2_decap_8 FILLER_14_1018 ();
 sg13g2_decap_8 FILLER_14_1025 ();
 sg13g2_fill_2 FILLER_14_1032 ();
 sg13g2_fill_2 FILLER_14_1065 ();
 sg13g2_decap_4 FILLER_14_1102 ();
 sg13g2_decap_8 FILLER_14_1120 ();
 sg13g2_fill_1 FILLER_14_1153 ();
 sg13g2_fill_2 FILLER_14_1210 ();
 sg13g2_decap_8 FILLER_14_1247 ();
 sg13g2_decap_8 FILLER_14_1254 ();
 sg13g2_decap_8 FILLER_14_1261 ();
 sg13g2_decap_8 FILLER_14_1268 ();
 sg13g2_decap_8 FILLER_14_1275 ();
 sg13g2_decap_8 FILLER_14_1282 ();
 sg13g2_decap_8 FILLER_14_1289 ();
 sg13g2_decap_8 FILLER_14_1296 ();
 sg13g2_decap_8 FILLER_14_1303 ();
 sg13g2_decap_8 FILLER_14_1310 ();
 sg13g2_decap_8 FILLER_14_1317 ();
 sg13g2_decap_8 FILLER_14_1324 ();
 sg13g2_decap_8 FILLER_14_1331 ();
 sg13g2_decap_8 FILLER_14_1338 ();
 sg13g2_decap_8 FILLER_14_1345 ();
 sg13g2_decap_8 FILLER_14_1352 ();
 sg13g2_decap_8 FILLER_14_1359 ();
 sg13g2_decap_8 FILLER_14_1366 ();
 sg13g2_decap_8 FILLER_14_1373 ();
 sg13g2_decap_8 FILLER_14_1380 ();
 sg13g2_decap_8 FILLER_14_1387 ();
 sg13g2_decap_8 FILLER_14_1394 ();
 sg13g2_decap_8 FILLER_14_1401 ();
 sg13g2_decap_8 FILLER_14_1408 ();
 sg13g2_decap_8 FILLER_14_1415 ();
 sg13g2_decap_8 FILLER_14_1422 ();
 sg13g2_decap_8 FILLER_14_1429 ();
 sg13g2_decap_8 FILLER_14_1436 ();
 sg13g2_decap_8 FILLER_14_1443 ();
 sg13g2_decap_8 FILLER_14_1450 ();
 sg13g2_decap_8 FILLER_14_1457 ();
 sg13g2_decap_8 FILLER_14_1464 ();
 sg13g2_decap_8 FILLER_14_1471 ();
 sg13g2_decap_8 FILLER_14_1478 ();
 sg13g2_decap_8 FILLER_14_1485 ();
 sg13g2_decap_8 FILLER_14_1492 ();
 sg13g2_decap_8 FILLER_14_1499 ();
 sg13g2_decap_8 FILLER_14_1506 ();
 sg13g2_decap_8 FILLER_14_1513 ();
 sg13g2_decap_8 FILLER_14_1520 ();
 sg13g2_decap_8 FILLER_14_1527 ();
 sg13g2_decap_8 FILLER_14_1534 ();
 sg13g2_decap_8 FILLER_14_1541 ();
 sg13g2_decap_8 FILLER_14_1548 ();
 sg13g2_decap_8 FILLER_14_1555 ();
 sg13g2_decap_8 FILLER_14_1562 ();
 sg13g2_decap_8 FILLER_14_1569 ();
 sg13g2_decap_8 FILLER_14_1576 ();
 sg13g2_decap_8 FILLER_14_1583 ();
 sg13g2_decap_8 FILLER_14_1590 ();
 sg13g2_decap_8 FILLER_14_1597 ();
 sg13g2_decap_8 FILLER_14_1604 ();
 sg13g2_decap_8 FILLER_14_1611 ();
 sg13g2_decap_8 FILLER_14_1618 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_fill_2 FILLER_15_394 ();
 sg13g2_fill_1 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_418 ();
 sg13g2_fill_1 FILLER_15_422 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_4 FILLER_15_525 ();
 sg13g2_fill_1 FILLER_15_529 ();
 sg13g2_decap_4 FILLER_15_534 ();
 sg13g2_fill_1 FILLER_15_567 ();
 sg13g2_fill_1 FILLER_15_589 ();
 sg13g2_decap_4 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_673 ();
 sg13g2_decap_8 FILLER_15_680 ();
 sg13g2_fill_1 FILLER_15_687 ();
 sg13g2_decap_4 FILLER_15_693 ();
 sg13g2_fill_1 FILLER_15_697 ();
 sg13g2_decap_8 FILLER_15_733 ();
 sg13g2_decap_8 FILLER_15_740 ();
 sg13g2_decap_8 FILLER_15_747 ();
 sg13g2_decap_8 FILLER_15_754 ();
 sg13g2_decap_8 FILLER_15_761 ();
 sg13g2_fill_2 FILLER_15_777 ();
 sg13g2_fill_2 FILLER_15_784 ();
 sg13g2_fill_1 FILLER_15_786 ();
 sg13g2_decap_8 FILLER_15_808 ();
 sg13g2_decap_4 FILLER_15_815 ();
 sg13g2_fill_1 FILLER_15_819 ();
 sg13g2_decap_4 FILLER_15_834 ();
 sg13g2_fill_2 FILLER_15_838 ();
 sg13g2_decap_4 FILLER_15_844 ();
 sg13g2_fill_2 FILLER_15_848 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_decap_8 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_15_868 ();
 sg13g2_decap_8 FILLER_15_875 ();
 sg13g2_fill_1 FILLER_15_882 ();
 sg13g2_decap_8 FILLER_15_888 ();
 sg13g2_decap_8 FILLER_15_895 ();
 sg13g2_decap_4 FILLER_15_902 ();
 sg13g2_fill_1 FILLER_15_906 ();
 sg13g2_fill_2 FILLER_15_958 ();
 sg13g2_fill_1 FILLER_15_986 ();
 sg13g2_decap_4 FILLER_15_1017 ();
 sg13g2_decap_8 FILLER_15_1046 ();
 sg13g2_decap_8 FILLER_15_1053 ();
 sg13g2_decap_8 FILLER_15_1060 ();
 sg13g2_decap_8 FILLER_15_1067 ();
 sg13g2_decap_8 FILLER_15_1074 ();
 sg13g2_decap_8 FILLER_15_1081 ();
 sg13g2_decap_8 FILLER_15_1088 ();
 sg13g2_decap_8 FILLER_15_1095 ();
 sg13g2_decap_4 FILLER_15_1102 ();
 sg13g2_fill_1 FILLER_15_1106 ();
 sg13g2_decap_4 FILLER_15_1111 ();
 sg13g2_fill_1 FILLER_15_1115 ();
 sg13g2_decap_8 FILLER_15_1137 ();
 sg13g2_decap_4 FILLER_15_1144 ();
 sg13g2_fill_1 FILLER_15_1148 ();
 sg13g2_decap_8 FILLER_15_1154 ();
 sg13g2_fill_2 FILLER_15_1161 ();
 sg13g2_fill_2 FILLER_15_1188 ();
 sg13g2_fill_1 FILLER_15_1190 ();
 sg13g2_decap_8 FILLER_15_1217 ();
 sg13g2_decap_8 FILLER_15_1224 ();
 sg13g2_decap_8 FILLER_15_1235 ();
 sg13g2_decap_8 FILLER_15_1242 ();
 sg13g2_decap_8 FILLER_15_1249 ();
 sg13g2_decap_8 FILLER_15_1256 ();
 sg13g2_decap_8 FILLER_15_1263 ();
 sg13g2_decap_8 FILLER_15_1270 ();
 sg13g2_decap_8 FILLER_15_1277 ();
 sg13g2_decap_8 FILLER_15_1284 ();
 sg13g2_decap_8 FILLER_15_1291 ();
 sg13g2_decap_8 FILLER_15_1298 ();
 sg13g2_decap_8 FILLER_15_1305 ();
 sg13g2_decap_8 FILLER_15_1312 ();
 sg13g2_decap_8 FILLER_15_1319 ();
 sg13g2_decap_8 FILLER_15_1326 ();
 sg13g2_decap_8 FILLER_15_1333 ();
 sg13g2_decap_8 FILLER_15_1340 ();
 sg13g2_decap_8 FILLER_15_1347 ();
 sg13g2_decap_8 FILLER_15_1354 ();
 sg13g2_decap_8 FILLER_15_1361 ();
 sg13g2_decap_8 FILLER_15_1368 ();
 sg13g2_decap_8 FILLER_15_1375 ();
 sg13g2_decap_8 FILLER_15_1382 ();
 sg13g2_decap_8 FILLER_15_1389 ();
 sg13g2_decap_8 FILLER_15_1396 ();
 sg13g2_decap_8 FILLER_15_1403 ();
 sg13g2_decap_8 FILLER_15_1410 ();
 sg13g2_decap_8 FILLER_15_1417 ();
 sg13g2_decap_8 FILLER_15_1424 ();
 sg13g2_decap_8 FILLER_15_1431 ();
 sg13g2_decap_8 FILLER_15_1438 ();
 sg13g2_decap_8 FILLER_15_1445 ();
 sg13g2_decap_8 FILLER_15_1452 ();
 sg13g2_decap_8 FILLER_15_1459 ();
 sg13g2_decap_8 FILLER_15_1466 ();
 sg13g2_decap_8 FILLER_15_1473 ();
 sg13g2_decap_8 FILLER_15_1480 ();
 sg13g2_decap_8 FILLER_15_1487 ();
 sg13g2_decap_8 FILLER_15_1494 ();
 sg13g2_decap_8 FILLER_15_1501 ();
 sg13g2_decap_8 FILLER_15_1508 ();
 sg13g2_decap_8 FILLER_15_1515 ();
 sg13g2_decap_8 FILLER_15_1522 ();
 sg13g2_decap_8 FILLER_15_1529 ();
 sg13g2_decap_8 FILLER_15_1536 ();
 sg13g2_decap_8 FILLER_15_1543 ();
 sg13g2_decap_8 FILLER_15_1550 ();
 sg13g2_decap_8 FILLER_15_1557 ();
 sg13g2_decap_8 FILLER_15_1564 ();
 sg13g2_decap_8 FILLER_15_1571 ();
 sg13g2_decap_8 FILLER_15_1578 ();
 sg13g2_decap_8 FILLER_15_1585 ();
 sg13g2_decap_8 FILLER_15_1592 ();
 sg13g2_decap_8 FILLER_15_1599 ();
 sg13g2_decap_8 FILLER_15_1606 ();
 sg13g2_decap_8 FILLER_15_1613 ();
 sg13g2_decap_4 FILLER_15_1620 ();
 sg13g2_fill_1 FILLER_15_1624 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_4 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_fill_2 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_355 ();
 sg13g2_fill_2 FILLER_16_381 ();
 sg13g2_fill_2 FILLER_16_409 ();
 sg13g2_fill_1 FILLER_16_411 ();
 sg13g2_fill_2 FILLER_16_421 ();
 sg13g2_fill_1 FILLER_16_423 ();
 sg13g2_decap_8 FILLER_16_459 ();
 sg13g2_decap_4 FILLER_16_466 ();
 sg13g2_decap_8 FILLER_16_474 ();
 sg13g2_decap_4 FILLER_16_507 ();
 sg13g2_fill_2 FILLER_16_511 ();
 sg13g2_fill_1 FILLER_16_523 ();
 sg13g2_fill_1 FILLER_16_528 ();
 sg13g2_fill_1 FILLER_16_581 ();
 sg13g2_fill_2 FILLER_16_592 ();
 sg13g2_fill_1 FILLER_16_594 ();
 sg13g2_fill_2 FILLER_16_600 ();
 sg13g2_decap_8 FILLER_16_636 ();
 sg13g2_fill_2 FILLER_16_643 ();
 sg13g2_fill_1 FILLER_16_645 ();
 sg13g2_fill_2 FILLER_16_681 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_730 ();
 sg13g2_decap_8 FILLER_16_794 ();
 sg13g2_decap_4 FILLER_16_801 ();
 sg13g2_decap_4 FILLER_16_831 ();
 sg13g2_fill_1 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_841 ();
 sg13g2_decap_4 FILLER_16_848 ();
 sg13g2_fill_1 FILLER_16_852 ();
 sg13g2_decap_4 FILLER_16_857 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_16_904 ();
 sg13g2_decap_8 FILLER_16_911 ();
 sg13g2_fill_1 FILLER_16_918 ();
 sg13g2_decap_8 FILLER_16_953 ();
 sg13g2_decap_4 FILLER_16_960 ();
 sg13g2_fill_1 FILLER_16_964 ();
 sg13g2_fill_1 FILLER_16_979 ();
 sg13g2_decap_8 FILLER_16_1026 ();
 sg13g2_fill_1 FILLER_16_1033 ();
 sg13g2_fill_2 FILLER_16_1081 ();
 sg13g2_fill_1 FILLER_16_1083 ();
 sg13g2_decap_8 FILLER_16_1088 ();
 sg13g2_decap_8 FILLER_16_1099 ();
 sg13g2_decap_8 FILLER_16_1106 ();
 sg13g2_fill_2 FILLER_16_1113 ();
 sg13g2_decap_4 FILLER_16_1136 ();
 sg13g2_fill_1 FILLER_16_1169 ();
 sg13g2_fill_2 FILLER_16_1200 ();
 sg13g2_fill_1 FILLER_16_1202 ();
 sg13g2_decap_8 FILLER_16_1207 ();
 sg13g2_fill_1 FILLER_16_1214 ();
 sg13g2_fill_1 FILLER_16_1224 ();
 sg13g2_decap_8 FILLER_16_1255 ();
 sg13g2_decap_8 FILLER_16_1262 ();
 sg13g2_decap_8 FILLER_16_1269 ();
 sg13g2_decap_8 FILLER_16_1276 ();
 sg13g2_decap_8 FILLER_16_1283 ();
 sg13g2_decap_8 FILLER_16_1290 ();
 sg13g2_decap_8 FILLER_16_1297 ();
 sg13g2_decap_8 FILLER_16_1304 ();
 sg13g2_decap_8 FILLER_16_1311 ();
 sg13g2_decap_8 FILLER_16_1318 ();
 sg13g2_decap_8 FILLER_16_1325 ();
 sg13g2_decap_8 FILLER_16_1332 ();
 sg13g2_decap_8 FILLER_16_1339 ();
 sg13g2_decap_8 FILLER_16_1346 ();
 sg13g2_decap_8 FILLER_16_1353 ();
 sg13g2_decap_8 FILLER_16_1360 ();
 sg13g2_decap_8 FILLER_16_1367 ();
 sg13g2_decap_8 FILLER_16_1374 ();
 sg13g2_decap_8 FILLER_16_1381 ();
 sg13g2_decap_8 FILLER_16_1388 ();
 sg13g2_decap_8 FILLER_16_1395 ();
 sg13g2_decap_8 FILLER_16_1402 ();
 sg13g2_decap_8 FILLER_16_1409 ();
 sg13g2_decap_8 FILLER_16_1416 ();
 sg13g2_decap_8 FILLER_16_1423 ();
 sg13g2_decap_8 FILLER_16_1430 ();
 sg13g2_decap_8 FILLER_16_1437 ();
 sg13g2_decap_8 FILLER_16_1444 ();
 sg13g2_decap_8 FILLER_16_1451 ();
 sg13g2_decap_8 FILLER_16_1458 ();
 sg13g2_decap_8 FILLER_16_1465 ();
 sg13g2_decap_8 FILLER_16_1472 ();
 sg13g2_decap_8 FILLER_16_1479 ();
 sg13g2_decap_8 FILLER_16_1486 ();
 sg13g2_decap_8 FILLER_16_1493 ();
 sg13g2_decap_8 FILLER_16_1500 ();
 sg13g2_decap_8 FILLER_16_1507 ();
 sg13g2_decap_8 FILLER_16_1514 ();
 sg13g2_decap_8 FILLER_16_1521 ();
 sg13g2_decap_8 FILLER_16_1528 ();
 sg13g2_decap_8 FILLER_16_1535 ();
 sg13g2_decap_8 FILLER_16_1542 ();
 sg13g2_decap_8 FILLER_16_1549 ();
 sg13g2_decap_8 FILLER_16_1556 ();
 sg13g2_decap_8 FILLER_16_1563 ();
 sg13g2_decap_8 FILLER_16_1570 ();
 sg13g2_decap_8 FILLER_16_1577 ();
 sg13g2_decap_8 FILLER_16_1584 ();
 sg13g2_decap_8 FILLER_16_1591 ();
 sg13g2_decap_8 FILLER_16_1598 ();
 sg13g2_decap_8 FILLER_16_1605 ();
 sg13g2_decap_8 FILLER_16_1612 ();
 sg13g2_decap_4 FILLER_16_1619 ();
 sg13g2_fill_2 FILLER_16_1623 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_4 FILLER_17_315 ();
 sg13g2_fill_1 FILLER_17_319 ();
 sg13g2_fill_1 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_fill_1 FILLER_17_435 ();
 sg13g2_fill_1 FILLER_17_462 ();
 sg13g2_decap_4 FILLER_17_489 ();
 sg13g2_fill_2 FILLER_17_493 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_fill_1 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_538 ();
 sg13g2_decap_4 FILLER_17_545 ();
 sg13g2_fill_2 FILLER_17_549 ();
 sg13g2_decap_8 FILLER_17_631 ();
 sg13g2_decap_8 FILLER_17_643 ();
 sg13g2_decap_4 FILLER_17_650 ();
 sg13g2_fill_1 FILLER_17_654 ();
 sg13g2_decap_8 FILLER_17_660 ();
 sg13g2_decap_8 FILLER_17_667 ();
 sg13g2_decap_8 FILLER_17_674 ();
 sg13g2_decap_8 FILLER_17_681 ();
 sg13g2_fill_2 FILLER_17_688 ();
 sg13g2_fill_2 FILLER_17_698 ();
 sg13g2_fill_2 FILLER_17_729 ();
 sg13g2_fill_1 FILLER_17_731 ();
 sg13g2_decap_8 FILLER_17_753 ();
 sg13g2_decap_8 FILLER_17_760 ();
 sg13g2_decap_8 FILLER_17_767 ();
 sg13g2_fill_1 FILLER_17_774 ();
 sg13g2_decap_8 FILLER_17_800 ();
 sg13g2_decap_4 FILLER_17_807 ();
 sg13g2_fill_1 FILLER_17_811 ();
 sg13g2_decap_8 FILLER_17_816 ();
 sg13g2_fill_1 FILLER_17_823 ();
 sg13g2_fill_2 FILLER_17_859 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_fill_2 FILLER_17_883 ();
 sg13g2_fill_2 FILLER_17_906 ();
 sg13g2_fill_1 FILLER_17_908 ();
 sg13g2_decap_8 FILLER_17_935 ();
 sg13g2_decap_4 FILLER_17_942 ();
 sg13g2_fill_1 FILLER_17_946 ();
 sg13g2_decap_8 FILLER_17_968 ();
 sg13g2_fill_1 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1023 ();
 sg13g2_fill_2 FILLER_17_1030 ();
 sg13g2_fill_1 FILLER_17_1032 ();
 sg13g2_decap_4 FILLER_17_1038 ();
 sg13g2_fill_1 FILLER_17_1042 ();
 sg13g2_decap_4 FILLER_17_1046 ();
 sg13g2_fill_1 FILLER_17_1050 ();
 sg13g2_decap_4 FILLER_17_1080 ();
 sg13g2_decap_8 FILLER_17_1136 ();
 sg13g2_fill_1 FILLER_17_1143 ();
 sg13g2_decap_8 FILLER_17_1170 ();
 sg13g2_fill_2 FILLER_17_1177 ();
 sg13g2_decap_4 FILLER_17_1208 ();
 sg13g2_decap_4 FILLER_17_1233 ();
 sg13g2_fill_1 FILLER_17_1237 ();
 sg13g2_decap_8 FILLER_17_1263 ();
 sg13g2_decap_8 FILLER_17_1270 ();
 sg13g2_decap_8 FILLER_17_1277 ();
 sg13g2_decap_8 FILLER_17_1284 ();
 sg13g2_decap_8 FILLER_17_1291 ();
 sg13g2_decap_8 FILLER_17_1298 ();
 sg13g2_decap_8 FILLER_17_1305 ();
 sg13g2_decap_8 FILLER_17_1312 ();
 sg13g2_decap_8 FILLER_17_1319 ();
 sg13g2_decap_8 FILLER_17_1326 ();
 sg13g2_decap_8 FILLER_17_1333 ();
 sg13g2_decap_8 FILLER_17_1340 ();
 sg13g2_decap_8 FILLER_17_1347 ();
 sg13g2_decap_8 FILLER_17_1354 ();
 sg13g2_decap_8 FILLER_17_1361 ();
 sg13g2_decap_8 FILLER_17_1368 ();
 sg13g2_decap_8 FILLER_17_1375 ();
 sg13g2_decap_8 FILLER_17_1382 ();
 sg13g2_decap_8 FILLER_17_1389 ();
 sg13g2_decap_8 FILLER_17_1396 ();
 sg13g2_decap_8 FILLER_17_1403 ();
 sg13g2_decap_8 FILLER_17_1410 ();
 sg13g2_decap_8 FILLER_17_1417 ();
 sg13g2_decap_8 FILLER_17_1424 ();
 sg13g2_decap_8 FILLER_17_1431 ();
 sg13g2_decap_8 FILLER_17_1438 ();
 sg13g2_decap_8 FILLER_17_1445 ();
 sg13g2_decap_8 FILLER_17_1452 ();
 sg13g2_decap_8 FILLER_17_1459 ();
 sg13g2_decap_8 FILLER_17_1466 ();
 sg13g2_decap_8 FILLER_17_1473 ();
 sg13g2_decap_8 FILLER_17_1480 ();
 sg13g2_decap_8 FILLER_17_1487 ();
 sg13g2_decap_8 FILLER_17_1494 ();
 sg13g2_decap_8 FILLER_17_1501 ();
 sg13g2_decap_8 FILLER_17_1508 ();
 sg13g2_decap_8 FILLER_17_1515 ();
 sg13g2_decap_8 FILLER_17_1522 ();
 sg13g2_decap_8 FILLER_17_1529 ();
 sg13g2_decap_8 FILLER_17_1536 ();
 sg13g2_decap_8 FILLER_17_1543 ();
 sg13g2_decap_8 FILLER_17_1550 ();
 sg13g2_decap_8 FILLER_17_1557 ();
 sg13g2_decap_8 FILLER_17_1564 ();
 sg13g2_decap_8 FILLER_17_1571 ();
 sg13g2_decap_8 FILLER_17_1578 ();
 sg13g2_decap_8 FILLER_17_1585 ();
 sg13g2_decap_8 FILLER_17_1592 ();
 sg13g2_decap_8 FILLER_17_1599 ();
 sg13g2_decap_8 FILLER_17_1606 ();
 sg13g2_decap_8 FILLER_17_1613 ();
 sg13g2_decap_4 FILLER_17_1620 ();
 sg13g2_fill_1 FILLER_17_1624 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_4 FILLER_18_329 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_decap_4 FILLER_18_338 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_fill_2 FILLER_18_361 ();
 sg13g2_fill_2 FILLER_18_403 ();
 sg13g2_decap_8 FILLER_18_409 ();
 sg13g2_decap_8 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_452 ();
 sg13g2_decap_8 FILLER_18_459 ();
 sg13g2_fill_2 FILLER_18_466 ();
 sg13g2_fill_2 FILLER_18_523 ();
 sg13g2_decap_8 FILLER_18_551 ();
 sg13g2_decap_8 FILLER_18_558 ();
 sg13g2_fill_1 FILLER_18_565 ();
 sg13g2_decap_8 FILLER_18_641 ();
 sg13g2_fill_1 FILLER_18_648 ();
 sg13g2_decap_4 FILLER_18_670 ();
 sg13g2_fill_2 FILLER_18_678 ();
 sg13g2_fill_1 FILLER_18_685 ();
 sg13g2_decap_8 FILLER_18_690 ();
 sg13g2_decap_8 FILLER_18_697 ();
 sg13g2_decap_8 FILLER_18_704 ();
 sg13g2_decap_4 FILLER_18_737 ();
 sg13g2_fill_2 FILLER_18_741 ();
 sg13g2_decap_4 FILLER_18_774 ();
 sg13g2_fill_1 FILLER_18_778 ();
 sg13g2_fill_2 FILLER_18_800 ();
 sg13g2_fill_1 FILLER_18_802 ();
 sg13g2_decap_4 FILLER_18_807 ();
 sg13g2_fill_1 FILLER_18_811 ();
 sg13g2_decap_8 FILLER_18_873 ();
 sg13g2_fill_2 FILLER_18_880 ();
 sg13g2_decap_8 FILLER_18_887 ();
 sg13g2_decap_8 FILLER_18_894 ();
 sg13g2_decap_8 FILLER_18_901 ();
 sg13g2_decap_8 FILLER_18_908 ();
 sg13g2_fill_2 FILLER_18_919 ();
 sg13g2_decap_8 FILLER_18_929 ();
 sg13g2_decap_8 FILLER_18_936 ();
 sg13g2_decap_4 FILLER_18_943 ();
 sg13g2_fill_1 FILLER_18_947 ();
 sg13g2_decap_8 FILLER_18_956 ();
 sg13g2_decap_8 FILLER_18_963 ();
 sg13g2_decap_8 FILLER_18_970 ();
 sg13g2_fill_1 FILLER_18_977 ();
 sg13g2_decap_4 FILLER_18_985 ();
 sg13g2_decap_8 FILLER_18_994 ();
 sg13g2_decap_8 FILLER_18_1001 ();
 sg13g2_decap_8 FILLER_18_1008 ();
 sg13g2_decap_8 FILLER_18_1015 ();
 sg13g2_decap_8 FILLER_18_1022 ();
 sg13g2_decap_8 FILLER_18_1029 ();
 sg13g2_fill_2 FILLER_18_1036 ();
 sg13g2_fill_2 FILLER_18_1068 ();
 sg13g2_fill_1 FILLER_18_1070 ();
 sg13g2_fill_1 FILLER_18_1092 ();
 sg13g2_fill_2 FILLER_18_1098 ();
 sg13g2_fill_1 FILLER_18_1100 ();
 sg13g2_decap_8 FILLER_18_1126 ();
 sg13g2_decap_8 FILLER_18_1133 ();
 sg13g2_decap_8 FILLER_18_1140 ();
 sg13g2_decap_4 FILLER_18_1147 ();
 sg13g2_decap_8 FILLER_18_1155 ();
 sg13g2_decap_8 FILLER_18_1162 ();
 sg13g2_decap_8 FILLER_18_1169 ();
 sg13g2_decap_8 FILLER_18_1176 ();
 sg13g2_decap_8 FILLER_18_1183 ();
 sg13g2_fill_1 FILLER_18_1216 ();
 sg13g2_fill_2 FILLER_18_1238 ();
 sg13g2_fill_1 FILLER_18_1240 ();
 sg13g2_decap_8 FILLER_18_1267 ();
 sg13g2_decap_8 FILLER_18_1274 ();
 sg13g2_decap_8 FILLER_18_1281 ();
 sg13g2_decap_8 FILLER_18_1288 ();
 sg13g2_decap_8 FILLER_18_1295 ();
 sg13g2_decap_8 FILLER_18_1302 ();
 sg13g2_decap_8 FILLER_18_1309 ();
 sg13g2_decap_8 FILLER_18_1316 ();
 sg13g2_decap_8 FILLER_18_1323 ();
 sg13g2_decap_8 FILLER_18_1330 ();
 sg13g2_decap_8 FILLER_18_1337 ();
 sg13g2_decap_8 FILLER_18_1344 ();
 sg13g2_decap_8 FILLER_18_1351 ();
 sg13g2_decap_8 FILLER_18_1358 ();
 sg13g2_decap_8 FILLER_18_1365 ();
 sg13g2_decap_8 FILLER_18_1372 ();
 sg13g2_decap_8 FILLER_18_1379 ();
 sg13g2_decap_8 FILLER_18_1386 ();
 sg13g2_decap_8 FILLER_18_1393 ();
 sg13g2_decap_8 FILLER_18_1400 ();
 sg13g2_decap_8 FILLER_18_1407 ();
 sg13g2_decap_8 FILLER_18_1414 ();
 sg13g2_decap_8 FILLER_18_1421 ();
 sg13g2_decap_8 FILLER_18_1428 ();
 sg13g2_decap_8 FILLER_18_1435 ();
 sg13g2_decap_8 FILLER_18_1442 ();
 sg13g2_decap_8 FILLER_18_1449 ();
 sg13g2_decap_8 FILLER_18_1456 ();
 sg13g2_decap_8 FILLER_18_1463 ();
 sg13g2_decap_8 FILLER_18_1470 ();
 sg13g2_decap_8 FILLER_18_1477 ();
 sg13g2_decap_8 FILLER_18_1484 ();
 sg13g2_decap_8 FILLER_18_1491 ();
 sg13g2_decap_8 FILLER_18_1498 ();
 sg13g2_decap_8 FILLER_18_1505 ();
 sg13g2_decap_8 FILLER_18_1512 ();
 sg13g2_decap_8 FILLER_18_1519 ();
 sg13g2_decap_8 FILLER_18_1526 ();
 sg13g2_decap_8 FILLER_18_1533 ();
 sg13g2_decap_8 FILLER_18_1540 ();
 sg13g2_decap_8 FILLER_18_1547 ();
 sg13g2_decap_8 FILLER_18_1554 ();
 sg13g2_decap_8 FILLER_18_1561 ();
 sg13g2_decap_8 FILLER_18_1568 ();
 sg13g2_decap_8 FILLER_18_1575 ();
 sg13g2_decap_8 FILLER_18_1582 ();
 sg13g2_decap_8 FILLER_18_1589 ();
 sg13g2_decap_8 FILLER_18_1596 ();
 sg13g2_decap_8 FILLER_18_1603 ();
 sg13g2_decap_8 FILLER_18_1610 ();
 sg13g2_decap_8 FILLER_18_1617 ();
 sg13g2_fill_1 FILLER_18_1624 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_fill_2 FILLER_19_322 ();
 sg13g2_fill_1 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_4 FILLER_19_370 ();
 sg13g2_fill_2 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_4 FILLER_19_387 ();
 sg13g2_fill_1 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_decap_4 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_19_442 ();
 sg13g2_decap_8 FILLER_19_449 ();
 sg13g2_decap_8 FILLER_19_456 ();
 sg13g2_decap_4 FILLER_19_463 ();
 sg13g2_decap_8 FILLER_19_480 ();
 sg13g2_decap_4 FILLER_19_487 ();
 sg13g2_fill_2 FILLER_19_491 ();
 sg13g2_decap_4 FILLER_19_514 ();
 sg13g2_fill_1 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_523 ();
 sg13g2_decap_4 FILLER_19_530 ();
 sg13g2_fill_2 FILLER_19_534 ();
 sg13g2_decap_8 FILLER_19_540 ();
 sg13g2_decap_4 FILLER_19_547 ();
 sg13g2_fill_2 FILLER_19_572 ();
 sg13g2_decap_4 FILLER_19_628 ();
 sg13g2_decap_8 FILLER_19_636 ();
 sg13g2_decap_8 FILLER_19_643 ();
 sg13g2_fill_2 FILLER_19_671 ();
 sg13g2_fill_2 FILLER_19_708 ();
 sg13g2_fill_2 FILLER_19_760 ();
 sg13g2_fill_1 FILLER_19_762 ();
 sg13g2_decap_8 FILLER_19_773 ();
 sg13g2_decap_8 FILLER_19_780 ();
 sg13g2_fill_2 FILLER_19_812 ();
 sg13g2_fill_1 FILLER_19_814 ();
 sg13g2_fill_1 FILLER_19_841 ();
 sg13g2_fill_2 FILLER_19_871 ();
 sg13g2_decap_8 FILLER_19_894 ();
 sg13g2_decap_8 FILLER_19_901 ();
 sg13g2_fill_2 FILLER_19_908 ();
 sg13g2_fill_1 FILLER_19_910 ();
 sg13g2_fill_2 FILLER_19_941 ();
 sg13g2_fill_1 FILLER_19_943 ();
 sg13g2_fill_2 FILLER_19_975 ();
 sg13g2_decap_8 FILLER_19_1010 ();
 sg13g2_decap_8 FILLER_19_1017 ();
 sg13g2_decap_8 FILLER_19_1024 ();
 sg13g2_fill_2 FILLER_19_1031 ();
 sg13g2_decap_4 FILLER_19_1038 ();
 sg13g2_fill_1 FILLER_19_1042 ();
 sg13g2_decap_4 FILLER_19_1140 ();
 sg13g2_fill_2 FILLER_19_1144 ();
 sg13g2_decap_8 FILLER_19_1150 ();
 sg13g2_decap_8 FILLER_19_1157 ();
 sg13g2_fill_2 FILLER_19_1164 ();
 sg13g2_fill_1 FILLER_19_1175 ();
 sg13g2_fill_2 FILLER_19_1213 ();
 sg13g2_fill_1 FILLER_19_1215 ();
 sg13g2_decap_4 FILLER_19_1221 ();
 sg13g2_fill_2 FILLER_19_1225 ();
 sg13g2_decap_8 FILLER_19_1231 ();
 sg13g2_decap_8 FILLER_19_1238 ();
 sg13g2_decap_8 FILLER_19_1245 ();
 sg13g2_fill_1 FILLER_19_1252 ();
 sg13g2_decap_8 FILLER_19_1286 ();
 sg13g2_decap_8 FILLER_19_1293 ();
 sg13g2_decap_8 FILLER_19_1300 ();
 sg13g2_decap_8 FILLER_19_1307 ();
 sg13g2_decap_8 FILLER_19_1314 ();
 sg13g2_decap_8 FILLER_19_1321 ();
 sg13g2_decap_8 FILLER_19_1328 ();
 sg13g2_decap_8 FILLER_19_1335 ();
 sg13g2_decap_8 FILLER_19_1342 ();
 sg13g2_decap_8 FILLER_19_1349 ();
 sg13g2_decap_8 FILLER_19_1356 ();
 sg13g2_decap_8 FILLER_19_1363 ();
 sg13g2_decap_8 FILLER_19_1370 ();
 sg13g2_decap_8 FILLER_19_1377 ();
 sg13g2_decap_8 FILLER_19_1384 ();
 sg13g2_decap_8 FILLER_19_1391 ();
 sg13g2_decap_8 FILLER_19_1398 ();
 sg13g2_decap_8 FILLER_19_1405 ();
 sg13g2_decap_8 FILLER_19_1412 ();
 sg13g2_decap_8 FILLER_19_1419 ();
 sg13g2_decap_8 FILLER_19_1426 ();
 sg13g2_decap_8 FILLER_19_1433 ();
 sg13g2_decap_8 FILLER_19_1440 ();
 sg13g2_decap_8 FILLER_19_1447 ();
 sg13g2_decap_8 FILLER_19_1454 ();
 sg13g2_decap_8 FILLER_19_1461 ();
 sg13g2_decap_8 FILLER_19_1468 ();
 sg13g2_decap_8 FILLER_19_1475 ();
 sg13g2_decap_8 FILLER_19_1482 ();
 sg13g2_decap_8 FILLER_19_1489 ();
 sg13g2_decap_8 FILLER_19_1496 ();
 sg13g2_decap_8 FILLER_19_1503 ();
 sg13g2_decap_8 FILLER_19_1510 ();
 sg13g2_decap_8 FILLER_19_1517 ();
 sg13g2_decap_8 FILLER_19_1524 ();
 sg13g2_decap_8 FILLER_19_1531 ();
 sg13g2_decap_8 FILLER_19_1538 ();
 sg13g2_decap_8 FILLER_19_1545 ();
 sg13g2_decap_8 FILLER_19_1552 ();
 sg13g2_decap_8 FILLER_19_1559 ();
 sg13g2_decap_8 FILLER_19_1566 ();
 sg13g2_decap_8 FILLER_19_1573 ();
 sg13g2_decap_8 FILLER_19_1580 ();
 sg13g2_decap_8 FILLER_19_1587 ();
 sg13g2_decap_8 FILLER_19_1594 ();
 sg13g2_decap_8 FILLER_19_1601 ();
 sg13g2_decap_8 FILLER_19_1608 ();
 sg13g2_decap_8 FILLER_19_1615 ();
 sg13g2_fill_2 FILLER_19_1622 ();
 sg13g2_fill_1 FILLER_19_1624 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_fill_2 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_fill_2 FILLER_20_383 ();
 sg13g2_fill_1 FILLER_20_385 ();
 sg13g2_decap_4 FILLER_20_412 ();
 sg13g2_fill_2 FILLER_20_416 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_fill_2 FILLER_20_456 ();
 sg13g2_fill_2 FILLER_20_484 ();
 sg13g2_fill_1 FILLER_20_486 ();
 sg13g2_decap_8 FILLER_20_491 ();
 sg13g2_decap_8 FILLER_20_498 ();
 sg13g2_decap_8 FILLER_20_505 ();
 sg13g2_decap_8 FILLER_20_512 ();
 sg13g2_fill_1 FILLER_20_519 ();
 sg13g2_decap_8 FILLER_20_524 ();
 sg13g2_decap_8 FILLER_20_531 ();
 sg13g2_decap_8 FILLER_20_538 ();
 sg13g2_fill_2 FILLER_20_545 ();
 sg13g2_fill_1 FILLER_20_547 ();
 sg13g2_decap_8 FILLER_20_552 ();
 sg13g2_decap_8 FILLER_20_559 ();
 sg13g2_decap_8 FILLER_20_566 ();
 sg13g2_fill_2 FILLER_20_573 ();
 sg13g2_fill_1 FILLER_20_575 ();
 sg13g2_decap_4 FILLER_20_633 ();
 sg13g2_fill_2 FILLER_20_637 ();
 sg13g2_decap_4 FILLER_20_643 ();
 sg13g2_decap_8 FILLER_20_652 ();
 sg13g2_decap_8 FILLER_20_659 ();
 sg13g2_decap_8 FILLER_20_666 ();
 sg13g2_fill_2 FILLER_20_673 ();
 sg13g2_fill_1 FILLER_20_675 ();
 sg13g2_fill_2 FILLER_20_705 ();
 sg13g2_fill_1 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_734 ();
 sg13g2_decap_4 FILLER_20_741 ();
 sg13g2_fill_2 FILLER_20_745 ();
 sg13g2_fill_2 FILLER_20_793 ();
 sg13g2_fill_1 FILLER_20_795 ();
 sg13g2_decap_8 FILLER_20_822 ();
 sg13g2_decap_8 FILLER_20_829 ();
 sg13g2_decap_4 FILLER_20_836 ();
 sg13g2_fill_1 FILLER_20_840 ();
 sg13g2_fill_2 FILLER_20_846 ();
 sg13g2_fill_1 FILLER_20_848 ();
 sg13g2_decap_4 FILLER_20_858 ();
 sg13g2_fill_1 FILLER_20_862 ();
 sg13g2_decap_4 FILLER_20_868 ();
 sg13g2_fill_1 FILLER_20_872 ();
 sg13g2_decap_8 FILLER_20_899 ();
 sg13g2_fill_2 FILLER_20_906 ();
 sg13g2_fill_1 FILLER_20_908 ();
 sg13g2_fill_2 FILLER_20_940 ();
 sg13g2_fill_1 FILLER_20_942 ();
 sg13g2_fill_2 FILLER_20_948 ();
 sg13g2_fill_1 FILLER_20_950 ();
 sg13g2_fill_2 FILLER_20_976 ();
 sg13g2_decap_4 FILLER_20_1004 ();
 sg13g2_fill_1 FILLER_20_1008 ();
 sg13g2_decap_8 FILLER_20_1014 ();
 sg13g2_fill_2 FILLER_20_1021 ();
 sg13g2_decap_8 FILLER_20_1044 ();
 sg13g2_decap_8 FILLER_20_1060 ();
 sg13g2_decap_8 FILLER_20_1067 ();
 sg13g2_decap_8 FILLER_20_1074 ();
 sg13g2_decap_4 FILLER_20_1081 ();
 sg13g2_decap_8 FILLER_20_1120 ();
 sg13g2_fill_2 FILLER_20_1127 ();
 sg13g2_decap_4 FILLER_20_1134 ();
 sg13g2_fill_2 FILLER_20_1138 ();
 sg13g2_fill_2 FILLER_20_1166 ();
 sg13g2_fill_1 FILLER_20_1219 ();
 sg13g2_fill_2 FILLER_20_1245 ();
 sg13g2_fill_2 FILLER_20_1273 ();
 sg13g2_decap_8 FILLER_20_1300 ();
 sg13g2_decap_8 FILLER_20_1307 ();
 sg13g2_decap_8 FILLER_20_1314 ();
 sg13g2_decap_8 FILLER_20_1321 ();
 sg13g2_decap_8 FILLER_20_1328 ();
 sg13g2_decap_8 FILLER_20_1335 ();
 sg13g2_decap_8 FILLER_20_1342 ();
 sg13g2_decap_8 FILLER_20_1349 ();
 sg13g2_decap_8 FILLER_20_1356 ();
 sg13g2_decap_8 FILLER_20_1363 ();
 sg13g2_decap_8 FILLER_20_1370 ();
 sg13g2_decap_8 FILLER_20_1377 ();
 sg13g2_decap_8 FILLER_20_1384 ();
 sg13g2_decap_8 FILLER_20_1391 ();
 sg13g2_decap_8 FILLER_20_1398 ();
 sg13g2_decap_8 FILLER_20_1405 ();
 sg13g2_decap_8 FILLER_20_1412 ();
 sg13g2_decap_8 FILLER_20_1419 ();
 sg13g2_decap_8 FILLER_20_1426 ();
 sg13g2_decap_8 FILLER_20_1433 ();
 sg13g2_decap_8 FILLER_20_1440 ();
 sg13g2_decap_8 FILLER_20_1447 ();
 sg13g2_decap_8 FILLER_20_1454 ();
 sg13g2_decap_8 FILLER_20_1461 ();
 sg13g2_decap_8 FILLER_20_1468 ();
 sg13g2_decap_8 FILLER_20_1475 ();
 sg13g2_decap_8 FILLER_20_1482 ();
 sg13g2_decap_8 FILLER_20_1489 ();
 sg13g2_decap_8 FILLER_20_1496 ();
 sg13g2_decap_8 FILLER_20_1503 ();
 sg13g2_decap_8 FILLER_20_1510 ();
 sg13g2_decap_8 FILLER_20_1517 ();
 sg13g2_decap_8 FILLER_20_1524 ();
 sg13g2_decap_8 FILLER_20_1531 ();
 sg13g2_decap_8 FILLER_20_1538 ();
 sg13g2_decap_8 FILLER_20_1545 ();
 sg13g2_decap_8 FILLER_20_1552 ();
 sg13g2_decap_8 FILLER_20_1559 ();
 sg13g2_decap_8 FILLER_20_1566 ();
 sg13g2_decap_8 FILLER_20_1573 ();
 sg13g2_decap_8 FILLER_20_1580 ();
 sg13g2_decap_8 FILLER_20_1587 ();
 sg13g2_decap_8 FILLER_20_1594 ();
 sg13g2_decap_8 FILLER_20_1601 ();
 sg13g2_decap_8 FILLER_20_1608 ();
 sg13g2_decap_8 FILLER_20_1615 ();
 sg13g2_fill_2 FILLER_20_1622 ();
 sg13g2_fill_1 FILLER_20_1624 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_fill_2 FILLER_21_404 ();
 sg13g2_decap_8 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_417 ();
 sg13g2_decap_4 FILLER_21_433 ();
 sg13g2_decap_4 FILLER_21_446 ();
 sg13g2_fill_1 FILLER_21_450 ();
 sg13g2_decap_8 FILLER_21_506 ();
 sg13g2_fill_1 FILLER_21_539 ();
 sg13g2_fill_1 FILLER_21_587 ();
 sg13g2_fill_2 FILLER_21_598 ();
 sg13g2_decap_4 FILLER_21_651 ();
 sg13g2_fill_2 FILLER_21_665 ();
 sg13g2_decap_4 FILLER_21_698 ();
 sg13g2_fill_1 FILLER_21_702 ();
 sg13g2_decap_8 FILLER_21_708 ();
 sg13g2_decap_4 FILLER_21_715 ();
 sg13g2_fill_2 FILLER_21_719 ();
 sg13g2_decap_4 FILLER_21_725 ();
 sg13g2_fill_1 FILLER_21_729 ();
 sg13g2_decap_8 FILLER_21_734 ();
 sg13g2_fill_2 FILLER_21_741 ();
 sg13g2_fill_1 FILLER_21_743 ();
 sg13g2_fill_1 FILLER_21_773 ();
 sg13g2_decap_8 FILLER_21_779 ();
 sg13g2_fill_1 FILLER_21_786 ();
 sg13g2_fill_2 FILLER_21_796 ();
 sg13g2_fill_2 FILLER_21_832 ();
 sg13g2_decap_4 FILLER_21_838 ();
 sg13g2_decap_8 FILLER_21_846 ();
 sg13g2_decap_8 FILLER_21_853 ();
 sg13g2_decap_8 FILLER_21_860 ();
 sg13g2_fill_1 FILLER_21_867 ();
 sg13g2_decap_4 FILLER_21_873 ();
 sg13g2_fill_2 FILLER_21_881 ();
 sg13g2_fill_1 FILLER_21_883 ();
 sg13g2_decap_8 FILLER_21_889 ();
 sg13g2_decap_4 FILLER_21_896 ();
 sg13g2_fill_2 FILLER_21_900 ();
 sg13g2_fill_1 FILLER_21_978 ();
 sg13g2_decap_8 FILLER_21_983 ();
 sg13g2_decap_8 FILLER_21_990 ();
 sg13g2_decap_4 FILLER_21_997 ();
 sg13g2_fill_1 FILLER_21_1001 ();
 sg13g2_decap_8 FILLER_21_1028 ();
 sg13g2_decap_8 FILLER_21_1035 ();
 sg13g2_fill_2 FILLER_21_1042 ();
 sg13g2_fill_1 FILLER_21_1044 ();
 sg13g2_decap_8 FILLER_21_1071 ();
 sg13g2_decap_4 FILLER_21_1078 ();
 sg13g2_fill_1 FILLER_21_1082 ();
 sg13g2_decap_8 FILLER_21_1087 ();
 sg13g2_decap_8 FILLER_21_1140 ();
 sg13g2_decap_8 FILLER_21_1147 ();
 sg13g2_fill_2 FILLER_21_1187 ();
 sg13g2_fill_2 FILLER_21_1215 ();
 sg13g2_fill_1 FILLER_21_1217 ();
 sg13g2_fill_2 FILLER_21_1269 ();
 sg13g2_fill_1 FILLER_21_1271 ();
 sg13g2_decap_8 FILLER_21_1298 ();
 sg13g2_decap_8 FILLER_21_1305 ();
 sg13g2_decap_8 FILLER_21_1312 ();
 sg13g2_decap_8 FILLER_21_1319 ();
 sg13g2_decap_8 FILLER_21_1326 ();
 sg13g2_decap_8 FILLER_21_1333 ();
 sg13g2_decap_8 FILLER_21_1340 ();
 sg13g2_decap_8 FILLER_21_1347 ();
 sg13g2_decap_8 FILLER_21_1354 ();
 sg13g2_decap_8 FILLER_21_1361 ();
 sg13g2_decap_8 FILLER_21_1368 ();
 sg13g2_decap_8 FILLER_21_1375 ();
 sg13g2_decap_8 FILLER_21_1382 ();
 sg13g2_decap_8 FILLER_21_1389 ();
 sg13g2_decap_8 FILLER_21_1396 ();
 sg13g2_decap_8 FILLER_21_1403 ();
 sg13g2_decap_8 FILLER_21_1410 ();
 sg13g2_decap_8 FILLER_21_1417 ();
 sg13g2_decap_8 FILLER_21_1424 ();
 sg13g2_decap_8 FILLER_21_1431 ();
 sg13g2_decap_8 FILLER_21_1438 ();
 sg13g2_decap_8 FILLER_21_1445 ();
 sg13g2_decap_8 FILLER_21_1452 ();
 sg13g2_decap_8 FILLER_21_1459 ();
 sg13g2_decap_8 FILLER_21_1466 ();
 sg13g2_decap_8 FILLER_21_1473 ();
 sg13g2_decap_8 FILLER_21_1480 ();
 sg13g2_decap_8 FILLER_21_1487 ();
 sg13g2_decap_8 FILLER_21_1494 ();
 sg13g2_decap_8 FILLER_21_1501 ();
 sg13g2_decap_8 FILLER_21_1508 ();
 sg13g2_decap_8 FILLER_21_1515 ();
 sg13g2_decap_8 FILLER_21_1522 ();
 sg13g2_decap_8 FILLER_21_1529 ();
 sg13g2_decap_8 FILLER_21_1536 ();
 sg13g2_decap_8 FILLER_21_1543 ();
 sg13g2_decap_8 FILLER_21_1550 ();
 sg13g2_decap_8 FILLER_21_1557 ();
 sg13g2_decap_8 FILLER_21_1564 ();
 sg13g2_decap_8 FILLER_21_1571 ();
 sg13g2_decap_8 FILLER_21_1578 ();
 sg13g2_decap_8 FILLER_21_1585 ();
 sg13g2_decap_8 FILLER_21_1592 ();
 sg13g2_decap_8 FILLER_21_1599 ();
 sg13g2_decap_8 FILLER_21_1606 ();
 sg13g2_decap_8 FILLER_21_1613 ();
 sg13g2_decap_4 FILLER_21_1620 ();
 sg13g2_fill_1 FILLER_21_1624 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_fill_2 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_fill_2 FILLER_22_301 ();
 sg13g2_decap_4 FILLER_22_307 ();
 sg13g2_fill_1 FILLER_22_311 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_fill_1 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_352 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_373 ();
 sg13g2_decap_4 FILLER_22_380 ();
 sg13g2_fill_2 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_fill_2 FILLER_22_397 ();
 sg13g2_fill_1 FILLER_22_399 ();
 sg13g2_decap_4 FILLER_22_426 ();
 sg13g2_decap_8 FILLER_22_439 ();
 sg13g2_decap_8 FILLER_22_446 ();
 sg13g2_decap_8 FILLER_22_453 ();
 sg13g2_fill_1 FILLER_22_460 ();
 sg13g2_decap_4 FILLER_22_465 ();
 sg13g2_fill_2 FILLER_22_469 ();
 sg13g2_decap_4 FILLER_22_476 ();
 sg13g2_fill_1 FILLER_22_480 ();
 sg13g2_fill_2 FILLER_22_485 ();
 sg13g2_decap_8 FILLER_22_491 ();
 sg13g2_decap_8 FILLER_22_498 ();
 sg13g2_decap_8 FILLER_22_505 ();
 sg13g2_decap_8 FILLER_22_517 ();
 sg13g2_fill_1 FILLER_22_591 ();
 sg13g2_decap_8 FILLER_22_622 ();
 sg13g2_decap_4 FILLER_22_629 ();
 sg13g2_decap_4 FILLER_22_643 ();
 sg13g2_fill_2 FILLER_22_647 ();
 sg13g2_fill_1 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_685 ();
 sg13g2_fill_1 FILLER_22_692 ();
 sg13g2_decap_4 FILLER_22_714 ();
 sg13g2_fill_2 FILLER_22_752 ();
 sg13g2_fill_2 FILLER_22_785 ();
 sg13g2_decap_4 FILLER_22_822 ();
 sg13g2_fill_1 FILLER_22_826 ();
 sg13g2_decap_4 FILLER_22_853 ();
 sg13g2_fill_1 FILLER_22_857 ();
 sg13g2_fill_2 FILLER_22_884 ();
 sg13g2_fill_1 FILLER_22_886 ();
 sg13g2_decap_8 FILLER_22_918 ();
 sg13g2_fill_1 FILLER_22_925 ();
 sg13g2_decap_8 FILLER_22_949 ();
 sg13g2_fill_2 FILLER_22_956 ();
 sg13g2_fill_2 FILLER_22_962 ();
 sg13g2_fill_1 FILLER_22_964 ();
 sg13g2_fill_2 FILLER_22_999 ();
 sg13g2_decap_4 FILLER_22_1027 ();
 sg13g2_fill_2 FILLER_22_1031 ();
 sg13g2_fill_2 FILLER_22_1047 ();
 sg13g2_fill_1 FILLER_22_1049 ();
 sg13g2_decap_4 FILLER_22_1071 ();
 sg13g2_fill_1 FILLER_22_1075 ();
 sg13g2_fill_1 FILLER_22_1102 ();
 sg13g2_decap_8 FILLER_22_1124 ();
 sg13g2_decap_8 FILLER_22_1131 ();
 sg13g2_fill_1 FILLER_22_1138 ();
 sg13g2_decap_8 FILLER_22_1143 ();
 sg13g2_decap_8 FILLER_22_1150 ();
 sg13g2_decap_4 FILLER_22_1157 ();
 sg13g2_decap_8 FILLER_22_1182 ();
 sg13g2_fill_2 FILLER_22_1189 ();
 sg13g2_decap_8 FILLER_22_1229 ();
 sg13g2_fill_1 FILLER_22_1236 ();
 sg13g2_fill_2 FILLER_22_1267 ();
 sg13g2_fill_1 FILLER_22_1269 ();
 sg13g2_decap_8 FILLER_22_1304 ();
 sg13g2_decap_8 FILLER_22_1311 ();
 sg13g2_decap_8 FILLER_22_1318 ();
 sg13g2_decap_8 FILLER_22_1325 ();
 sg13g2_decap_8 FILLER_22_1332 ();
 sg13g2_decap_8 FILLER_22_1339 ();
 sg13g2_decap_8 FILLER_22_1346 ();
 sg13g2_decap_8 FILLER_22_1353 ();
 sg13g2_decap_8 FILLER_22_1360 ();
 sg13g2_decap_8 FILLER_22_1367 ();
 sg13g2_decap_8 FILLER_22_1374 ();
 sg13g2_decap_8 FILLER_22_1381 ();
 sg13g2_decap_8 FILLER_22_1388 ();
 sg13g2_decap_8 FILLER_22_1395 ();
 sg13g2_decap_8 FILLER_22_1402 ();
 sg13g2_decap_8 FILLER_22_1409 ();
 sg13g2_decap_8 FILLER_22_1416 ();
 sg13g2_decap_8 FILLER_22_1423 ();
 sg13g2_decap_8 FILLER_22_1430 ();
 sg13g2_decap_8 FILLER_22_1437 ();
 sg13g2_decap_8 FILLER_22_1444 ();
 sg13g2_decap_8 FILLER_22_1451 ();
 sg13g2_decap_8 FILLER_22_1458 ();
 sg13g2_decap_8 FILLER_22_1465 ();
 sg13g2_decap_8 FILLER_22_1472 ();
 sg13g2_decap_8 FILLER_22_1479 ();
 sg13g2_decap_8 FILLER_22_1486 ();
 sg13g2_decap_8 FILLER_22_1493 ();
 sg13g2_decap_8 FILLER_22_1500 ();
 sg13g2_decap_8 FILLER_22_1507 ();
 sg13g2_decap_8 FILLER_22_1514 ();
 sg13g2_decap_8 FILLER_22_1521 ();
 sg13g2_decap_8 FILLER_22_1528 ();
 sg13g2_decap_8 FILLER_22_1535 ();
 sg13g2_decap_8 FILLER_22_1542 ();
 sg13g2_decap_8 FILLER_22_1549 ();
 sg13g2_decap_8 FILLER_22_1556 ();
 sg13g2_decap_8 FILLER_22_1563 ();
 sg13g2_decap_8 FILLER_22_1570 ();
 sg13g2_decap_8 FILLER_22_1577 ();
 sg13g2_decap_8 FILLER_22_1584 ();
 sg13g2_decap_8 FILLER_22_1591 ();
 sg13g2_decap_8 FILLER_22_1598 ();
 sg13g2_decap_8 FILLER_22_1605 ();
 sg13g2_decap_8 FILLER_22_1612 ();
 sg13g2_decap_4 FILLER_22_1619 ();
 sg13g2_fill_2 FILLER_22_1623 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_fill_1 FILLER_23_342 ();
 sg13g2_decap_4 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_8 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_410 ();
 sg13g2_fill_1 FILLER_23_412 ();
 sg13g2_decap_8 FILLER_23_417 ();
 sg13g2_fill_2 FILLER_23_424 ();
 sg13g2_fill_1 FILLER_23_426 ();
 sg13g2_fill_1 FILLER_23_453 ();
 sg13g2_decap_8 FILLER_23_531 ();
 sg13g2_decap_4 FILLER_23_538 ();
 sg13g2_fill_2 FILLER_23_542 ();
 sg13g2_fill_2 FILLER_23_549 ();
 sg13g2_decap_8 FILLER_23_559 ();
 sg13g2_fill_1 FILLER_23_566 ();
 sg13g2_decap_8 FILLER_23_572 ();
 sg13g2_decap_8 FILLER_23_579 ();
 sg13g2_decap_4 FILLER_23_586 ();
 sg13g2_fill_2 FILLER_23_590 ();
 sg13g2_fill_2 FILLER_23_597 ();
 sg13g2_decap_4 FILLER_23_639 ();
 sg13g2_decap_8 FILLER_23_648 ();
 sg13g2_decap_8 FILLER_23_655 ();
 sg13g2_decap_8 FILLER_23_662 ();
 sg13g2_decap_8 FILLER_23_669 ();
 sg13g2_decap_8 FILLER_23_676 ();
 sg13g2_decap_8 FILLER_23_683 ();
 sg13g2_decap_4 FILLER_23_690 ();
 sg13g2_fill_1 FILLER_23_694 ();
 sg13g2_decap_8 FILLER_23_716 ();
 sg13g2_decap_8 FILLER_23_723 ();
 sg13g2_decap_8 FILLER_23_730 ();
 sg13g2_fill_2 FILLER_23_737 ();
 sg13g2_fill_1 FILLER_23_739 ();
 sg13g2_decap_4 FILLER_23_794 ();
 sg13g2_fill_2 FILLER_23_862 ();
 sg13g2_fill_1 FILLER_23_868 ();
 sg13g2_fill_1 FILLER_23_895 ();
 sg13g2_decap_8 FILLER_23_913 ();
 sg13g2_fill_2 FILLER_23_920 ();
 sg13g2_fill_1 FILLER_23_922 ();
 sg13g2_fill_2 FILLER_23_949 ();
 sg13g2_fill_2 FILLER_23_956 ();
 sg13g2_decap_8 FILLER_23_997 ();
 sg13g2_decap_8 FILLER_23_1004 ();
 sg13g2_fill_2 FILLER_23_1018 ();
 sg13g2_decap_8 FILLER_23_1046 ();
 sg13g2_decap_8 FILLER_23_1053 ();
 sg13g2_decap_8 FILLER_23_1060 ();
 sg13g2_decap_8 FILLER_23_1067 ();
 sg13g2_decap_4 FILLER_23_1074 ();
 sg13g2_fill_2 FILLER_23_1078 ();
 sg13g2_decap_4 FILLER_23_1089 ();
 sg13g2_fill_1 FILLER_23_1093 ();
 sg13g2_fill_2 FILLER_23_1124 ();
 sg13g2_fill_1 FILLER_23_1126 ();
 sg13g2_decap_8 FILLER_23_1158 ();
 sg13g2_decap_8 FILLER_23_1165 ();
 sg13g2_decap_4 FILLER_23_1172 ();
 sg13g2_fill_1 FILLER_23_1176 ();
 sg13g2_decap_4 FILLER_23_1198 ();
 sg13g2_decap_8 FILLER_23_1223 ();
 sg13g2_decap_4 FILLER_23_1230 ();
 sg13g2_fill_2 FILLER_23_1234 ();
 sg13g2_fill_2 FILLER_23_1241 ();
 sg13g2_fill_1 FILLER_23_1243 ();
 sg13g2_fill_1 FILLER_23_1269 ();
 sg13g2_fill_2 FILLER_23_1279 ();
 sg13g2_fill_1 FILLER_23_1281 ();
 sg13g2_decap_8 FILLER_23_1308 ();
 sg13g2_decap_8 FILLER_23_1315 ();
 sg13g2_decap_8 FILLER_23_1322 ();
 sg13g2_decap_8 FILLER_23_1329 ();
 sg13g2_decap_8 FILLER_23_1336 ();
 sg13g2_decap_8 FILLER_23_1343 ();
 sg13g2_decap_8 FILLER_23_1350 ();
 sg13g2_decap_8 FILLER_23_1357 ();
 sg13g2_decap_8 FILLER_23_1364 ();
 sg13g2_decap_8 FILLER_23_1371 ();
 sg13g2_decap_8 FILLER_23_1378 ();
 sg13g2_decap_8 FILLER_23_1385 ();
 sg13g2_decap_8 FILLER_23_1392 ();
 sg13g2_decap_8 FILLER_23_1399 ();
 sg13g2_decap_8 FILLER_23_1406 ();
 sg13g2_decap_8 FILLER_23_1413 ();
 sg13g2_decap_8 FILLER_23_1420 ();
 sg13g2_decap_8 FILLER_23_1427 ();
 sg13g2_decap_8 FILLER_23_1434 ();
 sg13g2_decap_8 FILLER_23_1441 ();
 sg13g2_decap_8 FILLER_23_1448 ();
 sg13g2_decap_8 FILLER_23_1455 ();
 sg13g2_decap_8 FILLER_23_1462 ();
 sg13g2_decap_8 FILLER_23_1469 ();
 sg13g2_decap_8 FILLER_23_1476 ();
 sg13g2_decap_8 FILLER_23_1483 ();
 sg13g2_decap_8 FILLER_23_1490 ();
 sg13g2_decap_8 FILLER_23_1497 ();
 sg13g2_decap_8 FILLER_23_1504 ();
 sg13g2_decap_8 FILLER_23_1511 ();
 sg13g2_decap_8 FILLER_23_1518 ();
 sg13g2_decap_8 FILLER_23_1525 ();
 sg13g2_decap_8 FILLER_23_1532 ();
 sg13g2_decap_8 FILLER_23_1539 ();
 sg13g2_decap_8 FILLER_23_1546 ();
 sg13g2_decap_8 FILLER_23_1553 ();
 sg13g2_decap_8 FILLER_23_1560 ();
 sg13g2_decap_8 FILLER_23_1567 ();
 sg13g2_decap_8 FILLER_23_1574 ();
 sg13g2_decap_8 FILLER_23_1581 ();
 sg13g2_decap_8 FILLER_23_1588 ();
 sg13g2_decap_8 FILLER_23_1595 ();
 sg13g2_decap_8 FILLER_23_1602 ();
 sg13g2_decap_8 FILLER_23_1609 ();
 sg13g2_decap_8 FILLER_23_1616 ();
 sg13g2_fill_2 FILLER_23_1623 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_4 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_4 FILLER_24_340 ();
 sg13g2_fill_2 FILLER_24_365 ();
 sg13g2_fill_1 FILLER_24_367 ();
 sg13g2_fill_2 FILLER_24_398 ();
 sg13g2_fill_1 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_433 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_4 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_527 ();
 sg13g2_decap_4 FILLER_24_534 ();
 sg13g2_decap_4 FILLER_24_564 ();
 sg13g2_decap_4 FILLER_24_577 ();
 sg13g2_fill_2 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_587 ();
 sg13g2_decap_4 FILLER_24_594 ();
 sg13g2_fill_2 FILLER_24_598 ();
 sg13g2_decap_8 FILLER_24_605 ();
 sg13g2_decap_8 FILLER_24_612 ();
 sg13g2_fill_2 FILLER_24_619 ();
 sg13g2_fill_1 FILLER_24_621 ();
 sg13g2_decap_8 FILLER_24_626 ();
 sg13g2_decap_4 FILLER_24_633 ();
 sg13g2_decap_8 FILLER_24_642 ();
 sg13g2_decap_8 FILLER_24_649 ();
 sg13g2_decap_4 FILLER_24_656 ();
 sg13g2_decap_4 FILLER_24_665 ();
 sg13g2_fill_1 FILLER_24_669 ();
 sg13g2_decap_8 FILLER_24_674 ();
 sg13g2_fill_2 FILLER_24_681 ();
 sg13g2_fill_1 FILLER_24_683 ();
 sg13g2_decap_4 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_701 ();
 sg13g2_decap_8 FILLER_24_708 ();
 sg13g2_fill_2 FILLER_24_715 ();
 sg13g2_fill_1 FILLER_24_722 ();
 sg13g2_fill_2 FILLER_24_727 ();
 sg13g2_fill_2 FILLER_24_733 ();
 sg13g2_fill_2 FILLER_24_740 ();
 sg13g2_fill_1 FILLER_24_742 ();
 sg13g2_fill_1 FILLER_24_752 ();
 sg13g2_decap_8 FILLER_24_757 ();
 sg13g2_decap_4 FILLER_24_769 ();
 sg13g2_fill_2 FILLER_24_773 ();
 sg13g2_fill_2 FILLER_24_837 ();
 sg13g2_fill_1 FILLER_24_890 ();
 sg13g2_fill_1 FILLER_24_916 ();
 sg13g2_fill_1 FILLER_24_963 ();
 sg13g2_fill_2 FILLER_24_993 ();
 sg13g2_fill_1 FILLER_24_1026 ();
 sg13g2_decap_8 FILLER_24_1031 ();
 sg13g2_fill_2 FILLER_24_1038 ();
 sg13g2_fill_2 FILLER_24_1045 ();
 sg13g2_decap_8 FILLER_24_1051 ();
 sg13g2_fill_1 FILLER_24_1058 ();
 sg13g2_decap_8 FILLER_24_1063 ();
 sg13g2_decap_8 FILLER_24_1070 ();
 sg13g2_decap_4 FILLER_24_1077 ();
 sg13g2_fill_1 FILLER_24_1081 ();
 sg13g2_decap_8 FILLER_24_1127 ();
 sg13g2_decap_8 FILLER_24_1147 ();
 sg13g2_decap_4 FILLER_24_1154 ();
 sg13g2_fill_1 FILLER_24_1158 ();
 sg13g2_decap_8 FILLER_24_1163 ();
 sg13g2_decap_4 FILLER_24_1170 ();
 sg13g2_fill_2 FILLER_24_1199 ();
 sg13g2_fill_1 FILLER_24_1201 ();
 sg13g2_decap_8 FILLER_24_1265 ();
 sg13g2_fill_2 FILLER_24_1272 ();
 sg13g2_fill_1 FILLER_24_1274 ();
 sg13g2_fill_1 FILLER_24_1279 ();
 sg13g2_fill_2 FILLER_24_1309 ();
 sg13g2_fill_1 FILLER_24_1311 ();
 sg13g2_decap_8 FILLER_24_1316 ();
 sg13g2_decap_8 FILLER_24_1323 ();
 sg13g2_decap_8 FILLER_24_1330 ();
 sg13g2_decap_8 FILLER_24_1337 ();
 sg13g2_decap_8 FILLER_24_1344 ();
 sg13g2_decap_8 FILLER_24_1351 ();
 sg13g2_decap_8 FILLER_24_1358 ();
 sg13g2_decap_8 FILLER_24_1365 ();
 sg13g2_decap_8 FILLER_24_1372 ();
 sg13g2_decap_8 FILLER_24_1379 ();
 sg13g2_decap_8 FILLER_24_1386 ();
 sg13g2_decap_8 FILLER_24_1393 ();
 sg13g2_decap_8 FILLER_24_1400 ();
 sg13g2_decap_8 FILLER_24_1407 ();
 sg13g2_decap_8 FILLER_24_1414 ();
 sg13g2_decap_8 FILLER_24_1421 ();
 sg13g2_decap_8 FILLER_24_1428 ();
 sg13g2_decap_4 FILLER_24_1435 ();
 sg13g2_fill_1 FILLER_24_1439 ();
 sg13g2_decap_8 FILLER_24_1444 ();
 sg13g2_decap_8 FILLER_24_1451 ();
 sg13g2_decap_8 FILLER_24_1458 ();
 sg13g2_decap_8 FILLER_24_1465 ();
 sg13g2_decap_8 FILLER_24_1472 ();
 sg13g2_decap_8 FILLER_24_1479 ();
 sg13g2_decap_4 FILLER_24_1486 ();
 sg13g2_decap_8 FILLER_24_1494 ();
 sg13g2_decap_8 FILLER_24_1526 ();
 sg13g2_decap_8 FILLER_24_1533 ();
 sg13g2_decap_8 FILLER_24_1540 ();
 sg13g2_decap_8 FILLER_24_1547 ();
 sg13g2_decap_8 FILLER_24_1554 ();
 sg13g2_decap_8 FILLER_24_1561 ();
 sg13g2_decap_8 FILLER_24_1568 ();
 sg13g2_decap_8 FILLER_24_1575 ();
 sg13g2_decap_8 FILLER_24_1582 ();
 sg13g2_decap_8 FILLER_24_1589 ();
 sg13g2_decap_8 FILLER_24_1596 ();
 sg13g2_decap_8 FILLER_24_1603 ();
 sg13g2_decap_8 FILLER_24_1610 ();
 sg13g2_decap_8 FILLER_24_1617 ();
 sg13g2_fill_1 FILLER_24_1624 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_4 FILLER_25_238 ();
 sg13g2_fill_1 FILLER_25_242 ();
 sg13g2_decap_8 FILLER_25_247 ();
 sg13g2_decap_8 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_263 ();
 sg13g2_decap_8 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_fill_1 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_fill_2 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_563 ();
 sg13g2_decap_4 FILLER_25_570 ();
 sg13g2_fill_1 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_601 ();
 sg13g2_decap_4 FILLER_25_608 ();
 sg13g2_fill_1 FILLER_25_612 ();
 sg13g2_decap_4 FILLER_25_643 ();
 sg13g2_fill_2 FILLER_25_647 ();
 sg13g2_decap_4 FILLER_25_710 ();
 sg13g2_fill_1 FILLER_25_714 ();
 sg13g2_fill_1 FILLER_25_719 ();
 sg13g2_fill_1 FILLER_25_772 ();
 sg13g2_fill_2 FILLER_25_778 ();
 sg13g2_fill_2 FILLER_25_784 ();
 sg13g2_fill_2 FILLER_25_790 ();
 sg13g2_fill_1 FILLER_25_792 ();
 sg13g2_fill_2 FILLER_25_848 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_decap_4 FILLER_25_870 ();
 sg13g2_fill_1 FILLER_25_900 ();
 sg13g2_fill_2 FILLER_25_927 ();
 sg13g2_fill_1 FILLER_25_929 ();
 sg13g2_decap_8 FILLER_25_951 ();
 sg13g2_fill_2 FILLER_25_958 ();
 sg13g2_fill_1 FILLER_25_960 ();
 sg13g2_decap_8 FILLER_25_996 ();
 sg13g2_decap_4 FILLER_25_1007 ();
 sg13g2_fill_1 FILLER_25_1011 ();
 sg13g2_decap_4 FILLER_25_1037 ();
 sg13g2_fill_1 FILLER_25_1041 ();
 sg13g2_fill_2 FILLER_25_1068 ();
 sg13g2_fill_1 FILLER_25_1070 ();
 sg13g2_decap_8 FILLER_25_1075 ();
 sg13g2_fill_2 FILLER_25_1111 ();
 sg13g2_fill_1 FILLER_25_1113 ();
 sg13g2_fill_1 FILLER_25_1128 ();
 sg13g2_decap_8 FILLER_25_1168 ();
 sg13g2_fill_2 FILLER_25_1175 ();
 sg13g2_decap_8 FILLER_25_1206 ();
 sg13g2_decap_8 FILLER_25_1213 ();
 sg13g2_decap_8 FILLER_25_1220 ();
 sg13g2_decap_8 FILLER_25_1227 ();
 sg13g2_decap_8 FILLER_25_1234 ();
 sg13g2_fill_2 FILLER_25_1241 ();
 sg13g2_fill_1 FILLER_25_1243 ();
 sg13g2_decap_8 FILLER_25_1265 ();
 sg13g2_fill_2 FILLER_25_1272 ();
 sg13g2_fill_1 FILLER_25_1274 ();
 sg13g2_fill_2 FILLER_25_1301 ();
 sg13g2_fill_1 FILLER_25_1303 ();
 sg13g2_decap_8 FILLER_25_1330 ();
 sg13g2_decap_8 FILLER_25_1337 ();
 sg13g2_decap_8 FILLER_25_1344 ();
 sg13g2_decap_8 FILLER_25_1351 ();
 sg13g2_decap_8 FILLER_25_1358 ();
 sg13g2_decap_8 FILLER_25_1365 ();
 sg13g2_decap_8 FILLER_25_1372 ();
 sg13g2_decap_8 FILLER_25_1379 ();
 sg13g2_decap_8 FILLER_25_1386 ();
 sg13g2_decap_8 FILLER_25_1393 ();
 sg13g2_decap_8 FILLER_25_1400 ();
 sg13g2_decap_8 FILLER_25_1407 ();
 sg13g2_decap_8 FILLER_25_1414 ();
 sg13g2_decap_8 FILLER_25_1421 ();
 sg13g2_fill_2 FILLER_25_1428 ();
 sg13g2_fill_1 FILLER_25_1430 ();
 sg13g2_decap_4 FILLER_25_1457 ();
 sg13g2_fill_2 FILLER_25_1461 ();
 sg13g2_decap_8 FILLER_25_1471 ();
 sg13g2_decap_4 FILLER_25_1478 ();
 sg13g2_fill_1 FILLER_25_1482 ();
 sg13g2_decap_8 FILLER_25_1509 ();
 sg13g2_fill_2 FILLER_25_1516 ();
 sg13g2_decap_8 FILLER_25_1522 ();
 sg13g2_decap_8 FILLER_25_1529 ();
 sg13g2_decap_8 FILLER_25_1536 ();
 sg13g2_decap_8 FILLER_25_1543 ();
 sg13g2_decap_8 FILLER_25_1550 ();
 sg13g2_decap_8 FILLER_25_1557 ();
 sg13g2_decap_8 FILLER_25_1564 ();
 sg13g2_decap_8 FILLER_25_1571 ();
 sg13g2_decap_8 FILLER_25_1578 ();
 sg13g2_decap_8 FILLER_25_1585 ();
 sg13g2_decap_8 FILLER_25_1592 ();
 sg13g2_decap_8 FILLER_25_1599 ();
 sg13g2_decap_8 FILLER_25_1606 ();
 sg13g2_decap_8 FILLER_25_1613 ();
 sg13g2_decap_4 FILLER_25_1620 ();
 sg13g2_fill_1 FILLER_25_1624 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_4 FILLER_26_231 ();
 sg13g2_fill_2 FILLER_26_235 ();
 sg13g2_fill_2 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_265 ();
 sg13g2_decap_4 FILLER_26_292 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_8 FILLER_26_404 ();
 sg13g2_decap_8 FILLER_26_411 ();
 sg13g2_decap_8 FILLER_26_418 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_2 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_26_436 ();
 sg13g2_decap_4 FILLER_26_443 ();
 sg13g2_fill_1 FILLER_26_447 ();
 sg13g2_fill_1 FILLER_26_479 ();
 sg13g2_decap_4 FILLER_26_493 ();
 sg13g2_fill_2 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_503 ();
 sg13g2_decap_4 FILLER_26_510 ();
 sg13g2_fill_2 FILLER_26_514 ();
 sg13g2_fill_1 FILLER_26_547 ();
 sg13g2_fill_2 FILLER_26_552 ();
 sg13g2_decap_8 FILLER_26_575 ();
 sg13g2_decap_8 FILLER_26_587 ();
 sg13g2_fill_1 FILLER_26_594 ();
 sg13g2_fill_2 FILLER_26_600 ();
 sg13g2_fill_2 FILLER_26_623 ();
 sg13g2_fill_1 FILLER_26_625 ();
 sg13g2_fill_2 FILLER_26_631 ();
 sg13g2_fill_1 FILLER_26_633 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_4 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_736 ();
 sg13g2_decap_8 FILLER_26_743 ();
 sg13g2_decap_8 FILLER_26_750 ();
 sg13g2_decap_8 FILLER_26_757 ();
 sg13g2_decap_8 FILLER_26_764 ();
 sg13g2_decap_8 FILLER_26_771 ();
 sg13g2_decap_8 FILLER_26_778 ();
 sg13g2_decap_8 FILLER_26_785 ();
 sg13g2_fill_2 FILLER_26_792 ();
 sg13g2_fill_1 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_839 ();
 sg13g2_fill_2 FILLER_26_846 ();
 sg13g2_fill_1 FILLER_26_848 ();
 sg13g2_decap_8 FILLER_26_880 ();
 sg13g2_decap_8 FILLER_26_887 ();
 sg13g2_fill_1 FILLER_26_894 ();
 sg13g2_decap_8 FILLER_26_934 ();
 sg13g2_decap_8 FILLER_26_977 ();
 sg13g2_decap_4 FILLER_26_984 ();
 sg13g2_fill_1 FILLER_26_988 ();
 sg13g2_fill_1 FILLER_26_1003 ();
 sg13g2_decap_8 FILLER_26_1008 ();
 sg13g2_decap_8 FILLER_26_1015 ();
 sg13g2_decap_8 FILLER_26_1022 ();
 sg13g2_fill_1 FILLER_26_1029 ();
 sg13g2_decap_4 FILLER_26_1035 ();
 sg13g2_decap_4 FILLER_26_1043 ();
 sg13g2_fill_2 FILLER_26_1047 ();
 sg13g2_decap_4 FILLER_26_1053 ();
 sg13g2_fill_2 FILLER_26_1057 ();
 sg13g2_fill_2 FILLER_26_1090 ();
 sg13g2_fill_1 FILLER_26_1092 ();
 sg13g2_fill_2 FILLER_26_1124 ();
 sg13g2_decap_4 FILLER_26_1181 ();
 sg13g2_fill_2 FILLER_26_1185 ();
 sg13g2_decap_4 FILLER_26_1218 ();
 sg13g2_decap_8 FILLER_26_1227 ();
 sg13g2_decap_8 FILLER_26_1234 ();
 sg13g2_fill_2 FILLER_26_1241 ();
 sg13g2_fill_1 FILLER_26_1243 ();
 sg13g2_fill_2 FILLER_26_1278 ();
 sg13g2_fill_1 FILLER_26_1280 ();
 sg13g2_decap_8 FILLER_26_1307 ();
 sg13g2_decap_8 FILLER_26_1314 ();
 sg13g2_fill_2 FILLER_26_1321 ();
 sg13g2_decap_8 FILLER_26_1327 ();
 sg13g2_decap_8 FILLER_26_1334 ();
 sg13g2_decap_8 FILLER_26_1341 ();
 sg13g2_fill_2 FILLER_26_1348 ();
 sg13g2_fill_1 FILLER_26_1350 ();
 sg13g2_decap_8 FILLER_26_1355 ();
 sg13g2_decap_8 FILLER_26_1362 ();
 sg13g2_decap_8 FILLER_26_1369 ();
 sg13g2_decap_8 FILLER_26_1376 ();
 sg13g2_decap_4 FILLER_26_1383 ();
 sg13g2_decap_8 FILLER_26_1391 ();
 sg13g2_decap_8 FILLER_26_1398 ();
 sg13g2_decap_8 FILLER_26_1405 ();
 sg13g2_decap_8 FILLER_26_1412 ();
 sg13g2_decap_8 FILLER_26_1419 ();
 sg13g2_decap_8 FILLER_26_1426 ();
 sg13g2_decap_4 FILLER_26_1433 ();
 sg13g2_decap_8 FILLER_26_1441 ();
 sg13g2_fill_2 FILLER_26_1448 ();
 sg13g2_decap_8 FILLER_26_1485 ();
 sg13g2_decap_8 FILLER_26_1492 ();
 sg13g2_fill_2 FILLER_26_1499 ();
 sg13g2_decap_4 FILLER_26_1505 ();
 sg13g2_fill_1 FILLER_26_1509 ();
 sg13g2_decap_8 FILLER_26_1536 ();
 sg13g2_decap_8 FILLER_26_1543 ();
 sg13g2_decap_8 FILLER_26_1550 ();
 sg13g2_decap_8 FILLER_26_1557 ();
 sg13g2_decap_8 FILLER_26_1564 ();
 sg13g2_decap_8 FILLER_26_1571 ();
 sg13g2_decap_8 FILLER_26_1578 ();
 sg13g2_decap_8 FILLER_26_1585 ();
 sg13g2_decap_8 FILLER_26_1592 ();
 sg13g2_decap_8 FILLER_26_1599 ();
 sg13g2_decap_8 FILLER_26_1606 ();
 sg13g2_decap_8 FILLER_26_1613 ();
 sg13g2_decap_4 FILLER_26_1620 ();
 sg13g2_fill_1 FILLER_26_1624 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_4 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_decap_4 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_253 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_4 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_decap_8 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_286 ();
 sg13g2_decap_8 FILLER_27_293 ();
 sg13g2_fill_2 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_307 ();
 sg13g2_decap_8 FILLER_27_314 ();
 sg13g2_decap_8 FILLER_27_321 ();
 sg13g2_fill_1 FILLER_27_328 ();
 sg13g2_decap_4 FILLER_27_334 ();
 sg13g2_fill_1 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_decap_4 FILLER_27_422 ();
 sg13g2_decap_4 FILLER_27_447 ();
 sg13g2_fill_1 FILLER_27_451 ();
 sg13g2_decap_8 FILLER_27_509 ();
 sg13g2_decap_8 FILLER_27_521 ();
 sg13g2_decap_8 FILLER_27_528 ();
 sg13g2_decap_8 FILLER_27_535 ();
 sg13g2_decap_8 FILLER_27_542 ();
 sg13g2_decap_8 FILLER_27_549 ();
 sg13g2_decap_4 FILLER_27_556 ();
 sg13g2_decap_8 FILLER_27_606 ();
 sg13g2_decap_8 FILLER_27_613 ();
 sg13g2_decap_8 FILLER_27_620 ();
 sg13g2_decap_4 FILLER_27_627 ();
 sg13g2_fill_2 FILLER_27_631 ();
 sg13g2_decap_8 FILLER_27_654 ();
 sg13g2_decap_4 FILLER_27_661 ();
 sg13g2_fill_1 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_676 ();
 sg13g2_fill_1 FILLER_27_683 ();
 sg13g2_fill_2 FILLER_27_687 ();
 sg13g2_decap_8 FILLER_27_706 ();
 sg13g2_decap_4 FILLER_27_713 ();
 sg13g2_fill_1 FILLER_27_717 ();
 sg13g2_decap_8 FILLER_27_747 ();
 sg13g2_decap_8 FILLER_27_754 ();
 sg13g2_decap_4 FILLER_27_761 ();
 sg13g2_fill_1 FILLER_27_765 ();
 sg13g2_fill_2 FILLER_27_770 ();
 sg13g2_fill_1 FILLER_27_772 ();
 sg13g2_fill_2 FILLER_27_778 ();
 sg13g2_fill_1 FILLER_27_811 ();
 sg13g2_decap_8 FILLER_27_837 ();
 sg13g2_decap_8 FILLER_27_844 ();
 sg13g2_decap_8 FILLER_27_851 ();
 sg13g2_decap_8 FILLER_27_858 ();
 sg13g2_fill_1 FILLER_27_865 ();
 sg13g2_decap_8 FILLER_27_870 ();
 sg13g2_decap_8 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_27_884 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_decap_4 FILLER_27_898 ();
 sg13g2_fill_2 FILLER_27_902 ();
 sg13g2_fill_2 FILLER_27_934 ();
 sg13g2_fill_1 FILLER_27_936 ();
 sg13g2_fill_2 FILLER_27_958 ();
 sg13g2_fill_1 FILLER_27_991 ();
 sg13g2_fill_2 FILLER_27_1018 ();
 sg13g2_fill_2 FILLER_27_1046 ();
 sg13g2_decap_8 FILLER_27_1052 ();
 sg13g2_fill_2 FILLER_27_1059 ();
 sg13g2_decap_4 FILLER_27_1099 ();
 sg13g2_fill_1 FILLER_27_1103 ();
 sg13g2_decap_8 FILLER_27_1143 ();
 sg13g2_decap_8 FILLER_27_1150 ();
 sg13g2_decap_4 FILLER_27_1157 ();
 sg13g2_fill_2 FILLER_27_1161 ();
 sg13g2_fill_2 FILLER_27_1184 ();
 sg13g2_fill_1 FILLER_27_1186 ();
 sg13g2_decap_8 FILLER_27_1200 ();
 sg13g2_fill_2 FILLER_27_1207 ();
 sg13g2_fill_1 FILLER_27_1209 ();
 sg13g2_fill_1 FILLER_27_1215 ();
 sg13g2_decap_8 FILLER_27_1242 ();
 sg13g2_decap_8 FILLER_27_1253 ();
 sg13g2_decap_8 FILLER_27_1260 ();
 sg13g2_decap_4 FILLER_27_1267 ();
 sg13g2_fill_2 FILLER_27_1271 ();
 sg13g2_decap_8 FILLER_27_1278 ();
 sg13g2_decap_4 FILLER_27_1285 ();
 sg13g2_decap_8 FILLER_27_1293 ();
 sg13g2_decap_8 FILLER_27_1300 ();
 sg13g2_fill_1 FILLER_27_1307 ();
 sg13g2_decap_8 FILLER_27_1369 ();
 sg13g2_fill_2 FILLER_27_1376 ();
 sg13g2_fill_1 FILLER_27_1378 ();
 sg13g2_decap_8 FILLER_27_1405 ();
 sg13g2_decap_8 FILLER_27_1412 ();
 sg13g2_decap_4 FILLER_27_1419 ();
 sg13g2_fill_1 FILLER_27_1423 ();
 sg13g2_fill_1 FILLER_27_1509 ();
 sg13g2_decap_4 FILLER_27_1519 ();
 sg13g2_decap_8 FILLER_27_1527 ();
 sg13g2_fill_2 FILLER_27_1534 ();
 sg13g2_decap_8 FILLER_27_1540 ();
 sg13g2_decap_8 FILLER_27_1547 ();
 sg13g2_fill_1 FILLER_27_1554 ();
 sg13g2_decap_8 FILLER_27_1559 ();
 sg13g2_fill_2 FILLER_27_1566 ();
 sg13g2_decap_8 FILLER_27_1572 ();
 sg13g2_decap_8 FILLER_27_1579 ();
 sg13g2_decap_8 FILLER_27_1586 ();
 sg13g2_decap_8 FILLER_27_1593 ();
 sg13g2_decap_8 FILLER_27_1600 ();
 sg13g2_decap_8 FILLER_27_1607 ();
 sg13g2_decap_8 FILLER_27_1614 ();
 sg13g2_decap_4 FILLER_27_1621 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_4 FILLER_28_245 ();
 sg13g2_decap_4 FILLER_28_254 ();
 sg13g2_decap_8 FILLER_28_262 ();
 sg13g2_decap_4 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_310 ();
 sg13g2_decap_4 FILLER_28_317 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_fill_1 FILLER_28_331 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_4 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_decap_4 FILLER_28_373 ();
 sg13g2_fill_2 FILLER_28_377 ();
 sg13g2_fill_1 FILLER_28_447 ();
 sg13g2_decap_8 FILLER_28_511 ();
 sg13g2_fill_2 FILLER_28_518 ();
 sg13g2_fill_1 FILLER_28_520 ();
 sg13g2_decap_8 FILLER_28_530 ();
 sg13g2_decap_4 FILLER_28_537 ();
 sg13g2_decap_4 FILLER_28_546 ();
 sg13g2_fill_1 FILLER_28_550 ();
 sg13g2_decap_8 FILLER_28_581 ();
 sg13g2_fill_2 FILLER_28_588 ();
 sg13g2_decap_8 FILLER_28_611 ();
 sg13g2_decap_8 FILLER_28_618 ();
 sg13g2_decap_8 FILLER_28_625 ();
 sg13g2_decap_8 FILLER_28_632 ();
 sg13g2_decap_8 FILLER_28_639 ();
 sg13g2_decap_8 FILLER_28_646 ();
 sg13g2_decap_8 FILLER_28_653 ();
 sg13g2_decap_8 FILLER_28_660 ();
 sg13g2_decap_4 FILLER_28_667 ();
 sg13g2_fill_2 FILLER_28_671 ();
 sg13g2_decap_8 FILLER_28_678 ();
 sg13g2_decap_4 FILLER_28_685 ();
 sg13g2_decap_8 FILLER_28_715 ();
 sg13g2_fill_2 FILLER_28_726 ();
 sg13g2_decap_4 FILLER_28_789 ();
 sg13g2_fill_1 FILLER_28_793 ();
 sg13g2_fill_2 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_fill_2 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_835 ();
 sg13g2_decap_4 FILLER_28_842 ();
 sg13g2_fill_1 FILLER_28_846 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_fill_2 FILLER_28_858 ();
 sg13g2_decap_4 FILLER_28_896 ();
 sg13g2_fill_2 FILLER_28_900 ();
 sg13g2_decap_4 FILLER_28_906 ();
 sg13g2_decap_8 FILLER_28_945 ();
 sg13g2_decap_8 FILLER_28_952 ();
 sg13g2_fill_1 FILLER_28_959 ();
 sg13g2_decap_8 FILLER_28_964 ();
 sg13g2_fill_2 FILLER_28_971 ();
 sg13g2_fill_1 FILLER_28_977 ();
 sg13g2_decap_8 FILLER_28_1007 ();
 sg13g2_decap_8 FILLER_28_1014 ();
 sg13g2_decap_4 FILLER_28_1021 ();
 sg13g2_fill_1 FILLER_28_1025 ();
 sg13g2_decap_8 FILLER_28_1095 ();
 sg13g2_decap_4 FILLER_28_1102 ();
 sg13g2_decap_8 FILLER_28_1143 ();
 sg13g2_decap_8 FILLER_28_1150 ();
 sg13g2_fill_1 FILLER_28_1157 ();
 sg13g2_decap_4 FILLER_28_1184 ();
 sg13g2_fill_1 FILLER_28_1214 ();
 sg13g2_decap_4 FILLER_28_1267 ();
 sg13g2_fill_2 FILLER_28_1276 ();
 sg13g2_fill_1 FILLER_28_1278 ();
 sg13g2_decap_8 FILLER_28_1284 ();
 sg13g2_fill_2 FILLER_28_1291 ();
 sg13g2_fill_1 FILLER_28_1293 ();
 sg13g2_decap_4 FILLER_28_1299 ();
 sg13g2_fill_1 FILLER_28_1303 ();
 sg13g2_decap_4 FILLER_28_1308 ();
 sg13g2_decap_8 FILLER_28_1316 ();
 sg13g2_decap_8 FILLER_28_1323 ();
 sg13g2_decap_4 FILLER_28_1334 ();
 sg13g2_fill_2 FILLER_28_1338 ();
 sg13g2_fill_1 FILLER_28_1349 ();
 sg13g2_fill_2 FILLER_28_1355 ();
 sg13g2_fill_1 FILLER_28_1357 ();
 sg13g2_decap_8 FILLER_28_1362 ();
 sg13g2_decap_4 FILLER_28_1369 ();
 sg13g2_fill_2 FILLER_28_1373 ();
 sg13g2_fill_1 FILLER_28_1384 ();
 sg13g2_decap_8 FILLER_28_1389 ();
 sg13g2_decap_8 FILLER_28_1396 ();
 sg13g2_decap_8 FILLER_28_1403 ();
 sg13g2_decap_8 FILLER_28_1410 ();
 sg13g2_decap_8 FILLER_28_1417 ();
 sg13g2_decap_8 FILLER_28_1429 ();
 sg13g2_fill_1 FILLER_28_1436 ();
 sg13g2_fill_2 FILLER_28_1462 ();
 sg13g2_fill_1 FILLER_28_1464 ();
 sg13g2_fill_2 FILLER_28_1491 ();
 sg13g2_fill_1 FILLER_28_1493 ();
 sg13g2_fill_2 FILLER_28_1520 ();
 sg13g2_fill_1 FILLER_28_1522 ();
 sg13g2_fill_1 FILLER_28_1554 ();
 sg13g2_decap_8 FILLER_28_1586 ();
 sg13g2_decap_8 FILLER_28_1593 ();
 sg13g2_decap_8 FILLER_28_1600 ();
 sg13g2_decap_8 FILLER_28_1607 ();
 sg13g2_decap_8 FILLER_28_1614 ();
 sg13g2_decap_4 FILLER_28_1621 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_4 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_decap_8 FILLER_29_272 ();
 sg13g2_decap_4 FILLER_29_279 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_decap_4 FILLER_29_310 ();
 sg13g2_fill_1 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_decap_4 FILLER_29_377 ();
 sg13g2_fill_2 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_4 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_457 ();
 sg13g2_fill_1 FILLER_29_459 ();
 sg13g2_fill_1 FILLER_29_485 ();
 sg13g2_fill_1 FILLER_29_512 ();
 sg13g2_decap_8 FILLER_29_578 ();
 sg13g2_fill_1 FILLER_29_585 ();
 sg13g2_fill_2 FILLER_29_590 ();
 sg13g2_decap_8 FILLER_29_613 ();
 sg13g2_decap_8 FILLER_29_620 ();
 sg13g2_decap_4 FILLER_29_627 ();
 sg13g2_fill_2 FILLER_29_631 ();
 sg13g2_decap_8 FILLER_29_654 ();
 sg13g2_fill_2 FILLER_29_661 ();
 sg13g2_fill_1 FILLER_29_663 ();
 sg13g2_fill_2 FILLER_29_702 ();
 sg13g2_fill_1 FILLER_29_704 ();
 sg13g2_decap_8 FILLER_29_740 ();
 sg13g2_decap_8 FILLER_29_747 ();
 sg13g2_decap_8 FILLER_29_754 ();
 sg13g2_fill_1 FILLER_29_761 ();
 sg13g2_fill_2 FILLER_29_765 ();
 sg13g2_fill_1 FILLER_29_767 ();
 sg13g2_fill_2 FILLER_29_866 ();
 sg13g2_fill_2 FILLER_29_894 ();
 sg13g2_decap_8 FILLER_29_930 ();
 sg13g2_decap_8 FILLER_29_937 ();
 sg13g2_decap_8 FILLER_29_944 ();
 sg13g2_decap_8 FILLER_29_951 ();
 sg13g2_decap_4 FILLER_29_968 ();
 sg13g2_fill_2 FILLER_29_972 ();
 sg13g2_decap_4 FILLER_29_1000 ();
 sg13g2_decap_8 FILLER_29_1025 ();
 sg13g2_decap_8 FILLER_29_1032 ();
 sg13g2_fill_2 FILLER_29_1039 ();
 sg13g2_decap_8 FILLER_29_1067 ();
 sg13g2_decap_8 FILLER_29_1074 ();
 sg13g2_decap_8 FILLER_29_1081 ();
 sg13g2_decap_8 FILLER_29_1088 ();
 sg13g2_decap_4 FILLER_29_1095 ();
 sg13g2_fill_2 FILLER_29_1099 ();
 sg13g2_decap_8 FILLER_29_1166 ();
 sg13g2_decap_8 FILLER_29_1173 ();
 sg13g2_decap_8 FILLER_29_1180 ();
 sg13g2_decap_4 FILLER_29_1187 ();
 sg13g2_fill_2 FILLER_29_1241 ();
 sg13g2_decap_8 FILLER_29_1250 ();
 sg13g2_decap_8 FILLER_29_1257 ();
 sg13g2_decap_4 FILLER_29_1264 ();
 sg13g2_fill_1 FILLER_29_1294 ();
 sg13g2_fill_1 FILLER_29_1350 ();
 sg13g2_fill_2 FILLER_29_1376 ();
 sg13g2_fill_2 FILLER_29_1404 ();
 sg13g2_fill_1 FILLER_29_1406 ();
 sg13g2_decap_4 FILLER_29_1411 ();
 sg13g2_fill_1 FILLER_29_1415 ();
 sg13g2_fill_2 FILLER_29_1420 ();
 sg13g2_fill_1 FILLER_29_1422 ();
 sg13g2_decap_4 FILLER_29_1454 ();
 sg13g2_fill_1 FILLER_29_1467 ();
 sg13g2_decap_8 FILLER_29_1472 ();
 sg13g2_decap_8 FILLER_29_1479 ();
 sg13g2_decap_8 FILLER_29_1486 ();
 sg13g2_decap_8 FILLER_29_1502 ();
 sg13g2_decap_8 FILLER_29_1509 ();
 sg13g2_decap_8 FILLER_29_1516 ();
 sg13g2_decap_8 FILLER_29_1523 ();
 sg13g2_decap_8 FILLER_29_1559 ();
 sg13g2_fill_1 FILLER_29_1566 ();
 sg13g2_decap_8 FILLER_29_1576 ();
 sg13g2_decap_8 FILLER_29_1583 ();
 sg13g2_decap_8 FILLER_29_1590 ();
 sg13g2_decap_8 FILLER_29_1597 ();
 sg13g2_decap_8 FILLER_29_1604 ();
 sg13g2_decap_8 FILLER_29_1611 ();
 sg13g2_decap_8 FILLER_29_1618 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_230 ();
 sg13g2_decap_8 FILLER_30_237 ();
 sg13g2_decap_4 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_decap_8 FILLER_30_254 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_decap_4 FILLER_30_309 ();
 sg13g2_decap_8 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_30_331 ();
 sg13g2_fill_1 FILLER_30_338 ();
 sg13g2_fill_2 FILLER_30_381 ();
 sg13g2_fill_1 FILLER_30_383 ();
 sg13g2_fill_2 FILLER_30_430 ();
 sg13g2_fill_1 FILLER_30_432 ();
 sg13g2_decap_4 FILLER_30_506 ();
 sg13g2_fill_1 FILLER_30_510 ();
 sg13g2_fill_2 FILLER_30_515 ();
 sg13g2_fill_2 FILLER_30_546 ();
 sg13g2_fill_1 FILLER_30_548 ();
 sg13g2_decap_4 FILLER_30_553 ();
 sg13g2_fill_1 FILLER_30_557 ();
 sg13g2_fill_1 FILLER_30_592 ();
 sg13g2_decap_8 FILLER_30_597 ();
 sg13g2_decap_4 FILLER_30_604 ();
 sg13g2_fill_2 FILLER_30_608 ();
 sg13g2_decap_8 FILLER_30_662 ();
 sg13g2_fill_2 FILLER_30_669 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_fill_2 FILLER_30_686 ();
 sg13g2_fill_1 FILLER_30_688 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_fill_1 FILLER_30_721 ();
 sg13g2_decap_4 FILLER_30_727 ();
 sg13g2_fill_1 FILLER_30_756 ();
 sg13g2_fill_2 FILLER_30_812 ();
 sg13g2_fill_1 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_841 ();
 sg13g2_decap_8 FILLER_30_848 ();
 sg13g2_fill_1 FILLER_30_855 ();
 sg13g2_fill_2 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_30_913 ();
 sg13g2_fill_2 FILLER_30_920 ();
 sg13g2_decap_8 FILLER_30_943 ();
 sg13g2_decap_8 FILLER_30_950 ();
 sg13g2_decap_8 FILLER_30_957 ();
 sg13g2_decap_8 FILLER_30_964 ();
 sg13g2_fill_1 FILLER_30_971 ();
 sg13g2_decap_8 FILLER_30_977 ();
 sg13g2_fill_2 FILLER_30_984 ();
 sg13g2_decap_4 FILLER_30_990 ();
 sg13g2_decap_4 FILLER_30_1003 ();
 sg13g2_fill_1 FILLER_30_1007 ();
 sg13g2_decap_8 FILLER_30_1033 ();
 sg13g2_decap_8 FILLER_30_1040 ();
 sg13g2_decap_8 FILLER_30_1047 ();
 sg13g2_decap_8 FILLER_30_1054 ();
 sg13g2_decap_4 FILLER_30_1061 ();
 sg13g2_fill_1 FILLER_30_1065 ();
 sg13g2_decap_8 FILLER_30_1071 ();
 sg13g2_decap_8 FILLER_30_1078 ();
 sg13g2_fill_2 FILLER_30_1085 ();
 sg13g2_fill_2 FILLER_30_1116 ();
 sg13g2_decap_8 FILLER_30_1174 ();
 sg13g2_decap_8 FILLER_30_1181 ();
 sg13g2_fill_2 FILLER_30_1188 ();
 sg13g2_decap_8 FILLER_30_1197 ();
 sg13g2_fill_2 FILLER_30_1204 ();
 sg13g2_fill_1 FILLER_30_1206 ();
 sg13g2_decap_4 FILLER_30_1232 ();
 sg13g2_fill_1 FILLER_30_1236 ();
 sg13g2_fill_2 FILLER_30_1242 ();
 sg13g2_decap_4 FILLER_30_1282 ();
 sg13g2_fill_2 FILLER_30_1315 ();
 sg13g2_fill_1 FILLER_30_1317 ();
 sg13g2_fill_1 FILLER_30_1349 ();
 sg13g2_decap_4 FILLER_30_1381 ();
 sg13g2_fill_1 FILLER_30_1385 ();
 sg13g2_fill_2 FILLER_30_1390 ();
 sg13g2_decap_4 FILLER_30_1396 ();
 sg13g2_fill_1 FILLER_30_1431 ();
 sg13g2_decap_4 FILLER_30_1436 ();
 sg13g2_fill_1 FILLER_30_1440 ();
 sg13g2_decap_4 FILLER_30_1471 ();
 sg13g2_fill_2 FILLER_30_1475 ();
 sg13g2_fill_2 FILLER_30_1482 ();
 sg13g2_decap_4 FILLER_30_1489 ();
 sg13g2_decap_4 FILLER_30_1497 ();
 sg13g2_fill_2 FILLER_30_1501 ();
 sg13g2_decap_4 FILLER_30_1524 ();
 sg13g2_fill_2 FILLER_30_1528 ();
 sg13g2_decap_4 FILLER_30_1556 ();
 sg13g2_fill_2 FILLER_30_1560 ();
 sg13g2_decap_8 FILLER_30_1591 ();
 sg13g2_decap_8 FILLER_30_1598 ();
 sg13g2_decap_8 FILLER_30_1605 ();
 sg13g2_decap_8 FILLER_30_1612 ();
 sg13g2_decap_4 FILLER_30_1619 ();
 sg13g2_fill_2 FILLER_30_1623 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_fill_2 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_decap_4 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_fill_2 FILLER_31_324 ();
 sg13g2_decap_8 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_fill_2 FILLER_31_369 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_fill_1 FILLER_31_404 ();
 sg13g2_fill_2 FILLER_31_415 ();
 sg13g2_fill_1 FILLER_31_417 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_fill_2 FILLER_31_462 ();
 sg13g2_fill_1 FILLER_31_528 ();
 sg13g2_decap_8 FILLER_31_585 ();
 sg13g2_decap_8 FILLER_31_601 ();
 sg13g2_decap_8 FILLER_31_608 ();
 sg13g2_decap_4 FILLER_31_615 ();
 sg13g2_fill_2 FILLER_31_619 ();
 sg13g2_decap_4 FILLER_31_625 ();
 sg13g2_fill_1 FILLER_31_629 ();
 sg13g2_decap_8 FILLER_31_639 ();
 sg13g2_decap_8 FILLER_31_646 ();
 sg13g2_decap_8 FILLER_31_653 ();
 sg13g2_fill_2 FILLER_31_660 ();
 sg13g2_fill_1 FILLER_31_662 ();
 sg13g2_decap_8 FILLER_31_668 ();
 sg13g2_fill_1 FILLER_31_675 ();
 sg13g2_decap_4 FILLER_31_680 ();
 sg13g2_decap_4 FILLER_31_723 ();
 sg13g2_fill_1 FILLER_31_736 ();
 sg13g2_fill_2 FILLER_31_742 ();
 sg13g2_fill_1 FILLER_31_744 ();
 sg13g2_fill_1 FILLER_31_754 ();
 sg13g2_decap_8 FILLER_31_781 ();
 sg13g2_decap_8 FILLER_31_788 ();
 sg13g2_decap_8 FILLER_31_795 ();
 sg13g2_decap_8 FILLER_31_802 ();
 sg13g2_decap_4 FILLER_31_809 ();
 sg13g2_fill_1 FILLER_31_813 ();
 sg13g2_decap_8 FILLER_31_870 ();
 sg13g2_fill_2 FILLER_31_877 ();
 sg13g2_decap_4 FILLER_31_883 ();
 sg13g2_fill_2 FILLER_31_918 ();
 sg13g2_fill_1 FILLER_31_920 ();
 sg13g2_decap_8 FILLER_31_973 ();
 sg13g2_fill_1 FILLER_31_980 ();
 sg13g2_fill_1 FILLER_31_1006 ();
 sg13g2_decap_8 FILLER_31_1047 ();
 sg13g2_decap_4 FILLER_31_1054 ();
 sg13g2_decap_4 FILLER_31_1063 ();
 sg13g2_fill_1 FILLER_31_1071 ();
 sg13g2_fill_2 FILLER_31_1077 ();
 sg13g2_fill_2 FILLER_31_1178 ();
 sg13g2_decap_8 FILLER_31_1220 ();
 sg13g2_decap_8 FILLER_31_1227 ();
 sg13g2_fill_2 FILLER_31_1234 ();
 sg13g2_fill_1 FILLER_31_1236 ();
 sg13g2_decap_8 FILLER_31_1263 ();
 sg13g2_fill_2 FILLER_31_1310 ();
 sg13g2_fill_1 FILLER_31_1312 ();
 sg13g2_decap_8 FILLER_31_1334 ();
 sg13g2_decap_8 FILLER_31_1341 ();
 sg13g2_fill_2 FILLER_31_1348 ();
 sg13g2_fill_1 FILLER_31_1350 ();
 sg13g2_decap_8 FILLER_31_1355 ();
 sg13g2_decap_8 FILLER_31_1362 ();
 sg13g2_fill_2 FILLER_31_1369 ();
 sg13g2_fill_2 FILLER_31_1422 ();
 sg13g2_decap_4 FILLER_31_1429 ();
 sg13g2_fill_2 FILLER_31_1433 ();
 sg13g2_decap_4 FILLER_31_1524 ();
 sg13g2_fill_2 FILLER_31_1528 ();
 sg13g2_decap_4 FILLER_31_1539 ();
 sg13g2_fill_2 FILLER_31_1543 ();
 sg13g2_decap_8 FILLER_31_1606 ();
 sg13g2_decap_8 FILLER_31_1613 ();
 sg13g2_decap_4 FILLER_31_1620 ();
 sg13g2_fill_1 FILLER_31_1624 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_fill_2 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_237 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_decap_4 FILLER_32_276 ();
 sg13g2_fill_2 FILLER_32_280 ();
 sg13g2_fill_2 FILLER_32_320 ();
 sg13g2_decap_4 FILLER_32_374 ();
 sg13g2_fill_1 FILLER_32_378 ();
 sg13g2_fill_2 FILLER_32_384 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_8 FILLER_32_404 ();
 sg13g2_fill_2 FILLER_32_411 ();
 sg13g2_fill_2 FILLER_32_418 ();
 sg13g2_fill_1 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_435 ();
 sg13g2_fill_2 FILLER_32_442 ();
 sg13g2_fill_1 FILLER_32_444 ();
 sg13g2_fill_2 FILLER_32_450 ();
 sg13g2_decap_8 FILLER_32_506 ();
 sg13g2_decap_8 FILLER_32_513 ();
 sg13g2_decap_8 FILLER_32_520 ();
 sg13g2_decap_8 FILLER_32_527 ();
 sg13g2_fill_2 FILLER_32_534 ();
 sg13g2_fill_1 FILLER_32_536 ();
 sg13g2_decap_8 FILLER_32_541 ();
 sg13g2_decap_4 FILLER_32_548 ();
 sg13g2_fill_2 FILLER_32_552 ();
 sg13g2_decap_8 FILLER_32_559 ();
 sg13g2_fill_1 FILLER_32_566 ();
 sg13g2_decap_4 FILLER_32_571 ();
 sg13g2_fill_1 FILLER_32_575 ();
 sg13g2_fill_1 FILLER_32_581 ();
 sg13g2_decap_4 FILLER_32_586 ();
 sg13g2_decap_8 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_fill_1 FILLER_32_630 ();
 sg13g2_decap_8 FILLER_32_636 ();
 sg13g2_fill_2 FILLER_32_643 ();
 sg13g2_fill_1 FILLER_32_645 ();
 sg13g2_fill_2 FILLER_32_650 ();
 sg13g2_decap_8 FILLER_32_657 ();
 sg13g2_decap_4 FILLER_32_695 ();
 sg13g2_fill_2 FILLER_32_725 ();
 sg13g2_decap_4 FILLER_32_758 ();
 sg13g2_fill_1 FILLER_32_762 ();
 sg13g2_decap_8 FILLER_32_768 ();
 sg13g2_decap_8 FILLER_32_775 ();
 sg13g2_decap_8 FILLER_32_786 ();
 sg13g2_fill_1 FILLER_32_793 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_fill_2 FILLER_32_819 ();
 sg13g2_fill_1 FILLER_32_821 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_893 ();
 sg13g2_fill_2 FILLER_32_909 ();
 sg13g2_fill_1 FILLER_32_911 ();
 sg13g2_decap_8 FILLER_32_916 ();
 sg13g2_decap_8 FILLER_32_923 ();
 sg13g2_decap_8 FILLER_32_930 ();
 sg13g2_decap_8 FILLER_32_937 ();
 sg13g2_decap_8 FILLER_32_944 ();
 sg13g2_fill_2 FILLER_32_951 ();
 sg13g2_fill_1 FILLER_32_953 ();
 sg13g2_fill_1 FILLER_32_989 ();
 sg13g2_fill_2 FILLER_32_1020 ();
 sg13g2_fill_1 FILLER_32_1090 ();
 sg13g2_fill_2 FILLER_32_1095 ();
 sg13g2_decap_8 FILLER_32_1158 ();
 sg13g2_decap_8 FILLER_32_1170 ();
 sg13g2_fill_2 FILLER_32_1177 ();
 sg13g2_decap_8 FILLER_32_1184 ();
 sg13g2_decap_4 FILLER_32_1195 ();
 sg13g2_fill_1 FILLER_32_1199 ();
 sg13g2_fill_1 FILLER_32_1205 ();
 sg13g2_decap_8 FILLER_32_1210 ();
 sg13g2_decap_4 FILLER_32_1217 ();
 sg13g2_fill_1 FILLER_32_1221 ();
 sg13g2_decap_4 FILLER_32_1227 ();
 sg13g2_fill_1 FILLER_32_1235 ();
 sg13g2_decap_8 FILLER_32_1241 ();
 sg13g2_decap_8 FILLER_32_1248 ();
 sg13g2_decap_8 FILLER_32_1255 ();
 sg13g2_decap_4 FILLER_32_1262 ();
 sg13g2_fill_2 FILLER_32_1266 ();
 sg13g2_fill_2 FILLER_32_1281 ();
 sg13g2_fill_1 FILLER_32_1283 ();
 sg13g2_decap_8 FILLER_32_1335 ();
 sg13g2_decap_4 FILLER_32_1342 ();
 sg13g2_decap_8 FILLER_32_1350 ();
 sg13g2_fill_2 FILLER_32_1357 ();
 sg13g2_fill_1 FILLER_32_1359 ();
 sg13g2_decap_8 FILLER_32_1441 ();
 sg13g2_decap_4 FILLER_32_1448 ();
 sg13g2_fill_1 FILLER_32_1456 ();
 sg13g2_decap_4 FILLER_32_1478 ();
 sg13g2_fill_2 FILLER_32_1482 ();
 sg13g2_fill_2 FILLER_32_1488 ();
 sg13g2_fill_1 FILLER_32_1490 ();
 sg13g2_decap_8 FILLER_32_1495 ();
 sg13g2_decap_8 FILLER_32_1502 ();
 sg13g2_decap_8 FILLER_32_1509 ();
 sg13g2_decap_8 FILLER_32_1516 ();
 sg13g2_decap_8 FILLER_32_1523 ();
 sg13g2_decap_8 FILLER_32_1530 ();
 sg13g2_decap_8 FILLER_32_1537 ();
 sg13g2_decap_8 FILLER_32_1544 ();
 sg13g2_decap_8 FILLER_32_1551 ();
 sg13g2_fill_2 FILLER_32_1558 ();
 sg13g2_fill_1 FILLER_32_1560 ();
 sg13g2_decap_8 FILLER_32_1565 ();
 sg13g2_decap_8 FILLER_32_1572 ();
 sg13g2_decap_8 FILLER_32_1579 ();
 sg13g2_decap_8 FILLER_32_1586 ();
 sg13g2_decap_8 FILLER_32_1593 ();
 sg13g2_decap_8 FILLER_32_1600 ();
 sg13g2_decap_8 FILLER_32_1607 ();
 sg13g2_decap_8 FILLER_32_1614 ();
 sg13g2_decap_4 FILLER_32_1621 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_fill_2 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_253 ();
 sg13g2_decap_8 FILLER_33_260 ();
 sg13g2_decap_8 FILLER_33_267 ();
 sg13g2_fill_2 FILLER_33_274 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_324 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_decap_8 FILLER_33_337 ();
 sg13g2_decap_8 FILLER_33_344 ();
 sg13g2_decap_8 FILLER_33_351 ();
 sg13g2_decap_8 FILLER_33_358 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_fill_2 FILLER_33_379 ();
 sg13g2_fill_1 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_426 ();
 sg13g2_decap_8 FILLER_33_433 ();
 sg13g2_decap_8 FILLER_33_440 ();
 sg13g2_decap_8 FILLER_33_473 ();
 sg13g2_decap_8 FILLER_33_501 ();
 sg13g2_decap_8 FILLER_33_508 ();
 sg13g2_fill_1 FILLER_33_515 ();
 sg13g2_decap_4 FILLER_33_520 ();
 sg13g2_fill_1 FILLER_33_524 ();
 sg13g2_decap_4 FILLER_33_557 ();
 sg13g2_fill_1 FILLER_33_561 ();
 sg13g2_fill_2 FILLER_33_613 ();
 sg13g2_fill_1 FILLER_33_615 ();
 sg13g2_decap_8 FILLER_33_620 ();
 sg13g2_fill_2 FILLER_33_627 ();
 sg13g2_decap_8 FILLER_33_664 ();
 sg13g2_fill_1 FILLER_33_671 ();
 sg13g2_decap_8 FILLER_33_676 ();
 sg13g2_decap_8 FILLER_33_683 ();
 sg13g2_decap_4 FILLER_33_690 ();
 sg13g2_fill_2 FILLER_33_694 ();
 sg13g2_decap_8 FILLER_33_729 ();
 sg13g2_decap_8 FILLER_33_736 ();
 sg13g2_decap_8 FILLER_33_743 ();
 sg13g2_decap_8 FILLER_33_750 ();
 sg13g2_decap_8 FILLER_33_757 ();
 sg13g2_decap_4 FILLER_33_764 ();
 sg13g2_fill_1 FILLER_33_768 ();
 sg13g2_decap_8 FILLER_33_774 ();
 sg13g2_fill_1 FILLER_33_781 ();
 sg13g2_fill_2 FILLER_33_813 ();
 sg13g2_decap_8 FILLER_33_841 ();
 sg13g2_fill_2 FILLER_33_848 ();
 sg13g2_fill_1 FILLER_33_850 ();
 sg13g2_decap_8 FILLER_33_855 ();
 sg13g2_decap_8 FILLER_33_862 ();
 sg13g2_decap_8 FILLER_33_869 ();
 sg13g2_fill_2 FILLER_33_876 ();
 sg13g2_fill_1 FILLER_33_878 ();
 sg13g2_decap_8 FILLER_33_883 ();
 sg13g2_decap_8 FILLER_33_890 ();
 sg13g2_decap_4 FILLER_33_897 ();
 sg13g2_fill_2 FILLER_33_901 ();
 sg13g2_fill_1 FILLER_33_929 ();
 sg13g2_decap_8 FILLER_33_934 ();
 sg13g2_decap_4 FILLER_33_941 ();
 sg13g2_fill_1 FILLER_33_945 ();
 sg13g2_decap_8 FILLER_33_950 ();
 sg13g2_decap_8 FILLER_33_957 ();
 sg13g2_decap_8 FILLER_33_964 ();
 sg13g2_decap_4 FILLER_33_975 ();
 sg13g2_fill_2 FILLER_33_979 ();
 sg13g2_decap_8 FILLER_33_984 ();
 sg13g2_decap_8 FILLER_33_991 ();
 sg13g2_decap_8 FILLER_33_998 ();
 sg13g2_decap_4 FILLER_33_1005 ();
 sg13g2_fill_2 FILLER_33_1009 ();
 sg13g2_decap_8 FILLER_33_1057 ();
 sg13g2_decap_8 FILLER_33_1064 ();
 sg13g2_decap_4 FILLER_33_1101 ();
 sg13g2_fill_2 FILLER_33_1105 ();
 sg13g2_decap_8 FILLER_33_1152 ();
 sg13g2_fill_2 FILLER_33_1159 ();
 sg13g2_fill_1 FILLER_33_1161 ();
 sg13g2_decap_8 FILLER_33_1166 ();
 sg13g2_fill_1 FILLER_33_1173 ();
 sg13g2_decap_8 FILLER_33_1178 ();
 sg13g2_decap_8 FILLER_33_1185 ();
 sg13g2_decap_4 FILLER_33_1192 ();
 sg13g2_fill_1 FILLER_33_1222 ();
 sg13g2_decap_4 FILLER_33_1249 ();
 sg13g2_fill_1 FILLER_33_1253 ();
 sg13g2_decap_4 FILLER_33_1258 ();
 sg13g2_fill_1 FILLER_33_1288 ();
 sg13g2_decap_8 FILLER_33_1314 ();
 sg13g2_decap_8 FILLER_33_1321 ();
 sg13g2_fill_1 FILLER_33_1333 ();
 sg13g2_decap_8 FILLER_33_1364 ();
 sg13g2_fill_1 FILLER_33_1371 ();
 sg13g2_decap_8 FILLER_33_1376 ();
 sg13g2_decap_8 FILLER_33_1383 ();
 sg13g2_fill_1 FILLER_33_1390 ();
 sg13g2_decap_8 FILLER_33_1395 ();
 sg13g2_decap_8 FILLER_33_1402 ();
 sg13g2_fill_2 FILLER_33_1409 ();
 sg13g2_fill_1 FILLER_33_1411 ();
 sg13g2_decap_8 FILLER_33_1441 ();
 sg13g2_decap_8 FILLER_33_1448 ();
 sg13g2_decap_8 FILLER_33_1455 ();
 sg13g2_decap_8 FILLER_33_1462 ();
 sg13g2_decap_8 FILLER_33_1469 ();
 sg13g2_decap_4 FILLER_33_1476 ();
 sg13g2_fill_1 FILLER_33_1553 ();
 sg13g2_decap_8 FILLER_33_1579 ();
 sg13g2_fill_1 FILLER_33_1586 ();
 sg13g2_decap_8 FILLER_33_1591 ();
 sg13g2_decap_8 FILLER_33_1598 ();
 sg13g2_decap_8 FILLER_33_1605 ();
 sg13g2_decap_8 FILLER_33_1612 ();
 sg13g2_decap_4 FILLER_33_1619 ();
 sg13g2_fill_2 FILLER_33_1623 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_254 ();
 sg13g2_decap_4 FILLER_34_261 ();
 sg13g2_fill_2 FILLER_34_265 ();
 sg13g2_decap_8 FILLER_34_271 ();
 sg13g2_decap_4 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_282 ();
 sg13g2_fill_2 FILLER_34_293 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_fill_2 FILLER_34_300 ();
 sg13g2_fill_1 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_324 ();
 sg13g2_decap_4 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_fill_1 FILLER_34_393 ();
 sg13g2_fill_1 FILLER_34_450 ();
 sg13g2_fill_1 FILLER_34_460 ();
 sg13g2_decap_4 FILLER_34_465 ();
 sg13g2_decap_8 FILLER_34_473 ();
 sg13g2_decap_8 FILLER_34_480 ();
 sg13g2_decap_8 FILLER_34_487 ();
 sg13g2_decap_4 FILLER_34_494 ();
 sg13g2_fill_1 FILLER_34_498 ();
 sg13g2_decap_8 FILLER_34_564 ();
 sg13g2_decap_8 FILLER_34_571 ();
 sg13g2_fill_2 FILLER_34_578 ();
 sg13g2_fill_1 FILLER_34_580 ();
 sg13g2_fill_1 FILLER_34_584 ();
 sg13g2_fill_2 FILLER_34_608 ();
 sg13g2_decap_8 FILLER_34_645 ();
 sg13g2_fill_2 FILLER_34_652 ();
 sg13g2_fill_1 FILLER_34_654 ();
 sg13g2_fill_1 FILLER_34_660 ();
 sg13g2_decap_4 FILLER_34_665 ();
 sg13g2_fill_2 FILLER_34_669 ();
 sg13g2_decap_4 FILLER_34_737 ();
 sg13g2_fill_2 FILLER_34_741 ();
 sg13g2_decap_4 FILLER_34_747 ();
 sg13g2_fill_2 FILLER_34_751 ();
 sg13g2_decap_8 FILLER_34_788 ();
 sg13g2_decap_4 FILLER_34_795 ();
 sg13g2_fill_2 FILLER_34_799 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_8 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_840 ();
 sg13g2_fill_1 FILLER_34_847 ();
 sg13g2_decap_8 FILLER_34_856 ();
 sg13g2_decap_8 FILLER_34_863 ();
 sg13g2_fill_2 FILLER_34_870 ();
 sg13g2_decap_8 FILLER_34_898 ();
 sg13g2_decap_4 FILLER_34_965 ();
 sg13g2_fill_1 FILLER_34_969 ();
 sg13g2_decap_8 FILLER_34_974 ();
 sg13g2_decap_8 FILLER_34_981 ();
 sg13g2_decap_4 FILLER_34_988 ();
 sg13g2_decap_4 FILLER_34_997 ();
 sg13g2_fill_2 FILLER_34_1001 ();
 sg13g2_decap_8 FILLER_34_1033 ();
 sg13g2_fill_2 FILLER_34_1040 ();
 sg13g2_decap_8 FILLER_34_1046 ();
 sg13g2_fill_1 FILLER_34_1053 ();
 sg13g2_decap_8 FILLER_34_1058 ();
 sg13g2_decap_8 FILLER_34_1065 ();
 sg13g2_fill_2 FILLER_34_1072 ();
 sg13g2_decap_8 FILLER_34_1115 ();
 sg13g2_decap_8 FILLER_34_1122 ();
 sg13g2_decap_8 FILLER_34_1129 ();
 sg13g2_decap_8 FILLER_34_1136 ();
 sg13g2_decap_4 FILLER_34_1143 ();
 sg13g2_fill_1 FILLER_34_1147 ();
 sg13g2_fill_2 FILLER_34_1157 ();
 sg13g2_fill_1 FILLER_34_1164 ();
 sg13g2_decap_8 FILLER_34_1195 ();
 sg13g2_fill_1 FILLER_34_1202 ();
 sg13g2_decap_8 FILLER_34_1207 ();
 sg13g2_decap_8 FILLER_34_1214 ();
 sg13g2_fill_1 FILLER_34_1221 ();
 sg13g2_decap_8 FILLER_34_1320 ();
 sg13g2_decap_8 FILLER_34_1332 ();
 sg13g2_decap_8 FILLER_34_1339 ();
 sg13g2_decap_8 FILLER_34_1346 ();
 sg13g2_decap_4 FILLER_34_1353 ();
 sg13g2_decap_4 FILLER_34_1362 ();
 sg13g2_decap_8 FILLER_34_1370 ();
 sg13g2_decap_8 FILLER_34_1377 ();
 sg13g2_fill_1 FILLER_34_1384 ();
 sg13g2_decap_8 FILLER_34_1402 ();
 sg13g2_decap_8 FILLER_34_1409 ();
 sg13g2_decap_4 FILLER_34_1416 ();
 sg13g2_fill_2 FILLER_34_1420 ();
 sg13g2_decap_4 FILLER_34_1426 ();
 sg13g2_fill_2 FILLER_34_1430 ();
 sg13g2_decap_8 FILLER_34_1457 ();
 sg13g2_decap_8 FILLER_34_1464 ();
 sg13g2_decap_8 FILLER_34_1471 ();
 sg13g2_decap_4 FILLER_34_1478 ();
 sg13g2_fill_1 FILLER_34_1482 ();
 sg13g2_fill_1 FILLER_34_1509 ();
 sg13g2_decap_4 FILLER_34_1565 ();
 sg13g2_decap_8 FILLER_34_1604 ();
 sg13g2_decap_8 FILLER_34_1611 ();
 sg13g2_decap_8 FILLER_34_1618 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_224 ();
 sg13g2_fill_1 FILLER_35_226 ();
 sg13g2_decap_4 FILLER_35_257 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_315 ();
 sg13g2_decap_4 FILLER_35_363 ();
 sg13g2_fill_2 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_4 FILLER_35_380 ();
 sg13g2_fill_1 FILLER_35_384 ();
 sg13g2_decap_4 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_410 ();
 sg13g2_decap_8 FILLER_35_415 ();
 sg13g2_fill_1 FILLER_35_448 ();
 sg13g2_decap_8 FILLER_35_479 ();
 sg13g2_decap_4 FILLER_35_486 ();
 sg13g2_decap_8 FILLER_35_494 ();
 sg13g2_decap_8 FILLER_35_501 ();
 sg13g2_decap_8 FILLER_35_508 ();
 sg13g2_decap_8 FILLER_35_515 ();
 sg13g2_fill_1 FILLER_35_544 ();
 sg13g2_decap_4 FILLER_35_578 ();
 sg13g2_fill_1 FILLER_35_582 ();
 sg13g2_decap_8 FILLER_35_609 ();
 sg13g2_decap_8 FILLER_35_620 ();
 sg13g2_fill_1 FILLER_35_627 ();
 sg13g2_fill_2 FILLER_35_679 ();
 sg13g2_fill_2 FILLER_35_685 ();
 sg13g2_decap_8 FILLER_35_691 ();
 sg13g2_decap_8 FILLER_35_706 ();
 sg13g2_decap_8 FILLER_35_713 ();
 sg13g2_decap_4 FILLER_35_720 ();
 sg13g2_fill_2 FILLER_35_724 ();
 sg13g2_decap_8 FILLER_35_761 ();
 sg13g2_fill_1 FILLER_35_768 ();
 sg13g2_decap_8 FILLER_35_773 ();
 sg13g2_decap_8 FILLER_35_780 ();
 sg13g2_fill_2 FILLER_35_787 ();
 sg13g2_decap_8 FILLER_35_820 ();
 sg13g2_decap_8 FILLER_35_827 ();
 sg13g2_decap_4 FILLER_35_834 ();
 sg13g2_fill_2 FILLER_35_838 ();
 sg13g2_fill_1 FILLER_35_876 ();
 sg13g2_decap_8 FILLER_35_881 ();
 sg13g2_decap_8 FILLER_35_888 ();
 sg13g2_decap_8 FILLER_35_895 ();
 sg13g2_decap_4 FILLER_35_902 ();
 sg13g2_decap_8 FILLER_35_932 ();
 sg13g2_decap_8 FILLER_35_939 ();
 sg13g2_decap_8 FILLER_35_946 ();
 sg13g2_fill_1 FILLER_35_953 ();
 sg13g2_decap_8 FILLER_35_1014 ();
 sg13g2_decap_8 FILLER_35_1021 ();
 sg13g2_decap_8 FILLER_35_1028 ();
 sg13g2_fill_2 FILLER_35_1035 ();
 sg13g2_decap_8 FILLER_35_1072 ();
 sg13g2_fill_2 FILLER_35_1079 ();
 sg13g2_fill_1 FILLER_35_1081 ();
 sg13g2_fill_2 FILLER_35_1089 ();
 sg13g2_decap_8 FILLER_35_1124 ();
 sg13g2_decap_8 FILLER_35_1131 ();
 sg13g2_fill_2 FILLER_35_1138 ();
 sg13g2_fill_1 FILLER_35_1140 ();
 sg13g2_decap_8 FILLER_35_1201 ();
 sg13g2_decap_8 FILLER_35_1208 ();
 sg13g2_decap_8 FILLER_35_1215 ();
 sg13g2_fill_2 FILLER_35_1299 ();
 sg13g2_fill_1 FILLER_35_1301 ();
 sg13g2_decap_8 FILLER_35_1328 ();
 sg13g2_fill_1 FILLER_35_1335 ();
 sg13g2_fill_1 FILLER_35_1357 ();
 sg13g2_fill_1 FILLER_35_1410 ();
 sg13g2_decap_4 FILLER_35_1416 ();
 sg13g2_fill_2 FILLER_35_1420 ();
 sg13g2_fill_1 FILLER_35_1430 ();
 sg13g2_decap_8 FILLER_35_1457 ();
 sg13g2_decap_8 FILLER_35_1464 ();
 sg13g2_decap_8 FILLER_35_1471 ();
 sg13g2_decap_8 FILLER_35_1478 ();
 sg13g2_fill_2 FILLER_35_1485 ();
 sg13g2_fill_1 FILLER_35_1487 ();
 sg13g2_fill_2 FILLER_35_1525 ();
 sg13g2_fill_1 FILLER_35_1527 ();
 sg13g2_decap_8 FILLER_35_1587 ();
 sg13g2_decap_8 FILLER_35_1594 ();
 sg13g2_decap_8 FILLER_35_1601 ();
 sg13g2_decap_8 FILLER_35_1608 ();
 sg13g2_decap_8 FILLER_35_1615 ();
 sg13g2_fill_2 FILLER_35_1622 ();
 sg13g2_fill_1 FILLER_35_1624 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_4 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_221 ();
 sg13g2_decap_8 FILLER_36_227 ();
 sg13g2_decap_4 FILLER_36_234 ();
 sg13g2_fill_2 FILLER_36_248 ();
 sg13g2_fill_1 FILLER_36_250 ();
 sg13g2_decap_4 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_276 ();
 sg13g2_fill_2 FILLER_36_283 ();
 sg13g2_fill_1 FILLER_36_285 ();
 sg13g2_decap_8 FILLER_36_290 ();
 sg13g2_decap_8 FILLER_36_297 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_4 FILLER_36_315 ();
 sg13g2_decap_4 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_fill_2 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_4 FILLER_36_387 ();
 sg13g2_decap_4 FILLER_36_396 ();
 sg13g2_fill_2 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_fill_1 FILLER_36_430 ();
 sg13g2_decap_8 FILLER_36_435 ();
 sg13g2_decap_4 FILLER_36_442 ();
 sg13g2_fill_1 FILLER_36_446 ();
 sg13g2_fill_2 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_509 ();
 sg13g2_decap_4 FILLER_36_516 ();
 sg13g2_fill_2 FILLER_36_591 ();
 sg13g2_decap_4 FILLER_36_605 ();
 sg13g2_fill_1 FILLER_36_640 ();
 sg13g2_fill_2 FILLER_36_646 ();
 sg13g2_fill_2 FILLER_36_652 ();
 sg13g2_decap_8 FILLER_36_696 ();
 sg13g2_decap_8 FILLER_36_724 ();
 sg13g2_decap_8 FILLER_36_731 ();
 sg13g2_decap_8 FILLER_36_738 ();
 sg13g2_decap_8 FILLER_36_745 ();
 sg13g2_decap_8 FILLER_36_752 ();
 sg13g2_decap_8 FILLER_36_759 ();
 sg13g2_fill_2 FILLER_36_766 ();
 sg13g2_fill_1 FILLER_36_768 ();
 sg13g2_decap_4 FILLER_36_782 ();
 sg13g2_fill_2 FILLER_36_815 ();
 sg13g2_fill_1 FILLER_36_817 ();
 sg13g2_fill_2 FILLER_36_839 ();
 sg13g2_decap_4 FILLER_36_896 ();
 sg13g2_fill_2 FILLER_36_900 ();
 sg13g2_decap_4 FILLER_36_907 ();
 sg13g2_fill_1 FILLER_36_911 ();
 sg13g2_decap_8 FILLER_36_921 ();
 sg13g2_decap_8 FILLER_36_928 ();
 sg13g2_decap_8 FILLER_36_935 ();
 sg13g2_decap_8 FILLER_36_942 ();
 sg13g2_decap_4 FILLER_36_949 ();
 sg13g2_fill_2 FILLER_36_953 ();
 sg13g2_decap_8 FILLER_36_984 ();
 sg13g2_decap_4 FILLER_36_991 ();
 sg13g2_fill_2 FILLER_36_999 ();
 sg13g2_fill_2 FILLER_36_1006 ();
 sg13g2_fill_1 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1013 ();
 sg13g2_decap_4 FILLER_36_1020 ();
 sg13g2_fill_2 FILLER_36_1024 ();
 sg13g2_decap_8 FILLER_36_1039 ();
 sg13g2_fill_2 FILLER_36_1046 ();
 sg13g2_fill_1 FILLER_36_1048 ();
 sg13g2_decap_4 FILLER_36_1087 ();
 sg13g2_fill_1 FILLER_36_1091 ();
 sg13g2_fill_2 FILLER_36_1118 ();
 sg13g2_fill_1 FILLER_36_1120 ();
 sg13g2_fill_1 FILLER_36_1168 ();
 sg13g2_fill_2 FILLER_36_1190 ();
 sg13g2_fill_1 FILLER_36_1192 ();
 sg13g2_fill_2 FILLER_36_1257 ();
 sg13g2_fill_1 FILLER_36_1284 ();
 sg13g2_decap_8 FILLER_36_1289 ();
 sg13g2_decap_4 FILLER_36_1325 ();
 sg13g2_fill_1 FILLER_36_1329 ();
 sg13g2_fill_2 FILLER_36_1335 ();
 sg13g2_fill_1 FILLER_36_1337 ();
 sg13g2_fill_1 FILLER_36_1359 ();
 sg13g2_fill_2 FILLER_36_1364 ();
 sg13g2_fill_2 FILLER_36_1442 ();
 sg13g2_decap_8 FILLER_36_1453 ();
 sg13g2_decap_8 FILLER_36_1460 ();
 sg13g2_decap_8 FILLER_36_1467 ();
 sg13g2_decap_8 FILLER_36_1474 ();
 sg13g2_fill_2 FILLER_36_1481 ();
 sg13g2_fill_1 FILLER_36_1553 ();
 sg13g2_fill_2 FILLER_36_1579 ();
 sg13g2_decap_8 FILLER_36_1606 ();
 sg13g2_decap_8 FILLER_36_1613 ();
 sg13g2_decap_4 FILLER_36_1620 ();
 sg13g2_fill_1 FILLER_36_1624 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_248 ();
 sg13g2_decap_4 FILLER_37_274 ();
 sg13g2_fill_1 FILLER_37_278 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_fill_2 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_404 ();
 sg13g2_decap_8 FILLER_37_411 ();
 sg13g2_fill_2 FILLER_37_418 ();
 sg13g2_decap_8 FILLER_37_425 ();
 sg13g2_fill_1 FILLER_37_432 ();
 sg13g2_decap_8 FILLER_37_437 ();
 sg13g2_fill_2 FILLER_37_444 ();
 sg13g2_fill_1 FILLER_37_446 ();
 sg13g2_fill_2 FILLER_37_473 ();
 sg13g2_decap_8 FILLER_37_484 ();
 sg13g2_decap_8 FILLER_37_491 ();
 sg13g2_decap_4 FILLER_37_498 ();
 sg13g2_decap_8 FILLER_37_619 ();
 sg13g2_decap_8 FILLER_37_626 ();
 sg13g2_fill_2 FILLER_37_633 ();
 sg13g2_fill_2 FILLER_37_639 ();
 sg13g2_fill_1 FILLER_37_641 ();
 sg13g2_decap_8 FILLER_37_668 ();
 sg13g2_fill_2 FILLER_37_701 ();
 sg13g2_fill_1 FILLER_37_703 ();
 sg13g2_decap_8 FILLER_37_725 ();
 sg13g2_fill_1 FILLER_37_732 ();
 sg13g2_decap_4 FILLER_37_754 ();
 sg13g2_fill_1 FILLER_37_789 ();
 sg13g2_fill_2 FILLER_37_816 ();
 sg13g2_fill_1 FILLER_37_839 ();
 sg13g2_decap_8 FILLER_37_871 ();
 sg13g2_decap_8 FILLER_37_878 ();
 sg13g2_decap_4 FILLER_37_885 ();
 sg13g2_fill_2 FILLER_37_889 ();
 sg13g2_decap_4 FILLER_37_912 ();
 sg13g2_decap_8 FILLER_37_958 ();
 sg13g2_decap_4 FILLER_37_965 ();
 sg13g2_decap_8 FILLER_37_1020 ();
 sg13g2_decap_4 FILLER_37_1053 ();
 sg13g2_fill_1 FILLER_37_1057 ();
 sg13g2_decap_8 FILLER_37_1083 ();
 sg13g2_fill_1 FILLER_37_1115 ();
 sg13g2_decap_8 FILLER_37_1121 ();
 sg13g2_fill_1 FILLER_37_1128 ();
 sg13g2_fill_2 FILLER_37_1150 ();
 sg13g2_decap_4 FILLER_37_1224 ();
 sg13g2_fill_2 FILLER_37_1228 ();
 sg13g2_decap_4 FILLER_37_1284 ();
 sg13g2_fill_1 FILLER_37_1288 ();
 sg13g2_fill_2 FILLER_37_1323 ();
 sg13g2_fill_1 FILLER_37_1325 ();
 sg13g2_decap_8 FILLER_37_1330 ();
 sg13g2_decap_8 FILLER_37_1337 ();
 sg13g2_decap_8 FILLER_37_1344 ();
 sg13g2_decap_4 FILLER_37_1351 ();
 sg13g2_fill_2 FILLER_37_1355 ();
 sg13g2_fill_1 FILLER_37_1422 ();
 sg13g2_fill_1 FILLER_37_1427 ();
 sg13g2_decap_8 FILLER_37_1453 ();
 sg13g2_decap_8 FILLER_37_1460 ();
 sg13g2_decap_8 FILLER_37_1467 ();
 sg13g2_fill_2 FILLER_37_1474 ();
 sg13g2_fill_2 FILLER_37_1506 ();
 sg13g2_decap_4 FILLER_37_1559 ();
 sg13g2_fill_1 FILLER_37_1563 ();
 sg13g2_fill_1 FILLER_37_1568 ();
 sg13g2_decap_8 FILLER_37_1600 ();
 sg13g2_decap_8 FILLER_37_1607 ();
 sg13g2_decap_8 FILLER_37_1614 ();
 sg13g2_decap_4 FILLER_37_1621 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_4 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_225 ();
 sg13g2_fill_2 FILLER_38_359 ();
 sg13g2_fill_1 FILLER_38_361 ();
 sg13g2_fill_1 FILLER_38_383 ();
 sg13g2_fill_2 FILLER_38_405 ();
 sg13g2_fill_1 FILLER_38_407 ();
 sg13g2_fill_2 FILLER_38_412 ();
 sg13g2_decap_4 FILLER_38_419 ();
 sg13g2_fill_2 FILLER_38_423 ();
 sg13g2_decap_8 FILLER_38_455 ();
 sg13g2_fill_2 FILLER_38_462 ();
 sg13g2_fill_2 FILLER_38_469 ();
 sg13g2_fill_1 FILLER_38_471 ();
 sg13g2_decap_4 FILLER_38_498 ();
 sg13g2_fill_1 FILLER_38_548 ();
 sg13g2_decap_8 FILLER_38_554 ();
 sg13g2_decap_4 FILLER_38_561 ();
 sg13g2_decap_8 FILLER_38_642 ();
 sg13g2_decap_8 FILLER_38_649 ();
 sg13g2_decap_8 FILLER_38_656 ();
 sg13g2_decap_8 FILLER_38_663 ();
 sg13g2_decap_8 FILLER_38_670 ();
 sg13g2_decap_8 FILLER_38_677 ();
 sg13g2_fill_2 FILLER_38_684 ();
 sg13g2_fill_2 FILLER_38_707 ();
 sg13g2_fill_1 FILLER_38_709 ();
 sg13g2_fill_2 FILLER_38_731 ();
 sg13g2_fill_1 FILLER_38_733 ();
 sg13g2_decap_8 FILLER_38_755 ();
 sg13g2_decap_4 FILLER_38_762 ();
 sg13g2_fill_2 FILLER_38_766 ();
 sg13g2_decap_8 FILLER_38_806 ();
 sg13g2_fill_2 FILLER_38_813 ();
 sg13g2_fill_1 FILLER_38_815 ();
 sg13g2_decap_8 FILLER_38_820 ();
 sg13g2_fill_1 FILLER_38_827 ();
 sg13g2_decap_8 FILLER_38_832 ();
 sg13g2_decap_8 FILLER_38_839 ();
 sg13g2_decap_4 FILLER_38_846 ();
 sg13g2_fill_2 FILLER_38_850 ();
 sg13g2_decap_8 FILLER_38_856 ();
 sg13g2_decap_8 FILLER_38_863 ();
 sg13g2_decap_8 FILLER_38_896 ();
 sg13g2_decap_4 FILLER_38_903 ();
 sg13g2_decap_8 FILLER_38_911 ();
 sg13g2_decap_8 FILLER_38_918 ();
 sg13g2_fill_1 FILLER_38_925 ();
 sg13g2_decap_4 FILLER_38_947 ();
 sg13g2_fill_2 FILLER_38_951 ();
 sg13g2_decap_8 FILLER_38_958 ();
 sg13g2_decap_8 FILLER_38_965 ();
 sg13g2_decap_8 FILLER_38_972 ();
 sg13g2_fill_1 FILLER_38_979 ();
 sg13g2_fill_1 FILLER_38_1030 ();
 sg13g2_decap_8 FILLER_38_1035 ();
 sg13g2_fill_1 FILLER_38_1042 ();
 sg13g2_decap_8 FILLER_38_1048 ();
 sg13g2_fill_1 FILLER_38_1055 ();
 sg13g2_decap_4 FILLER_38_1060 ();
 sg13g2_fill_2 FILLER_38_1078 ();
 sg13g2_fill_2 FILLER_38_1090 ();
 sg13g2_fill_1 FILLER_38_1092 ();
 sg13g2_decap_8 FILLER_38_1097 ();
 sg13g2_decap_8 FILLER_38_1104 ();
 sg13g2_decap_8 FILLER_38_1111 ();
 sg13g2_decap_8 FILLER_38_1118 ();
 sg13g2_fill_2 FILLER_38_1125 ();
 sg13g2_decap_8 FILLER_38_1131 ();
 sg13g2_decap_4 FILLER_38_1138 ();
 sg13g2_decap_8 FILLER_38_1163 ();
 sg13g2_decap_8 FILLER_38_1170 ();
 sg13g2_decap_8 FILLER_38_1177 ();
 sg13g2_decap_8 FILLER_38_1184 ();
 sg13g2_decap_8 FILLER_38_1191 ();
 sg13g2_decap_8 FILLER_38_1198 ();
 sg13g2_fill_1 FILLER_38_1205 ();
 sg13g2_decap_8 FILLER_38_1210 ();
 sg13g2_decap_4 FILLER_38_1217 ();
 sg13g2_decap_4 FILLER_38_1226 ();
 sg13g2_fill_2 FILLER_38_1234 ();
 sg13g2_decap_8 FILLER_38_1272 ();
 sg13g2_fill_1 FILLER_38_1279 ();
 sg13g2_fill_2 FILLER_38_1310 ();
 sg13g2_decap_8 FILLER_38_1343 ();
 sg13g2_decap_4 FILLER_38_1350 ();
 sg13g2_fill_1 FILLER_38_1432 ();
 sg13g2_fill_2 FILLER_38_1437 ();
 sg13g2_fill_1 FILLER_38_1439 ();
 sg13g2_fill_2 FILLER_38_1482 ();
 sg13g2_fill_1 FILLER_38_1539 ();
 sg13g2_decap_8 FILLER_38_1599 ();
 sg13g2_decap_8 FILLER_38_1606 ();
 sg13g2_decap_8 FILLER_38_1613 ();
 sg13g2_decap_4 FILLER_38_1620 ();
 sg13g2_fill_1 FILLER_38_1624 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_4 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_183 ();
 sg13g2_decap_8 FILLER_39_190 ();
 sg13g2_decap_8 FILLER_39_197 ();
 sg13g2_decap_8 FILLER_39_204 ();
 sg13g2_decap_4 FILLER_39_211 ();
 sg13g2_fill_1 FILLER_39_274 ();
 sg13g2_fill_1 FILLER_39_288 ();
 sg13g2_decap_8 FILLER_39_331 ();
 sg13g2_decap_8 FILLER_39_338 ();
 sg13g2_decap_8 FILLER_39_345 ();
 sg13g2_decap_8 FILLER_39_352 ();
 sg13g2_decap_8 FILLER_39_359 ();
 sg13g2_decap_8 FILLER_39_366 ();
 sg13g2_fill_2 FILLER_39_373 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_fill_1 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_426 ();
 sg13g2_decap_4 FILLER_39_433 ();
 sg13g2_fill_2 FILLER_39_437 ();
 sg13g2_decap_8 FILLER_39_444 ();
 sg13g2_decap_8 FILLER_39_451 ();
 sg13g2_decap_8 FILLER_39_458 ();
 sg13g2_decap_4 FILLER_39_465 ();
 sg13g2_fill_1 FILLER_39_469 ();
 sg13g2_decap_4 FILLER_39_473 ();
 sg13g2_decap_8 FILLER_39_486 ();
 sg13g2_decap_8 FILLER_39_493 ();
 sg13g2_fill_2 FILLER_39_500 ();
 sg13g2_fill_2 FILLER_39_512 ();
 sg13g2_fill_1 FILLER_39_514 ();
 sg13g2_fill_2 FILLER_39_524 ();
 sg13g2_fill_1 FILLER_39_526 ();
 sg13g2_decap_8 FILLER_39_565 ();
 sg13g2_decap_4 FILLER_39_572 ();
 sg13g2_fill_2 FILLER_39_597 ();
 sg13g2_fill_1 FILLER_39_599 ();
 sg13g2_decap_4 FILLER_39_634 ();
 sg13g2_fill_1 FILLER_39_638 ();
 sg13g2_decap_8 FILLER_39_681 ();
 sg13g2_decap_8 FILLER_39_688 ();
 sg13g2_decap_8 FILLER_39_695 ();
 sg13g2_decap_8 FILLER_39_712 ();
 sg13g2_decap_8 FILLER_39_719 ();
 sg13g2_decap_8 FILLER_39_726 ();
 sg13g2_decap_8 FILLER_39_733 ();
 sg13g2_fill_2 FILLER_39_749 ();
 sg13g2_decap_8 FILLER_39_755 ();
 sg13g2_decap_8 FILLER_39_762 ();
 sg13g2_decap_8 FILLER_39_769 ();
 sg13g2_fill_1 FILLER_39_776 ();
 sg13g2_fill_2 FILLER_39_786 ();
 sg13g2_decap_4 FILLER_39_793 ();
 sg13g2_fill_2 FILLER_39_801 ();
 sg13g2_fill_1 FILLER_39_803 ();
 sg13g2_fill_1 FILLER_39_835 ();
 sg13g2_decap_4 FILLER_39_841 ();
 sg13g2_fill_1 FILLER_39_845 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_fill_2 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_39_868 ();
 sg13g2_decap_4 FILLER_39_875 ();
 sg13g2_decap_8 FILLER_39_883 ();
 sg13g2_fill_2 FILLER_39_890 ();
 sg13g2_fill_1 FILLER_39_936 ();
 sg13g2_decap_8 FILLER_39_941 ();
 sg13g2_decap_8 FILLER_39_948 ();
 sg13g2_decap_8 FILLER_39_955 ();
 sg13g2_fill_1 FILLER_39_962 ();
 sg13g2_decap_8 FILLER_39_968 ();
 sg13g2_decap_8 FILLER_39_975 ();
 sg13g2_decap_8 FILLER_39_982 ();
 sg13g2_decap_8 FILLER_39_989 ();
 sg13g2_decap_4 FILLER_39_996 ();
 sg13g2_fill_2 FILLER_39_1000 ();
 sg13g2_decap_8 FILLER_39_1006 ();
 sg13g2_decap_4 FILLER_39_1013 ();
 sg13g2_fill_2 FILLER_39_1017 ();
 sg13g2_decap_8 FILLER_39_1079 ();
 sg13g2_fill_1 FILLER_39_1086 ();
 sg13g2_fill_1 FILLER_39_1118 ();
 sg13g2_decap_8 FILLER_39_1145 ();
 sg13g2_decap_8 FILLER_39_1152 ();
 sg13g2_decap_4 FILLER_39_1159 ();
 sg13g2_fill_1 FILLER_39_1163 ();
 sg13g2_decap_8 FILLER_39_1185 ();
 sg13g2_decap_8 FILLER_39_1192 ();
 sg13g2_fill_2 FILLER_39_1199 ();
 sg13g2_decap_8 FILLER_39_1205 ();
 sg13g2_decap_4 FILLER_39_1212 ();
 sg13g2_fill_2 FILLER_39_1216 ();
 sg13g2_decap_8 FILLER_39_1258 ();
 sg13g2_decap_4 FILLER_39_1265 ();
 sg13g2_decap_8 FILLER_39_1290 ();
 sg13g2_decap_4 FILLER_39_1297 ();
 sg13g2_decap_4 FILLER_39_1310 ();
 sg13g2_decap_8 FILLER_39_1318 ();
 sg13g2_decap_8 FILLER_39_1325 ();
 sg13g2_fill_2 FILLER_39_1332 ();
 sg13g2_fill_1 FILLER_39_1338 ();
 sg13g2_fill_1 FILLER_39_1348 ();
 sg13g2_fill_1 FILLER_39_1416 ();
 sg13g2_decap_8 FILLER_39_1464 ();
 sg13g2_decap_8 FILLER_39_1471 ();
 sg13g2_decap_4 FILLER_39_1478 ();
 sg13g2_fill_2 FILLER_39_1482 ();
 sg13g2_fill_1 FILLER_39_1492 ();
 sg13g2_fill_1 FILLER_39_1497 ();
 sg13g2_decap_8 FILLER_39_1599 ();
 sg13g2_decap_8 FILLER_39_1606 ();
 sg13g2_decap_8 FILLER_39_1613 ();
 sg13g2_decap_4 FILLER_39_1620 ();
 sg13g2_fill_1 FILLER_39_1624 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_4 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_198 ();
 sg13g2_decap_8 FILLER_40_205 ();
 sg13g2_decap_4 FILLER_40_212 ();
 sg13g2_fill_2 FILLER_40_216 ();
 sg13g2_decap_8 FILLER_40_225 ();
 sg13g2_fill_1 FILLER_40_232 ();
 sg13g2_fill_2 FILLER_40_288 ();
 sg13g2_decap_8 FILLER_40_326 ();
 sg13g2_decap_4 FILLER_40_333 ();
 sg13g2_fill_1 FILLER_40_337 ();
 sg13g2_fill_1 FILLER_40_342 ();
 sg13g2_fill_2 FILLER_40_356 ();
 sg13g2_decap_8 FILLER_40_363 ();
 sg13g2_decap_4 FILLER_40_370 ();
 sg13g2_fill_2 FILLER_40_374 ();
 sg13g2_fill_2 FILLER_40_385 ();
 sg13g2_decap_4 FILLER_40_391 ();
 sg13g2_fill_1 FILLER_40_395 ();
 sg13g2_decap_8 FILLER_40_405 ();
 sg13g2_fill_1 FILLER_40_412 ();
 sg13g2_decap_8 FILLER_40_426 ();
 sg13g2_decap_4 FILLER_40_433 ();
 sg13g2_fill_1 FILLER_40_437 ();
 sg13g2_decap_8 FILLER_40_442 ();
 sg13g2_decap_8 FILLER_40_449 ();
 sg13g2_fill_2 FILLER_40_456 ();
 sg13g2_fill_1 FILLER_40_458 ();
 sg13g2_fill_1 FILLER_40_464 ();
 sg13g2_fill_1 FILLER_40_469 ();
 sg13g2_decap_4 FILLER_40_495 ();
 sg13g2_fill_2 FILLER_40_499 ();
 sg13g2_decap_8 FILLER_40_509 ();
 sg13g2_decap_4 FILLER_40_516 ();
 sg13g2_fill_1 FILLER_40_520 ();
 sg13g2_fill_1 FILLER_40_547 ();
 sg13g2_decap_4 FILLER_40_569 ();
 sg13g2_fill_1 FILLER_40_619 ();
 sg13g2_fill_1 FILLER_40_641 ();
 sg13g2_fill_1 FILLER_40_663 ();
 sg13g2_decap_8 FILLER_40_685 ();
 sg13g2_decap_8 FILLER_40_692 ();
 sg13g2_decap_8 FILLER_40_699 ();
 sg13g2_decap_8 FILLER_40_706 ();
 sg13g2_decap_8 FILLER_40_717 ();
 sg13g2_fill_2 FILLER_40_724 ();
 sg13g2_fill_1 FILLER_40_726 ();
 sg13g2_decap_4 FILLER_40_737 ();
 sg13g2_fill_2 FILLER_40_741 ();
 sg13g2_fill_2 FILLER_40_769 ();
 sg13g2_fill_1 FILLER_40_771 ();
 sg13g2_decap_4 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_807 ();
 sg13g2_decap_8 FILLER_40_814 ();
 sg13g2_decap_8 FILLER_40_821 ();
 sg13g2_fill_1 FILLER_40_828 ();
 sg13g2_decap_4 FILLER_40_834 ();
 sg13g2_fill_1 FILLER_40_838 ();
 sg13g2_decap_4 FILLER_40_891 ();
 sg13g2_fill_1 FILLER_40_895 ();
 sg13g2_fill_2 FILLER_40_906 ();
 sg13g2_decap_4 FILLER_40_921 ();
 sg13g2_fill_1 FILLER_40_925 ();
 sg13g2_decap_4 FILLER_40_952 ();
 sg13g2_fill_1 FILLER_40_956 ();
 sg13g2_decap_8 FILLER_40_975 ();
 sg13g2_decap_8 FILLER_40_982 ();
 sg13g2_fill_2 FILLER_40_989 ();
 sg13g2_fill_1 FILLER_40_991 ();
 sg13g2_fill_2 FILLER_40_1001 ();
 sg13g2_fill_1 FILLER_40_1003 ();
 sg13g2_decap_4 FILLER_40_1008 ();
 sg13g2_fill_2 FILLER_40_1012 ();
 sg13g2_fill_2 FILLER_40_1049 ();
 sg13g2_decap_8 FILLER_40_1060 ();
 sg13g2_decap_8 FILLER_40_1067 ();
 sg13g2_decap_8 FILLER_40_1074 ();
 sg13g2_fill_1 FILLER_40_1081 ();
 sg13g2_fill_2 FILLER_40_1119 ();
 sg13g2_fill_1 FILLER_40_1121 ();
 sg13g2_decap_8 FILLER_40_1131 ();
 sg13g2_decap_8 FILLER_40_1138 ();
 sg13g2_fill_2 FILLER_40_1145 ();
 sg13g2_fill_2 FILLER_40_1151 ();
 sg13g2_fill_2 FILLER_40_1162 ();
 sg13g2_decap_4 FILLER_40_1220 ();
 sg13g2_decap_4 FILLER_40_1262 ();
 sg13g2_fill_1 FILLER_40_1266 ();
 sg13g2_decap_8 FILLER_40_1288 ();
 sg13g2_fill_2 FILLER_40_1321 ();
 sg13g2_decap_8 FILLER_40_1449 ();
 sg13g2_decap_8 FILLER_40_1456 ();
 sg13g2_decap_8 FILLER_40_1463 ();
 sg13g2_decap_8 FILLER_40_1470 ();
 sg13g2_fill_2 FILLER_40_1477 ();
 sg13g2_fill_1 FILLER_40_1479 ();
 sg13g2_fill_2 FILLER_40_1566 ();
 sg13g2_decap_8 FILLER_40_1573 ();
 sg13g2_decap_8 FILLER_40_1580 ();
 sg13g2_decap_8 FILLER_40_1587 ();
 sg13g2_decap_8 FILLER_40_1594 ();
 sg13g2_decap_8 FILLER_40_1601 ();
 sg13g2_decap_8 FILLER_40_1608 ();
 sg13g2_decap_8 FILLER_40_1615 ();
 sg13g2_fill_2 FILLER_40_1622 ();
 sg13g2_fill_1 FILLER_40_1624 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_4 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_201 ();
 sg13g2_decap_4 FILLER_41_208 ();
 sg13g2_fill_1 FILLER_41_293 ();
 sg13g2_fill_2 FILLER_41_319 ();
 sg13g2_decap_4 FILLER_41_403 ();
 sg13g2_decap_4 FILLER_41_484 ();
 sg13g2_fill_1 FILLER_41_488 ();
 sg13g2_fill_2 FILLER_41_520 ();
 sg13g2_fill_1 FILLER_41_522 ();
 sg13g2_fill_2 FILLER_41_579 ();
 sg13g2_fill_1 FILLER_41_581 ();
 sg13g2_decap_8 FILLER_41_586 ();
 sg13g2_decap_4 FILLER_41_593 ();
 sg13g2_fill_2 FILLER_41_597 ();
 sg13g2_decap_8 FILLER_41_629 ();
 sg13g2_decap_8 FILLER_41_636 ();
 sg13g2_decap_8 FILLER_41_643 ();
 sg13g2_decap_8 FILLER_41_650 ();
 sg13g2_decap_8 FILLER_41_657 ();
 sg13g2_decap_8 FILLER_41_664 ();
 sg13g2_decap_8 FILLER_41_671 ();
 sg13g2_decap_8 FILLER_41_678 ();
 sg13g2_fill_2 FILLER_41_685 ();
 sg13g2_decap_8 FILLER_41_692 ();
 sg13g2_fill_2 FILLER_41_699 ();
 sg13g2_fill_1 FILLER_41_705 ();
 sg13g2_decap_8 FILLER_41_732 ();
 sg13g2_decap_8 FILLER_41_739 ();
 sg13g2_decap_8 FILLER_41_746 ();
 sg13g2_fill_1 FILLER_41_753 ();
 sg13g2_decap_8 FILLER_41_757 ();
 sg13g2_decap_8 FILLER_41_764 ();
 sg13g2_decap_8 FILLER_41_776 ();
 sg13g2_decap_4 FILLER_41_783 ();
 sg13g2_fill_2 FILLER_41_787 ();
 sg13g2_decap_8 FILLER_41_793 ();
 sg13g2_decap_8 FILLER_41_800 ();
 sg13g2_decap_4 FILLER_41_807 ();
 sg13g2_fill_1 FILLER_41_811 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_4 FILLER_41_847 ();
 sg13g2_fill_1 FILLER_41_851 ();
 sg13g2_fill_2 FILLER_41_856 ();
 sg13g2_decap_8 FILLER_41_863 ();
 sg13g2_fill_2 FILLER_41_870 ();
 sg13g2_decap_8 FILLER_41_876 ();
 sg13g2_decap_8 FILLER_41_883 ();
 sg13g2_decap_8 FILLER_41_890 ();
 sg13g2_decap_8 FILLER_41_897 ();
 sg13g2_decap_8 FILLER_41_904 ();
 sg13g2_fill_2 FILLER_41_911 ();
 sg13g2_decap_8 FILLER_41_943 ();
 sg13g2_decap_8 FILLER_41_950 ();
 sg13g2_decap_4 FILLER_41_957 ();
 sg13g2_fill_2 FILLER_41_961 ();
 sg13g2_fill_2 FILLER_41_989 ();
 sg13g2_decap_8 FILLER_41_1022 ();
 sg13g2_decap_8 FILLER_41_1029 ();
 sg13g2_decap_8 FILLER_41_1036 ();
 sg13g2_fill_1 FILLER_41_1043 ();
 sg13g2_decap_8 FILLER_41_1069 ();
 sg13g2_fill_1 FILLER_41_1120 ();
 sg13g2_decap_8 FILLER_41_1125 ();
 sg13g2_fill_1 FILLER_41_1132 ();
 sg13g2_fill_2 FILLER_41_1138 ();
 sg13g2_decap_8 FILLER_41_1166 ();
 sg13g2_decap_8 FILLER_41_1173 ();
 sg13g2_decap_4 FILLER_41_1180 ();
 sg13g2_decap_4 FILLER_41_1238 ();
 sg13g2_fill_1 FILLER_41_1310 ();
 sg13g2_fill_2 FILLER_41_1363 ();
 sg13g2_fill_2 FILLER_41_1416 ();
 sg13g2_decap_8 FILLER_41_1447 ();
 sg13g2_decap_8 FILLER_41_1454 ();
 sg13g2_fill_2 FILLER_41_1461 ();
 sg13g2_fill_2 FILLER_41_1484 ();
 sg13g2_fill_1 FILLER_41_1486 ();
 sg13g2_decap_4 FILLER_41_1491 ();
 sg13g2_fill_2 FILLER_41_1495 ();
 sg13g2_fill_2 FILLER_41_1543 ();
 sg13g2_decap_8 FILLER_41_1575 ();
 sg13g2_decap_8 FILLER_41_1582 ();
 sg13g2_decap_8 FILLER_41_1589 ();
 sg13g2_decap_8 FILLER_41_1596 ();
 sg13g2_decap_8 FILLER_41_1603 ();
 sg13g2_decap_8 FILLER_41_1610 ();
 sg13g2_decap_8 FILLER_41_1617 ();
 sg13g2_fill_1 FILLER_41_1624 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_fill_2 FILLER_42_168 ();
 sg13g2_fill_1 FILLER_42_170 ();
 sg13g2_decap_8 FILLER_42_197 ();
 sg13g2_decap_4 FILLER_42_208 ();
 sg13g2_fill_2 FILLER_42_212 ();
 sg13g2_fill_2 FILLER_42_240 ();
 sg13g2_fill_1 FILLER_42_242 ();
 sg13g2_fill_2 FILLER_42_247 ();
 sg13g2_fill_2 FILLER_42_254 ();
 sg13g2_decap_4 FILLER_42_260 ();
 sg13g2_fill_2 FILLER_42_320 ();
 sg13g2_fill_1 FILLER_42_327 ();
 sg13g2_fill_1 FILLER_42_332 ();
 sg13g2_fill_1 FILLER_42_437 ();
 sg13g2_fill_1 FILLER_42_447 ();
 sg13g2_decap_8 FILLER_42_452 ();
 sg13g2_decap_4 FILLER_42_459 ();
 sg13g2_fill_2 FILLER_42_467 ();
 sg13g2_decap_8 FILLER_42_482 ();
 sg13g2_decap_4 FILLER_42_489 ();
 sg13g2_fill_1 FILLER_42_523 ();
 sg13g2_fill_2 FILLER_42_561 ();
 sg13g2_fill_1 FILLER_42_572 ();
 sg13g2_fill_2 FILLER_42_624 ();
 sg13g2_fill_1 FILLER_42_626 ();
 sg13g2_decap_8 FILLER_42_648 ();
 sg13g2_fill_2 FILLER_42_655 ();
 sg13g2_fill_1 FILLER_42_657 ();
 sg13g2_decap_8 FILLER_42_662 ();
 sg13g2_decap_8 FILLER_42_669 ();
 sg13g2_decap_8 FILLER_42_676 ();
 sg13g2_decap_4 FILLER_42_683 ();
 sg13g2_decap_8 FILLER_42_726 ();
 sg13g2_decap_8 FILLER_42_733 ();
 sg13g2_decap_4 FILLER_42_740 ();
 sg13g2_fill_1 FILLER_42_744 ();
 sg13g2_decap_8 FILLER_42_783 ();
 sg13g2_fill_1 FILLER_42_790 ();
 sg13g2_fill_1 FILLER_42_801 ();
 sg13g2_decap_8 FILLER_42_831 ();
 sg13g2_fill_2 FILLER_42_838 ();
 sg13g2_fill_1 FILLER_42_840 ();
 sg13g2_decap_4 FILLER_42_871 ();
 sg13g2_fill_2 FILLER_42_875 ();
 sg13g2_decap_4 FILLER_42_882 ();
 sg13g2_fill_2 FILLER_42_886 ();
 sg13g2_decap_8 FILLER_42_898 ();
 sg13g2_decap_4 FILLER_42_926 ();
 sg13g2_fill_2 FILLER_42_930 ();
 sg13g2_fill_2 FILLER_42_953 ();
 sg13g2_fill_2 FILLER_42_960 ();
 sg13g2_decap_8 FILLER_42_972 ();
 sg13g2_fill_2 FILLER_42_979 ();
 sg13g2_fill_1 FILLER_42_981 ();
 sg13g2_decap_4 FILLER_42_987 ();
 sg13g2_fill_1 FILLER_42_991 ();
 sg13g2_decap_8 FILLER_42_1001 ();
 sg13g2_decap_8 FILLER_42_1008 ();
 sg13g2_decap_8 FILLER_42_1015 ();
 sg13g2_decap_8 FILLER_42_1026 ();
 sg13g2_decap_8 FILLER_42_1072 ();
 sg13g2_fill_1 FILLER_42_1079 ();
 sg13g2_decap_8 FILLER_42_1084 ();
 sg13g2_decap_4 FILLER_42_1091 ();
 sg13g2_fill_2 FILLER_42_1099 ();
 sg13g2_decap_8 FILLER_42_1137 ();
 sg13g2_fill_2 FILLER_42_1144 ();
 sg13g2_fill_2 FILLER_42_1151 ();
 sg13g2_fill_1 FILLER_42_1163 ();
 sg13g2_fill_2 FILLER_42_1168 ();
 sg13g2_fill_1 FILLER_42_1174 ();
 sg13g2_fill_2 FILLER_42_1216 ();
 sg13g2_decap_8 FILLER_42_1273 ();
 sg13g2_decap_8 FILLER_42_1280 ();
 sg13g2_decap_8 FILLER_42_1287 ();
 sg13g2_decap_4 FILLER_42_1294 ();
 sg13g2_fill_1 FILLER_42_1298 ();
 sg13g2_decap_8 FILLER_42_1304 ();
 sg13g2_decap_4 FILLER_42_1311 ();
 sg13g2_decap_8 FILLER_42_1336 ();
 sg13g2_decap_8 FILLER_42_1343 ();
 sg13g2_decap_4 FILLER_42_1350 ();
 sg13g2_fill_2 FILLER_42_1354 ();
 sg13g2_fill_2 FILLER_42_1361 ();
 sg13g2_decap_8 FILLER_42_1410 ();
 sg13g2_decap_4 FILLER_42_1417 ();
 sg13g2_fill_2 FILLER_42_1421 ();
 sg13g2_decap_4 FILLER_42_1432 ();
 sg13g2_decap_8 FILLER_42_1440 ();
 sg13g2_decap_4 FILLER_42_1447 ();
 sg13g2_decap_8 FILLER_42_1472 ();
 sg13g2_decap_4 FILLER_42_1479 ();
 sg13g2_decap_8 FILLER_42_1488 ();
 sg13g2_fill_2 FILLER_42_1499 ();
 sg13g2_fill_1 FILLER_42_1501 ();
 sg13g2_decap_8 FILLER_42_1528 ();
 sg13g2_fill_1 FILLER_42_1539 ();
 sg13g2_decap_8 FILLER_42_1570 ();
 sg13g2_decap_8 FILLER_42_1577 ();
 sg13g2_decap_8 FILLER_42_1584 ();
 sg13g2_decap_8 FILLER_42_1591 ();
 sg13g2_decap_8 FILLER_42_1598 ();
 sg13g2_decap_8 FILLER_42_1605 ();
 sg13g2_decap_8 FILLER_42_1612 ();
 sg13g2_decap_4 FILLER_42_1619 ();
 sg13g2_fill_2 FILLER_42_1623 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_fill_1 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_159 ();
 sg13g2_decap_8 FILLER_43_166 ();
 sg13g2_decap_4 FILLER_43_173 ();
 sg13g2_fill_2 FILLER_43_177 ();
 sg13g2_decap_4 FILLER_43_184 ();
 sg13g2_decap_4 FILLER_43_192 ();
 sg13g2_fill_1 FILLER_43_196 ();
 sg13g2_fill_2 FILLER_43_228 ();
 sg13g2_fill_1 FILLER_43_230 ();
 sg13g2_fill_2 FILLER_43_285 ();
 sg13g2_fill_1 FILLER_43_321 ();
 sg13g2_decap_4 FILLER_43_327 ();
 sg13g2_fill_2 FILLER_43_335 ();
 sg13g2_fill_1 FILLER_43_337 ();
 sg13g2_decap_8 FILLER_43_418 ();
 sg13g2_decap_8 FILLER_43_425 ();
 sg13g2_decap_8 FILLER_43_432 ();
 sg13g2_fill_2 FILLER_43_439 ();
 sg13g2_fill_2 FILLER_43_466 ();
 sg13g2_fill_1 FILLER_43_468 ();
 sg13g2_fill_2 FILLER_43_495 ();
 sg13g2_decap_4 FILLER_43_527 ();
 sg13g2_fill_2 FILLER_43_531 ();
 sg13g2_decap_4 FILLER_43_559 ();
 sg13g2_fill_2 FILLER_43_563 ();
 sg13g2_decap_4 FILLER_43_593 ();
 sg13g2_decap_4 FILLER_43_610 ();
 sg13g2_fill_2 FILLER_43_614 ();
 sg13g2_fill_2 FILLER_43_624 ();
 sg13g2_decap_8 FILLER_43_647 ();
 sg13g2_decap_8 FILLER_43_680 ();
 sg13g2_fill_1 FILLER_43_738 ();
 sg13g2_fill_1 FILLER_43_843 ();
 sg13g2_decap_4 FILLER_43_870 ();
 sg13g2_fill_1 FILLER_43_874 ();
 sg13g2_decap_8 FILLER_43_880 ();
 sg13g2_decap_4 FILLER_43_887 ();
 sg13g2_fill_2 FILLER_43_891 ();
 sg13g2_fill_1 FILLER_43_918 ();
 sg13g2_fill_1 FILLER_43_924 ();
 sg13g2_fill_2 FILLER_43_929 ();
 sg13g2_fill_1 FILLER_43_931 ();
 sg13g2_decap_8 FILLER_43_957 ();
 sg13g2_fill_2 FILLER_43_964 ();
 sg13g2_decap_8 FILLER_43_970 ();
 sg13g2_decap_8 FILLER_43_977 ();
 sg13g2_fill_1 FILLER_43_984 ();
 sg13g2_fill_2 FILLER_43_1070 ();
 sg13g2_fill_1 FILLER_43_1077 ();
 sg13g2_fill_1 FILLER_43_1103 ();
 sg13g2_decap_8 FILLER_43_1129 ();
 sg13g2_decap_8 FILLER_43_1136 ();
 sg13g2_fill_1 FILLER_43_1143 ();
 sg13g2_fill_1 FILLER_43_1149 ();
 sg13g2_decap_8 FILLER_43_1175 ();
 sg13g2_decap_8 FILLER_43_1182 ();
 sg13g2_fill_2 FILLER_43_1189 ();
 sg13g2_fill_1 FILLER_43_1191 ();
 sg13g2_decap_4 FILLER_43_1226 ();
 sg13g2_decap_8 FILLER_43_1276 ();
 sg13g2_decap_8 FILLER_43_1283 ();
 sg13g2_decap_8 FILLER_43_1290 ();
 sg13g2_decap_8 FILLER_43_1297 ();
 sg13g2_decap_8 FILLER_43_1304 ();
 sg13g2_decap_8 FILLER_43_1311 ();
 sg13g2_fill_2 FILLER_43_1318 ();
 sg13g2_fill_1 FILLER_43_1320 ();
 sg13g2_decap_8 FILLER_43_1326 ();
 sg13g2_decap_4 FILLER_43_1333 ();
 sg13g2_decap_8 FILLER_43_1342 ();
 sg13g2_decap_4 FILLER_43_1366 ();
 sg13g2_fill_2 FILLER_43_1395 ();
 sg13g2_fill_1 FILLER_43_1397 ();
 sg13g2_decap_8 FILLER_43_1419 ();
 sg13g2_fill_1 FILLER_43_1426 ();
 sg13g2_decap_8 FILLER_43_1432 ();
 sg13g2_fill_2 FILLER_43_1439 ();
 sg13g2_fill_1 FILLER_43_1441 ();
 sg13g2_fill_2 FILLER_43_1446 ();
 sg13g2_fill_1 FILLER_43_1448 ();
 sg13g2_decap_8 FILLER_43_1470 ();
 sg13g2_fill_2 FILLER_43_1477 ();
 sg13g2_decap_4 FILLER_43_1526 ();
 sg13g2_decap_8 FILLER_43_1534 ();
 sg13g2_fill_1 FILLER_43_1541 ();
 sg13g2_fill_2 FILLER_43_1546 ();
 sg13g2_fill_1 FILLER_43_1548 ();
 sg13g2_decap_8 FILLER_43_1591 ();
 sg13g2_decap_8 FILLER_43_1598 ();
 sg13g2_decap_8 FILLER_43_1605 ();
 sg13g2_decap_8 FILLER_43_1612 ();
 sg13g2_decap_4 FILLER_43_1619 ();
 sg13g2_fill_2 FILLER_43_1623 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_fill_2 FILLER_44_147 ();
 sg13g2_fill_2 FILLER_44_175 ();
 sg13g2_fill_1 FILLER_44_177 ();
 sg13g2_decap_8 FILLER_44_199 ();
 sg13g2_decap_4 FILLER_44_206 ();
 sg13g2_fill_1 FILLER_44_210 ();
 sg13g2_fill_2 FILLER_44_216 ();
 sg13g2_fill_2 FILLER_44_222 ();
 sg13g2_decap_4 FILLER_44_228 ();
 sg13g2_decap_8 FILLER_44_263 ();
 sg13g2_decap_8 FILLER_44_270 ();
 sg13g2_decap_4 FILLER_44_277 ();
 sg13g2_fill_2 FILLER_44_337 ();
 sg13g2_fill_1 FILLER_44_339 ();
 sg13g2_fill_1 FILLER_44_365 ();
 sg13g2_fill_2 FILLER_44_439 ();
 sg13g2_decap_8 FILLER_44_467 ();
 sg13g2_decap_8 FILLER_44_474 ();
 sg13g2_decap_8 FILLER_44_481 ();
 sg13g2_decap_8 FILLER_44_488 ();
 sg13g2_fill_2 FILLER_44_495 ();
 sg13g2_decap_8 FILLER_44_528 ();
 sg13g2_fill_2 FILLER_44_535 ();
 sg13g2_fill_1 FILLER_44_537 ();
 sg13g2_decap_8 FILLER_44_542 ();
 sg13g2_decap_8 FILLER_44_549 ();
 sg13g2_fill_1 FILLER_44_556 ();
 sg13g2_fill_1 FILLER_44_566 ();
 sg13g2_decap_8 FILLER_44_571 ();
 sg13g2_decap_4 FILLER_44_583 ();
 sg13g2_fill_2 FILLER_44_592 ();
 sg13g2_fill_1 FILLER_44_599 ();
 sg13g2_decap_4 FILLER_44_626 ();
 sg13g2_fill_1 FILLER_44_630 ();
 sg13g2_decap_8 FILLER_44_640 ();
 sg13g2_decap_8 FILLER_44_647 ();
 sg13g2_fill_2 FILLER_44_659 ();
 sg13g2_fill_1 FILLER_44_661 ();
 sg13g2_decap_8 FILLER_44_666 ();
 sg13g2_decap_8 FILLER_44_673 ();
 sg13g2_decap_8 FILLER_44_680 ();
 sg13g2_decap_8 FILLER_44_687 ();
 sg13g2_decap_4 FILLER_44_710 ();
 sg13g2_fill_1 FILLER_44_714 ();
 sg13g2_fill_2 FILLER_44_736 ();
 sg13g2_fill_1 FILLER_44_738 ();
 sg13g2_decap_8 FILLER_44_744 ();
 sg13g2_decap_4 FILLER_44_751 ();
 sg13g2_decap_8 FILLER_44_763 ();
 sg13g2_decap_4 FILLER_44_770 ();
 sg13g2_decap_4 FILLER_44_778 ();
 sg13g2_fill_2 FILLER_44_782 ();
 sg13g2_decap_8 FILLER_44_809 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_decap_4 FILLER_44_823 ();
 sg13g2_fill_1 FILLER_44_827 ();
 sg13g2_fill_2 FILLER_44_833 ();
 sg13g2_fill_1 FILLER_44_840 ();
 sg13g2_fill_2 FILLER_44_846 ();
 sg13g2_fill_1 FILLER_44_848 ();
 sg13g2_decap_8 FILLER_44_853 ();
 sg13g2_fill_2 FILLER_44_860 ();
 sg13g2_fill_1 FILLER_44_862 ();
 sg13g2_decap_4 FILLER_44_868 ();
 sg13g2_decap_8 FILLER_44_897 ();
 sg13g2_fill_2 FILLER_44_904 ();
 sg13g2_fill_1 FILLER_44_906 ();
 sg13g2_decap_8 FILLER_44_933 ();
 sg13g2_fill_1 FILLER_44_940 ();
 sg13g2_decap_8 FILLER_44_946 ();
 sg13g2_fill_2 FILLER_44_984 ();
 sg13g2_fill_2 FILLER_44_1017 ();
 sg13g2_fill_2 FILLER_44_1023 ();
 sg13g2_fill_1 FILLER_44_1025 ();
 sg13g2_decap_4 FILLER_44_1137 ();
 sg13g2_decap_8 FILLER_44_1177 ();
 sg13g2_fill_2 FILLER_44_1184 ();
 sg13g2_fill_1 FILLER_44_1186 ();
 sg13g2_fill_1 FILLER_44_1217 ();
 sg13g2_decap_8 FILLER_44_1223 ();
 sg13g2_decap_8 FILLER_44_1230 ();
 sg13g2_decap_8 FILLER_44_1237 ();
 sg13g2_decap_4 FILLER_44_1244 ();
 sg13g2_decap_8 FILLER_44_1269 ();
 sg13g2_decap_8 FILLER_44_1276 ();
 sg13g2_decap_8 FILLER_44_1283 ();
 sg13g2_decap_8 FILLER_44_1290 ();
 sg13g2_decap_4 FILLER_44_1297 ();
 sg13g2_fill_1 FILLER_44_1301 ();
 sg13g2_decap_4 FILLER_44_1312 ();
 sg13g2_fill_2 FILLER_44_1316 ();
 sg13g2_fill_2 FILLER_44_1323 ();
 sg13g2_fill_1 FILLER_44_1325 ();
 sg13g2_fill_2 FILLER_44_1347 ();
 sg13g2_fill_1 FILLER_44_1349 ();
 sg13g2_decap_8 FILLER_44_1385 ();
 sg13g2_decap_8 FILLER_44_1392 ();
 sg13g2_decap_4 FILLER_44_1399 ();
 sg13g2_fill_1 FILLER_44_1403 ();
 sg13g2_fill_2 FILLER_44_1425 ();
 sg13g2_fill_1 FILLER_44_1427 ();
 sg13g2_fill_2 FILLER_44_1454 ();
 sg13g2_decap_8 FILLER_44_1460 ();
 sg13g2_decap_8 FILLER_44_1471 ();
 sg13g2_decap_8 FILLER_44_1478 ();
 sg13g2_fill_1 FILLER_44_1485 ();
 sg13g2_fill_2 FILLER_44_1490 ();
 sg13g2_fill_1 FILLER_44_1492 ();
 sg13g2_decap_8 FILLER_44_1498 ();
 sg13g2_decap_4 FILLER_44_1505 ();
 sg13g2_fill_2 FILLER_44_1509 ();
 sg13g2_decap_8 FILLER_44_1515 ();
 sg13g2_fill_2 FILLER_44_1522 ();
 sg13g2_fill_1 FILLER_44_1528 ();
 sg13g2_decap_8 FILLER_44_1560 ();
 sg13g2_decap_8 FILLER_44_1567 ();
 sg13g2_decap_8 FILLER_44_1574 ();
 sg13g2_decap_8 FILLER_44_1581 ();
 sg13g2_decap_8 FILLER_44_1588 ();
 sg13g2_decap_8 FILLER_44_1595 ();
 sg13g2_decap_8 FILLER_44_1602 ();
 sg13g2_decap_8 FILLER_44_1609 ();
 sg13g2_decap_8 FILLER_44_1616 ();
 sg13g2_fill_2 FILLER_44_1623 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_fill_2 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_139 ();
 sg13g2_decap_8 FILLER_45_146 ();
 sg13g2_fill_2 FILLER_45_153 ();
 sg13g2_fill_1 FILLER_45_160 ();
 sg13g2_decap_8 FILLER_45_165 ();
 sg13g2_decap_8 FILLER_45_172 ();
 sg13g2_fill_2 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_181 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_4 FILLER_45_238 ();
 sg13g2_fill_1 FILLER_45_242 ();
 sg13g2_decap_8 FILLER_45_248 ();
 sg13g2_decap_8 FILLER_45_255 ();
 sg13g2_fill_2 FILLER_45_267 ();
 sg13g2_fill_1 FILLER_45_269 ();
 sg13g2_fill_2 FILLER_45_313 ();
 sg13g2_decap_8 FILLER_45_348 ();
 sg13g2_fill_1 FILLER_45_355 ();
 sg13g2_fill_2 FILLER_45_394 ();
 sg13g2_fill_1 FILLER_45_396 ();
 sg13g2_decap_4 FILLER_45_401 ();
 sg13g2_decap_8 FILLER_45_410 ();
 sg13g2_fill_2 FILLER_45_417 ();
 sg13g2_decap_4 FILLER_45_440 ();
 sg13g2_fill_2 FILLER_45_444 ();
 sg13g2_fill_2 FILLER_45_451 ();
 sg13g2_fill_1 FILLER_45_453 ();
 sg13g2_decap_8 FILLER_45_458 ();
 sg13g2_decap_4 FILLER_45_465 ();
 sg13g2_fill_1 FILLER_45_490 ();
 sg13g2_decap_4 FILLER_45_496 ();
 sg13g2_fill_1 FILLER_45_500 ();
 sg13g2_fill_1 FILLER_45_509 ();
 sg13g2_decap_8 FILLER_45_514 ();
 sg13g2_decap_8 FILLER_45_521 ();
 sg13g2_decap_8 FILLER_45_528 ();
 sg13g2_fill_1 FILLER_45_535 ();
 sg13g2_decap_8 FILLER_45_540 ();
 sg13g2_decap_4 FILLER_45_547 ();
 sg13g2_fill_2 FILLER_45_551 ();
 sg13g2_decap_8 FILLER_45_584 ();
 sg13g2_decap_8 FILLER_45_591 ();
 sg13g2_decap_4 FILLER_45_598 ();
 sg13g2_fill_2 FILLER_45_610 ();
 sg13g2_fill_2 FILLER_45_622 ();
 sg13g2_decap_4 FILLER_45_650 ();
 sg13g2_decap_8 FILLER_45_663 ();
 sg13g2_fill_1 FILLER_45_670 ();
 sg13g2_decap_4 FILLER_45_675 ();
 sg13g2_fill_2 FILLER_45_679 ();
 sg13g2_decap_4 FILLER_45_684 ();
 sg13g2_fill_2 FILLER_45_688 ();
 sg13g2_decap_8 FILLER_45_725 ();
 sg13g2_decap_8 FILLER_45_732 ();
 sg13g2_decap_4 FILLER_45_739 ();
 sg13g2_fill_1 FILLER_45_748 ();
 sg13g2_fill_1 FILLER_45_759 ();
 sg13g2_fill_2 FILLER_45_790 ();
 sg13g2_fill_1 FILLER_45_792 ();
 sg13g2_fill_2 FILLER_45_816 ();
 sg13g2_fill_1 FILLER_45_818 ();
 sg13g2_decap_8 FILLER_45_844 ();
 sg13g2_fill_2 FILLER_45_851 ();
 sg13g2_decap_8 FILLER_45_900 ();
 sg13g2_decap_8 FILLER_45_907 ();
 sg13g2_decap_8 FILLER_45_919 ();
 sg13g2_decap_8 FILLER_45_926 ();
 sg13g2_fill_1 FILLER_45_933 ();
 sg13g2_decap_8 FILLER_45_960 ();
 sg13g2_decap_8 FILLER_45_967 ();
 sg13g2_fill_2 FILLER_45_974 ();
 sg13g2_fill_1 FILLER_45_976 ();
 sg13g2_decap_8 FILLER_45_982 ();
 sg13g2_decap_4 FILLER_45_989 ();
 sg13g2_decap_8 FILLER_45_997 ();
 sg13g2_decap_4 FILLER_45_1004 ();
 sg13g2_fill_1 FILLER_45_1008 ();
 sg13g2_fill_1 FILLER_45_1030 ();
 sg13g2_decap_8 FILLER_45_1110 ();
 sg13g2_decap_4 FILLER_45_1117 ();
 sg13g2_fill_2 FILLER_45_1121 ();
 sg13g2_decap_4 FILLER_45_1152 ();
 sg13g2_fill_2 FILLER_45_1156 ();
 sg13g2_decap_4 FILLER_45_1162 ();
 sg13g2_fill_1 FILLER_45_1179 ();
 sg13g2_decap_8 FILLER_45_1209 ();
 sg13g2_decap_8 FILLER_45_1216 ();
 sg13g2_decap_4 FILLER_45_1233 ();
 sg13g2_fill_1 FILLER_45_1237 ();
 sg13g2_decap_8 FILLER_45_1242 ();
 sg13g2_decap_4 FILLER_45_1249 ();
 sg13g2_fill_1 FILLER_45_1253 ();
 sg13g2_decap_8 FILLER_45_1258 ();
 sg13g2_decap_8 FILLER_45_1301 ();
 sg13g2_decap_4 FILLER_45_1308 ();
 sg13g2_decap_8 FILLER_45_1316 ();
 sg13g2_decap_8 FILLER_45_1323 ();
 sg13g2_fill_2 FILLER_45_1330 ();
 sg13g2_decap_4 FILLER_45_1342 ();
 sg13g2_fill_2 FILLER_45_1346 ();
 sg13g2_decap_8 FILLER_45_1374 ();
 sg13g2_decap_8 FILLER_45_1381 ();
 sg13g2_fill_2 FILLER_45_1388 ();
 sg13g2_decap_8 FILLER_45_1425 ();
 sg13g2_fill_2 FILLER_45_1432 ();
 sg13g2_fill_1 FILLER_45_1434 ();
 sg13g2_decap_8 FILLER_45_1439 ();
 sg13g2_decap_8 FILLER_45_1446 ();
 sg13g2_fill_1 FILLER_45_1453 ();
 sg13g2_fill_1 FILLER_45_1510 ();
 sg13g2_decap_4 FILLER_45_1545 ();
 sg13g2_decap_8 FILLER_45_1591 ();
 sg13g2_decap_8 FILLER_45_1598 ();
 sg13g2_decap_8 FILLER_45_1605 ();
 sg13g2_decap_8 FILLER_45_1612 ();
 sg13g2_decap_4 FILLER_45_1619 ();
 sg13g2_fill_2 FILLER_45_1623 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_fill_2 FILLER_46_126 ();
 sg13g2_fill_2 FILLER_46_159 ();
 sg13g2_fill_1 FILLER_46_165 ();
 sg13g2_decap_8 FILLER_46_170 ();
 sg13g2_decap_8 FILLER_46_177 ();
 sg13g2_decap_8 FILLER_46_184 ();
 sg13g2_fill_1 FILLER_46_191 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_fill_2 FILLER_46_203 ();
 sg13g2_fill_1 FILLER_46_205 ();
 sg13g2_fill_2 FILLER_46_211 ();
 sg13g2_fill_1 FILLER_46_213 ();
 sg13g2_decap_8 FILLER_46_235 ();
 sg13g2_fill_2 FILLER_46_242 ();
 sg13g2_decap_8 FILLER_46_257 ();
 sg13g2_decap_4 FILLER_46_264 ();
 sg13g2_fill_1 FILLER_46_268 ();
 sg13g2_fill_2 FILLER_46_295 ();
 sg13g2_fill_2 FILLER_46_318 ();
 sg13g2_decap_8 FILLER_46_351 ();
 sg13g2_fill_2 FILLER_46_358 ();
 sg13g2_fill_1 FILLER_46_360 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_fill_1 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_426 ();
 sg13g2_decap_8 FILLER_46_433 ();
 sg13g2_fill_1 FILLER_46_440 ();
 sg13g2_decap_8 FILLER_46_446 ();
 sg13g2_decap_4 FILLER_46_458 ();
 sg13g2_fill_1 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_484 ();
 sg13g2_decap_8 FILLER_46_491 ();
 sg13g2_decap_8 FILLER_46_559 ();
 sg13g2_decap_8 FILLER_46_566 ();
 sg13g2_decap_8 FILLER_46_573 ();
 sg13g2_decap_8 FILLER_46_580 ();
 sg13g2_decap_4 FILLER_46_587 ();
 sg13g2_decap_4 FILLER_46_596 ();
 sg13g2_fill_1 FILLER_46_600 ();
 sg13g2_fill_1 FILLER_46_606 ();
 sg13g2_decap_8 FILLER_46_642 ();
 sg13g2_decap_8 FILLER_46_649 ();
 sg13g2_fill_2 FILLER_46_656 ();
 sg13g2_fill_2 FILLER_46_689 ();
 sg13g2_fill_2 FILLER_46_696 ();
 sg13g2_decap_8 FILLER_46_731 ();
 sg13g2_decap_8 FILLER_46_738 ();
 sg13g2_fill_2 FILLER_46_745 ();
 sg13g2_fill_2 FILLER_46_799 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_decap_8 FILLER_46_864 ();
 sg13g2_decap_8 FILLER_46_871 ();
 sg13g2_decap_4 FILLER_46_878 ();
 sg13g2_decap_8 FILLER_46_886 ();
 sg13g2_fill_1 FILLER_46_893 ();
 sg13g2_decap_8 FILLER_46_898 ();
 sg13g2_decap_8 FILLER_46_905 ();
 sg13g2_fill_2 FILLER_46_912 ();
 sg13g2_decap_4 FILLER_46_919 ();
 sg13g2_fill_1 FILLER_46_923 ();
 sg13g2_decap_8 FILLER_46_953 ();
 sg13g2_decap_8 FILLER_46_960 ();
 sg13g2_decap_4 FILLER_46_967 ();
 sg13g2_decap_8 FILLER_46_975 ();
 sg13g2_decap_8 FILLER_46_982 ();
 sg13g2_decap_8 FILLER_46_989 ();
 sg13g2_decap_8 FILLER_46_996 ();
 sg13g2_fill_2 FILLER_46_1003 ();
 sg13g2_fill_2 FILLER_46_1031 ();
 sg13g2_fill_1 FILLER_46_1033 ();
 sg13g2_fill_2 FILLER_46_1074 ();
 sg13g2_fill_1 FILLER_46_1076 ();
 sg13g2_decap_8 FILLER_46_1086 ();
 sg13g2_decap_8 FILLER_46_1093 ();
 sg13g2_decap_4 FILLER_46_1100 ();
 sg13g2_decap_8 FILLER_46_1151 ();
 sg13g2_fill_1 FILLER_46_1158 ();
 sg13g2_decap_4 FILLER_46_1190 ();
 sg13g2_fill_1 FILLER_46_1199 ();
 sg13g2_fill_1 FILLER_46_1205 ();
 sg13g2_decap_8 FILLER_46_1262 ();
 sg13g2_decap_8 FILLER_46_1269 ();
 sg13g2_fill_1 FILLER_46_1276 ();
 sg13g2_decap_4 FILLER_46_1281 ();
 sg13g2_fill_1 FILLER_46_1285 ();
 sg13g2_decap_4 FILLER_46_1290 ();
 sg13g2_decap_8 FILLER_46_1330 ();
 sg13g2_decap_8 FILLER_46_1337 ();
 sg13g2_decap_4 FILLER_46_1344 ();
 sg13g2_fill_2 FILLER_46_1348 ();
 sg13g2_decap_8 FILLER_46_1375 ();
 sg13g2_decap_8 FILLER_46_1382 ();
 sg13g2_fill_2 FILLER_46_1389 ();
 sg13g2_fill_1 FILLER_46_1391 ();
 sg13g2_decap_8 FILLER_46_1413 ();
 sg13g2_decap_8 FILLER_46_1430 ();
 sg13g2_fill_1 FILLER_46_1437 ();
 sg13g2_decap_8 FILLER_46_1451 ();
 sg13g2_decap_8 FILLER_46_1458 ();
 sg13g2_decap_8 FILLER_46_1465 ();
 sg13g2_fill_2 FILLER_46_1472 ();
 sg13g2_fill_1 FILLER_46_1474 ();
 sg13g2_decap_8 FILLER_46_1510 ();
 sg13g2_decap_8 FILLER_46_1517 ();
 sg13g2_fill_1 FILLER_46_1529 ();
 sg13g2_decap_8 FILLER_46_1555 ();
 sg13g2_decap_8 FILLER_46_1562 ();
 sg13g2_fill_1 FILLER_46_1569 ();
 sg13g2_decap_8 FILLER_46_1591 ();
 sg13g2_decap_8 FILLER_46_1598 ();
 sg13g2_decap_8 FILLER_46_1605 ();
 sg13g2_decap_8 FILLER_46_1612 ();
 sg13g2_decap_4 FILLER_46_1619 ();
 sg13g2_fill_2 FILLER_46_1623 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_4 FILLER_47_155 ();
 sg13g2_fill_1 FILLER_47_185 ();
 sg13g2_fill_2 FILLER_47_212 ();
 sg13g2_decap_8 FILLER_47_235 ();
 sg13g2_fill_2 FILLER_47_242 ();
 sg13g2_fill_1 FILLER_47_244 ();
 sg13g2_decap_8 FILLER_47_271 ();
 sg13g2_decap_8 FILLER_47_278 ();
 sg13g2_decap_8 FILLER_47_285 ();
 sg13g2_decap_8 FILLER_47_292 ();
 sg13g2_decap_8 FILLER_47_299 ();
 sg13g2_decap_8 FILLER_47_306 ();
 sg13g2_decap_8 FILLER_47_313 ();
 sg13g2_decap_8 FILLER_47_320 ();
 sg13g2_decap_8 FILLER_47_327 ();
 sg13g2_decap_8 FILLER_47_334 ();
 sg13g2_decap_8 FILLER_47_341 ();
 sg13g2_decap_8 FILLER_47_358 ();
 sg13g2_fill_1 FILLER_47_365 ();
 sg13g2_decap_4 FILLER_47_379 ();
 sg13g2_fill_1 FILLER_47_383 ();
 sg13g2_fill_2 FILLER_47_410 ();
 sg13g2_fill_1 FILLER_47_412 ();
 sg13g2_decap_4 FILLER_47_426 ();
 sg13g2_fill_2 FILLER_47_430 ();
 sg13g2_fill_1 FILLER_47_437 ();
 sg13g2_decap_4 FILLER_47_443 ();
 sg13g2_fill_1 FILLER_47_456 ();
 sg13g2_decap_8 FILLER_47_461 ();
 sg13g2_fill_2 FILLER_47_468 ();
 sg13g2_fill_2 FILLER_47_475 ();
 sg13g2_decap_8 FILLER_47_482 ();
 sg13g2_decap_8 FILLER_47_489 ();
 sg13g2_decap_8 FILLER_47_496 ();
 sg13g2_decap_4 FILLER_47_503 ();
 sg13g2_fill_1 FILLER_47_507 ();
 sg13g2_decap_8 FILLER_47_533 ();
 sg13g2_decap_8 FILLER_47_570 ();
 sg13g2_decap_8 FILLER_47_577 ();
 sg13g2_fill_1 FILLER_47_584 ();
 sg13g2_decap_4 FILLER_47_611 ();
 sg13g2_fill_1 FILLER_47_615 ();
 sg13g2_fill_1 FILLER_47_626 ();
 sg13g2_fill_2 FILLER_47_631 ();
 sg13g2_fill_1 FILLER_47_633 ();
 sg13g2_decap_8 FILLER_47_669 ();
 sg13g2_decap_4 FILLER_47_676 ();
 sg13g2_fill_1 FILLER_47_680 ();
 sg13g2_decap_4 FILLER_47_747 ();
 sg13g2_fill_2 FILLER_47_792 ();
 sg13g2_fill_2 FILLER_47_807 ();
 sg13g2_decap_8 FILLER_47_813 ();
 sg13g2_decap_8 FILLER_47_820 ();
 sg13g2_fill_2 FILLER_47_827 ();
 sg13g2_fill_1 FILLER_47_829 ();
 sg13g2_fill_2 FILLER_47_838 ();
 sg13g2_decap_8 FILLER_47_845 ();
 sg13g2_decap_4 FILLER_47_852 ();
 sg13g2_fill_1 FILLER_47_856 ();
 sg13g2_fill_1 FILLER_47_865 ();
 sg13g2_fill_2 FILLER_47_874 ();
 sg13g2_decap_4 FILLER_47_912 ();
 sg13g2_fill_2 FILLER_47_921 ();
 sg13g2_fill_1 FILLER_47_923 ();
 sg13g2_decap_4 FILLER_47_928 ();
 sg13g2_fill_2 FILLER_47_932 ();
 sg13g2_decap_8 FILLER_47_943 ();
 sg13g2_decap_8 FILLER_47_959 ();
 sg13g2_fill_2 FILLER_47_966 ();
 sg13g2_decap_4 FILLER_47_999 ();
 sg13g2_fill_1 FILLER_47_1003 ();
 sg13g2_decap_8 FILLER_47_1009 ();
 sg13g2_decap_8 FILLER_47_1016 ();
 sg13g2_decap_8 FILLER_47_1023 ();
 sg13g2_fill_2 FILLER_47_1030 ();
 sg13g2_decap_8 FILLER_47_1096 ();
 sg13g2_fill_2 FILLER_47_1103 ();
 sg13g2_fill_1 FILLER_47_1105 ();
 sg13g2_decap_8 FILLER_47_1152 ();
 sg13g2_decap_8 FILLER_47_1159 ();
 sg13g2_decap_8 FILLER_47_1166 ();
 sg13g2_decap_8 FILLER_47_1178 ();
 sg13g2_decap_8 FILLER_47_1185 ();
 sg13g2_fill_1 FILLER_47_1192 ();
 sg13g2_decap_8 FILLER_47_1197 ();
 sg13g2_decap_8 FILLER_47_1204 ();
 sg13g2_decap_4 FILLER_47_1211 ();
 sg13g2_fill_2 FILLER_47_1219 ();
 sg13g2_decap_8 FILLER_47_1246 ();
 sg13g2_decap_8 FILLER_47_1253 ();
 sg13g2_decap_4 FILLER_47_1265 ();
 sg13g2_fill_2 FILLER_47_1269 ();
 sg13g2_fill_1 FILLER_47_1276 ();
 sg13g2_decap_8 FILLER_47_1282 ();
 sg13g2_decap_8 FILLER_47_1289 ();
 sg13g2_fill_2 FILLER_47_1296 ();
 sg13g2_fill_1 FILLER_47_1298 ();
 sg13g2_fill_1 FILLER_47_1308 ();
 sg13g2_decap_4 FILLER_47_1355 ();
 sg13g2_fill_1 FILLER_47_1359 ();
 sg13g2_decap_8 FILLER_47_1364 ();
 sg13g2_fill_1 FILLER_47_1371 ();
 sg13g2_decap_8 FILLER_47_1376 ();
 sg13g2_decap_4 FILLER_47_1383 ();
 sg13g2_fill_2 FILLER_47_1387 ();
 sg13g2_decap_4 FILLER_47_1410 ();
 sg13g2_fill_2 FILLER_47_1414 ();
 sg13g2_decap_4 FILLER_47_1420 ();
 sg13g2_fill_1 FILLER_47_1424 ();
 sg13g2_decap_4 FILLER_47_1430 ();
 sg13g2_fill_1 FILLER_47_1434 ();
 sg13g2_decap_8 FILLER_47_1461 ();
 sg13g2_decap_4 FILLER_47_1468 ();
 sg13g2_decap_8 FILLER_47_1476 ();
 sg13g2_decap_8 FILLER_47_1483 ();
 sg13g2_decap_8 FILLER_47_1494 ();
 sg13g2_fill_2 FILLER_47_1501 ();
 sg13g2_fill_1 FILLER_47_1503 ();
 sg13g2_decap_4 FILLER_47_1509 ();
 sg13g2_fill_1 FILLER_47_1513 ();
 sg13g2_fill_2 FILLER_47_1543 ();
 sg13g2_fill_1 FILLER_47_1545 ();
 sg13g2_decap_8 FILLER_47_1567 ();
 sg13g2_decap_8 FILLER_47_1574 ();
 sg13g2_decap_8 FILLER_47_1581 ();
 sg13g2_decap_8 FILLER_47_1588 ();
 sg13g2_decap_8 FILLER_47_1595 ();
 sg13g2_decap_8 FILLER_47_1602 ();
 sg13g2_decap_8 FILLER_47_1609 ();
 sg13g2_decap_8 FILLER_47_1616 ();
 sg13g2_fill_2 FILLER_47_1623 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_4 FILLER_48_119 ();
 sg13g2_fill_2 FILLER_48_149 ();
 sg13g2_fill_1 FILLER_48_151 ();
 sg13g2_fill_1 FILLER_48_157 ();
 sg13g2_decap_8 FILLER_48_167 ();
 sg13g2_decap_8 FILLER_48_178 ();
 sg13g2_decap_8 FILLER_48_185 ();
 sg13g2_fill_1 FILLER_48_192 ();
 sg13g2_fill_1 FILLER_48_222 ();
 sg13g2_decap_4 FILLER_48_228 ();
 sg13g2_decap_8 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_285 ();
 sg13g2_fill_1 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_293 ();
 sg13g2_decap_4 FILLER_48_300 ();
 sg13g2_fill_2 FILLER_48_304 ();
 sg13g2_fill_1 FILLER_48_310 ();
 sg13g2_decap_4 FILLER_48_316 ();
 sg13g2_fill_1 FILLER_48_320 ();
 sg13g2_decap_8 FILLER_48_330 ();
 sg13g2_decap_8 FILLER_48_337 ();
 sg13g2_decap_8 FILLER_48_344 ();
 sg13g2_decap_4 FILLER_48_351 ();
 sg13g2_fill_2 FILLER_48_386 ();
 sg13g2_fill_1 FILLER_48_388 ();
 sg13g2_fill_2 FILLER_48_398 ();
 sg13g2_fill_1 FILLER_48_400 ();
 sg13g2_decap_4 FILLER_48_440 ();
 sg13g2_decap_8 FILLER_48_475 ();
 sg13g2_fill_2 FILLER_48_482 ();
 sg13g2_decap_8 FILLER_48_488 ();
 sg13g2_decap_8 FILLER_48_495 ();
 sg13g2_decap_4 FILLER_48_502 ();
 sg13g2_fill_1 FILLER_48_506 ();
 sg13g2_decap_8 FILLER_48_528 ();
 sg13g2_decap_8 FILLER_48_535 ();
 sg13g2_decap_4 FILLER_48_542 ();
 sg13g2_fill_2 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_fill_2 FILLER_48_588 ();
 sg13g2_fill_1 FILLER_48_590 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_609 ();
 sg13g2_fill_1 FILLER_48_616 ();
 sg13g2_decap_4 FILLER_48_622 ();
 sg13g2_fill_2 FILLER_48_626 ();
 sg13g2_decap_8 FILLER_48_632 ();
 sg13g2_decap_8 FILLER_48_639 ();
 sg13g2_decap_4 FILLER_48_646 ();
 sg13g2_decap_8 FILLER_48_654 ();
 sg13g2_decap_4 FILLER_48_661 ();
 sg13g2_fill_2 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_fill_2 FILLER_48_679 ();
 sg13g2_fill_2 FILLER_48_686 ();
 sg13g2_fill_1 FILLER_48_688 ();
 sg13g2_fill_2 FILLER_48_728 ();
 sg13g2_fill_1 FILLER_48_785 ();
 sg13g2_decap_8 FILLER_48_811 ();
 sg13g2_decap_8 FILLER_48_818 ();
 sg13g2_decap_8 FILLER_48_825 ();
 sg13g2_fill_2 FILLER_48_842 ();
 sg13g2_fill_2 FILLER_48_852 ();
 sg13g2_fill_1 FILLER_48_885 ();
 sg13g2_decap_8 FILLER_48_890 ();
 sg13g2_decap_8 FILLER_48_897 ();
 sg13g2_fill_2 FILLER_48_904 ();
 sg13g2_fill_1 FILLER_48_906 ();
 sg13g2_decap_4 FILLER_48_912 ();
 sg13g2_fill_1 FILLER_48_916 ();
 sg13g2_fill_2 FILLER_48_943 ();
 sg13g2_fill_1 FILLER_48_945 ();
 sg13g2_decap_4 FILLER_48_972 ();
 sg13g2_fill_1 FILLER_48_976 ();
 sg13g2_fill_1 FILLER_48_1007 ();
 sg13g2_decap_4 FILLER_48_1092 ();
 sg13g2_fill_1 FILLER_48_1096 ();
 sg13g2_fill_1 FILLER_48_1101 ();
 sg13g2_fill_1 FILLER_48_1123 ();
 sg13g2_fill_2 FILLER_48_1129 ();
 sg13g2_fill_1 FILLER_48_1131 ();
 sg13g2_decap_4 FILLER_48_1162 ();
 sg13g2_decap_8 FILLER_48_1170 ();
 sg13g2_decap_8 FILLER_48_1177 ();
 sg13g2_fill_1 FILLER_48_1184 ();
 sg13g2_fill_1 FILLER_48_1190 ();
 sg13g2_decap_8 FILLER_48_1195 ();
 sg13g2_fill_2 FILLER_48_1237 ();
 sg13g2_fill_1 FILLER_48_1239 ();
 sg13g2_decap_4 FILLER_48_1244 ();
 sg13g2_fill_2 FILLER_48_1248 ();
 sg13g2_fill_2 FILLER_48_1307 ();
 sg13g2_fill_1 FILLER_48_1309 ();
 sg13g2_decap_8 FILLER_48_1336 ();
 sg13g2_decap_4 FILLER_48_1343 ();
 sg13g2_fill_1 FILLER_48_1347 ();
 sg13g2_fill_1 FILLER_48_1379 ();
 sg13g2_fill_1 FILLER_48_1385 ();
 sg13g2_decap_8 FILLER_48_1394 ();
 sg13g2_decap_8 FILLER_48_1401 ();
 sg13g2_decap_8 FILLER_48_1434 ();
 sg13g2_fill_2 FILLER_48_1441 ();
 sg13g2_fill_2 FILLER_48_1456 ();
 sg13g2_fill_1 FILLER_48_1458 ();
 sg13g2_decap_4 FILLER_48_1490 ();
 sg13g2_fill_2 FILLER_48_1499 ();
 sg13g2_fill_1 FILLER_48_1501 ();
 sg13g2_decap_4 FILLER_48_1575 ();
 sg13g2_fill_2 FILLER_48_1579 ();
 sg13g2_decap_8 FILLER_48_1607 ();
 sg13g2_decap_8 FILLER_48_1614 ();
 sg13g2_decap_4 FILLER_48_1621 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_4 FILLER_49_112 ();
 sg13g2_fill_1 FILLER_49_116 ();
 sg13g2_decap_4 FILLER_49_121 ();
 sg13g2_fill_1 FILLER_49_125 ();
 sg13g2_fill_1 FILLER_49_197 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_decap_8 FILLER_49_239 ();
 sg13g2_fill_1 FILLER_49_246 ();
 sg13g2_fill_1 FILLER_49_324 ();
 sg13g2_decap_4 FILLER_49_351 ();
 sg13g2_fill_2 FILLER_49_355 ();
 sg13g2_fill_2 FILLER_49_412 ();
 sg13g2_decap_8 FILLER_49_435 ();
 sg13g2_decap_4 FILLER_49_442 ();
 sg13g2_fill_2 FILLER_49_446 ();
 sg13g2_decap_8 FILLER_49_504 ();
 sg13g2_decap_8 FILLER_49_511 ();
 sg13g2_fill_2 FILLER_49_518 ();
 sg13g2_fill_2 FILLER_49_564 ();
 sg13g2_fill_1 FILLER_49_566 ();
 sg13g2_decap_4 FILLER_49_606 ();
 sg13g2_decap_8 FILLER_49_641 ();
 sg13g2_decap_8 FILLER_49_648 ();
 sg13g2_fill_2 FILLER_49_655 ();
 sg13g2_decap_8 FILLER_49_662 ();
 sg13g2_decap_8 FILLER_49_669 ();
 sg13g2_fill_2 FILLER_49_676 ();
 sg13g2_decap_4 FILLER_49_733 ();
 sg13g2_fill_1 FILLER_49_737 ();
 sg13g2_fill_2 FILLER_49_815 ();
 sg13g2_fill_1 FILLER_49_823 ();
 sg13g2_fill_1 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_894 ();
 sg13g2_decap_8 FILLER_49_901 ();
 sg13g2_decap_8 FILLER_49_908 ();
 sg13g2_fill_2 FILLER_49_915 ();
 sg13g2_fill_1 FILLER_49_917 ();
 sg13g2_fill_2 FILLER_49_922 ();
 sg13g2_fill_2 FILLER_49_928 ();
 sg13g2_decap_8 FILLER_49_964 ();
 sg13g2_decap_4 FILLER_49_979 ();
 sg13g2_decap_4 FILLER_49_1004 ();
 sg13g2_fill_1 FILLER_49_1008 ();
 sg13g2_fill_2 FILLER_49_1030 ();
 sg13g2_fill_1 FILLER_49_1032 ();
 sg13g2_decap_8 FILLER_49_1037 ();
 sg13g2_decap_8 FILLER_49_1044 ();
 sg13g2_decap_8 FILLER_49_1051 ();
 sg13g2_fill_2 FILLER_49_1058 ();
 sg13g2_decap_8 FILLER_49_1121 ();
 sg13g2_decap_8 FILLER_49_1128 ();
 sg13g2_fill_2 FILLER_49_1135 ();
 sg13g2_fill_1 FILLER_49_1137 ();
 sg13g2_fill_1 FILLER_49_1185 ();
 sg13g2_decap_8 FILLER_49_1212 ();
 sg13g2_fill_2 FILLER_49_1223 ();
 sg13g2_decap_8 FILLER_49_1272 ();
 sg13g2_fill_2 FILLER_49_1279 ();
 sg13g2_decap_8 FILLER_49_1306 ();
 sg13g2_decap_8 FILLER_49_1313 ();
 sg13g2_decap_8 FILLER_49_1320 ();
 sg13g2_decap_8 FILLER_49_1327 ();
 sg13g2_decap_8 FILLER_49_1334 ();
 sg13g2_decap_8 FILLER_49_1341 ();
 sg13g2_fill_1 FILLER_49_1348 ();
 sg13g2_fill_2 FILLER_49_1405 ();
 sg13g2_decap_8 FILLER_49_1419 ();
 sg13g2_decap_8 FILLER_49_1431 ();
 sg13g2_decap_8 FILLER_49_1438 ();
 sg13g2_fill_2 FILLER_49_1450 ();
 sg13g2_fill_2 FILLER_49_1482 ();
 sg13g2_fill_1 FILLER_49_1484 ();
 sg13g2_fill_1 FILLER_49_1522 ();
 sg13g2_decap_8 FILLER_49_1527 ();
 sg13g2_fill_2 FILLER_49_1534 ();
 sg13g2_decap_8 FILLER_49_1540 ();
 sg13g2_fill_1 FILLER_49_1547 ();
 sg13g2_decap_8 FILLER_49_1569 ();
 sg13g2_decap_8 FILLER_49_1576 ();
 sg13g2_decap_4 FILLER_49_1583 ();
 sg13g2_decap_8 FILLER_49_1591 ();
 sg13g2_decap_8 FILLER_49_1598 ();
 sg13g2_decap_8 FILLER_49_1605 ();
 sg13g2_decap_8 FILLER_49_1612 ();
 sg13g2_decap_4 FILLER_49_1619 ();
 sg13g2_fill_2 FILLER_49_1623 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_4 FILLER_50_105 ();
 sg13g2_fill_2 FILLER_50_109 ();
 sg13g2_decap_4 FILLER_50_172 ();
 sg13g2_fill_1 FILLER_50_200 ();
 sg13g2_decap_4 FILLER_50_205 ();
 sg13g2_decap_8 FILLER_50_213 ();
 sg13g2_fill_2 FILLER_50_220 ();
 sg13g2_fill_1 FILLER_50_222 ();
 sg13g2_fill_2 FILLER_50_249 ();
 sg13g2_fill_1 FILLER_50_251 ();
 sg13g2_decap_4 FILLER_50_282 ();
 sg13g2_decap_8 FILLER_50_319 ();
 sg13g2_decap_8 FILLER_50_326 ();
 sg13g2_fill_1 FILLER_50_333 ();
 sg13g2_decap_8 FILLER_50_338 ();
 sg13g2_fill_2 FILLER_50_345 ();
 sg13g2_fill_1 FILLER_50_347 ();
 sg13g2_decap_4 FILLER_50_361 ();
 sg13g2_fill_1 FILLER_50_365 ();
 sg13g2_decap_4 FILLER_50_401 ();
 sg13g2_decap_8 FILLER_50_430 ();
 sg13g2_decap_4 FILLER_50_437 ();
 sg13g2_fill_2 FILLER_50_471 ();
 sg13g2_fill_1 FILLER_50_473 ();
 sg13g2_decap_8 FILLER_50_478 ();
 sg13g2_decap_4 FILLER_50_485 ();
 sg13g2_fill_1 FILLER_50_489 ();
 sg13g2_decap_8 FILLER_50_511 ();
 sg13g2_decap_8 FILLER_50_518 ();
 sg13g2_decap_8 FILLER_50_525 ();
 sg13g2_decap_4 FILLER_50_532 ();
 sg13g2_fill_1 FILLER_50_536 ();
 sg13g2_decap_8 FILLER_50_541 ();
 sg13g2_decap_8 FILLER_50_548 ();
 sg13g2_fill_2 FILLER_50_576 ();
 sg13g2_decap_8 FILLER_50_612 ();
 sg13g2_fill_2 FILLER_50_619 ();
 sg13g2_fill_1 FILLER_50_621 ();
 sg13g2_decap_8 FILLER_50_630 ();
 sg13g2_decap_4 FILLER_50_637 ();
 sg13g2_decap_8 FILLER_50_728 ();
 sg13g2_fill_2 FILLER_50_735 ();
 sg13g2_fill_1 FILLER_50_737 ();
 sg13g2_fill_2 FILLER_50_763 ();
 sg13g2_fill_1 FILLER_50_765 ();
 sg13g2_decap_8 FILLER_50_796 ();
 sg13g2_decap_8 FILLER_50_803 ();
 sg13g2_decap_8 FILLER_50_810 ();
 sg13g2_fill_2 FILLER_50_817 ();
 sg13g2_fill_1 FILLER_50_819 ();
 sg13g2_decap_4 FILLER_50_826 ();
 sg13g2_decap_4 FILLER_50_886 ();
 sg13g2_fill_2 FILLER_50_890 ();
 sg13g2_fill_2 FILLER_50_918 ();
 sg13g2_fill_1 FILLER_50_959 ();
 sg13g2_decap_8 FILLER_50_998 ();
 sg13g2_decap_8 FILLER_50_1005 ();
 sg13g2_decap_8 FILLER_50_1064 ();
 sg13g2_decap_4 FILLER_50_1071 ();
 sg13g2_decap_8 FILLER_50_1113 ();
 sg13g2_fill_2 FILLER_50_1120 ();
 sg13g2_fill_1 FILLER_50_1122 ();
 sg13g2_decap_8 FILLER_50_1144 ();
 sg13g2_decap_4 FILLER_50_1151 ();
 sg13g2_fill_2 FILLER_50_1155 ();
 sg13g2_decap_8 FILLER_50_1161 ();
 sg13g2_decap_8 FILLER_50_1168 ();
 sg13g2_decap_8 FILLER_50_1184 ();
 sg13g2_decap_8 FILLER_50_1191 ();
 sg13g2_decap_8 FILLER_50_1198 ();
 sg13g2_decap_8 FILLER_50_1205 ();
 sg13g2_decap_8 FILLER_50_1212 ();
 sg13g2_decap_8 FILLER_50_1219 ();
 sg13g2_decap_8 FILLER_50_1226 ();
 sg13g2_decap_8 FILLER_50_1233 ();
 sg13g2_decap_8 FILLER_50_1240 ();
 sg13g2_decap_4 FILLER_50_1247 ();
 sg13g2_fill_1 FILLER_50_1251 ();
 sg13g2_decap_8 FILLER_50_1281 ();
 sg13g2_decap_8 FILLER_50_1288 ();
 sg13g2_decap_8 FILLER_50_1295 ();
 sg13g2_decap_8 FILLER_50_1306 ();
 sg13g2_decap_8 FILLER_50_1313 ();
 sg13g2_decap_4 FILLER_50_1320 ();
 sg13g2_fill_1 FILLER_50_1324 ();
 sg13g2_decap_8 FILLER_50_1338 ();
 sg13g2_decap_8 FILLER_50_1345 ();
 sg13g2_decap_8 FILLER_50_1352 ();
 sg13g2_fill_2 FILLER_50_1385 ();
 sg13g2_fill_1 FILLER_50_1387 ();
 sg13g2_decap_4 FILLER_50_1392 ();
 sg13g2_fill_2 FILLER_50_1396 ();
 sg13g2_fill_1 FILLER_50_1407 ();
 sg13g2_fill_2 FILLER_50_1468 ();
 sg13g2_fill_2 FILLER_50_1496 ();
 sg13g2_fill_1 FILLER_50_1498 ();
 sg13g2_fill_2 FILLER_50_1525 ();
 sg13g2_decap_8 FILLER_50_1556 ();
 sg13g2_decap_4 FILLER_50_1563 ();
 sg13g2_fill_2 FILLER_50_1567 ();
 sg13g2_decap_8 FILLER_50_1590 ();
 sg13g2_decap_8 FILLER_50_1597 ();
 sg13g2_decap_8 FILLER_50_1604 ();
 sg13g2_decap_8 FILLER_50_1611 ();
 sg13g2_decap_8 FILLER_50_1618 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_4 FILLER_51_119 ();
 sg13g2_fill_2 FILLER_51_127 ();
 sg13g2_decap_8 FILLER_51_158 ();
 sg13g2_decap_8 FILLER_51_165 ();
 sg13g2_fill_1 FILLER_51_172 ();
 sg13g2_fill_2 FILLER_51_228 ();
 sg13g2_decap_4 FILLER_51_234 ();
 sg13g2_decap_8 FILLER_51_272 ();
 sg13g2_decap_8 FILLER_51_279 ();
 sg13g2_decap_4 FILLER_51_286 ();
 sg13g2_fill_2 FILLER_51_290 ();
 sg13g2_fill_2 FILLER_51_296 ();
 sg13g2_fill_1 FILLER_51_298 ();
 sg13g2_decap_8 FILLER_51_308 ();
 sg13g2_decap_8 FILLER_51_315 ();
 sg13g2_decap_8 FILLER_51_327 ();
 sg13g2_decap_8 FILLER_51_334 ();
 sg13g2_decap_8 FILLER_51_341 ();
 sg13g2_fill_2 FILLER_51_348 ();
 sg13g2_fill_1 FILLER_51_376 ();
 sg13g2_decap_8 FILLER_51_381 ();
 sg13g2_fill_2 FILLER_51_388 ();
 sg13g2_fill_1 FILLER_51_390 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_fill_2 FILLER_51_403 ();
 sg13g2_decap_8 FILLER_51_409 ();
 sg13g2_fill_1 FILLER_51_416 ();
 sg13g2_decap_4 FILLER_51_485 ();
 sg13g2_fill_2 FILLER_51_489 ();
 sg13g2_fill_2 FILLER_51_517 ();
 sg13g2_decap_8 FILLER_51_532 ();
 sg13g2_decap_8 FILLER_51_539 ();
 sg13g2_decap_8 FILLER_51_546 ();
 sg13g2_decap_4 FILLER_51_553 ();
 sg13g2_decap_8 FILLER_51_578 ();
 sg13g2_decap_4 FILLER_51_585 ();
 sg13g2_fill_1 FILLER_51_589 ();
 sg13g2_fill_2 FILLER_51_616 ();
 sg13g2_decap_8 FILLER_51_644 ();
 sg13g2_decap_4 FILLER_51_659 ();
 sg13g2_fill_2 FILLER_51_663 ();
 sg13g2_decap_4 FILLER_51_674 ();
 sg13g2_decap_4 FILLER_51_682 ();
 sg13g2_fill_1 FILLER_51_686 ();
 sg13g2_fill_1 FILLER_51_696 ();
 sg13g2_fill_1 FILLER_51_777 ();
 sg13g2_decap_8 FILLER_51_783 ();
 sg13g2_decap_8 FILLER_51_790 ();
 sg13g2_fill_2 FILLER_51_797 ();
 sg13g2_decap_8 FILLER_51_803 ();
 sg13g2_decap_8 FILLER_51_810 ();
 sg13g2_decap_4 FILLER_51_817 ();
 sg13g2_fill_2 FILLER_51_838 ();
 sg13g2_fill_1 FILLER_51_856 ();
 sg13g2_fill_2 FILLER_51_882 ();
 sg13g2_fill_2 FILLER_51_889 ();
 sg13g2_decap_8 FILLER_51_990 ();
 sg13g2_decap_8 FILLER_51_997 ();
 sg13g2_decap_8 FILLER_51_1004 ();
 sg13g2_decap_4 FILLER_51_1011 ();
 sg13g2_decap_4 FILLER_51_1036 ();
 sg13g2_decap_8 FILLER_51_1049 ();
 sg13g2_fill_2 FILLER_51_1056 ();
 sg13g2_fill_1 FILLER_51_1058 ();
 sg13g2_decap_4 FILLER_51_1063 ();
 sg13g2_fill_2 FILLER_51_1067 ();
 sg13g2_fill_2 FILLER_51_1074 ();
 sg13g2_decap_8 FILLER_51_1123 ();
 sg13g2_decap_4 FILLER_51_1130 ();
 sg13g2_fill_2 FILLER_51_1148 ();
 sg13g2_fill_1 FILLER_51_1150 ();
 sg13g2_decap_8 FILLER_51_1155 ();
 sg13g2_decap_8 FILLER_51_1162 ();
 sg13g2_fill_1 FILLER_51_1169 ();
 sg13g2_fill_1 FILLER_51_1195 ();
 sg13g2_decap_4 FILLER_51_1201 ();
 sg13g2_fill_2 FILLER_51_1209 ();
 sg13g2_fill_1 FILLER_51_1211 ();
 sg13g2_fill_2 FILLER_51_1216 ();
 sg13g2_decap_4 FILLER_51_1239 ();
 sg13g2_decap_8 FILLER_51_1248 ();
 sg13g2_decap_8 FILLER_51_1255 ();
 sg13g2_fill_2 FILLER_51_1262 ();
 sg13g2_fill_1 FILLER_51_1264 ();
 sg13g2_fill_2 FILLER_51_1352 ();
 sg13g2_decap_4 FILLER_51_1359 ();
 sg13g2_fill_2 FILLER_51_1363 ();
 sg13g2_fill_1 FILLER_51_1369 ();
 sg13g2_fill_2 FILLER_51_1404 ();
 sg13g2_fill_1 FILLER_51_1406 ();
 sg13g2_decap_8 FILLER_51_1433 ();
 sg13g2_decap_8 FILLER_51_1440 ();
 sg13g2_fill_2 FILLER_51_1447 ();
 sg13g2_decap_8 FILLER_51_1453 ();
 sg13g2_decap_8 FILLER_51_1460 ();
 sg13g2_fill_2 FILLER_51_1467 ();
 sg13g2_decap_4 FILLER_51_1473 ();
 sg13g2_fill_1 FILLER_51_1477 ();
 sg13g2_decap_8 FILLER_51_1482 ();
 sg13g2_decap_8 FILLER_51_1489 ();
 sg13g2_decap_8 FILLER_51_1496 ();
 sg13g2_decap_8 FILLER_51_1503 ();
 sg13g2_decap_4 FILLER_51_1510 ();
 sg13g2_fill_2 FILLER_51_1514 ();
 sg13g2_decap_8 FILLER_51_1551 ();
 sg13g2_decap_8 FILLER_51_1558 ();
 sg13g2_decap_8 FILLER_51_1565 ();
 sg13g2_decap_8 FILLER_51_1572 ();
 sg13g2_decap_8 FILLER_51_1579 ();
 sg13g2_decap_8 FILLER_51_1586 ();
 sg13g2_decap_8 FILLER_51_1593 ();
 sg13g2_decap_8 FILLER_51_1600 ();
 sg13g2_decap_8 FILLER_51_1607 ();
 sg13g2_decap_8 FILLER_51_1614 ();
 sg13g2_decap_4 FILLER_51_1621 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_4 FILLER_52_112 ();
 sg13g2_fill_2 FILLER_52_142 ();
 sg13g2_decap_8 FILLER_52_152 ();
 sg13g2_fill_1 FILLER_52_192 ();
 sg13g2_decap_8 FILLER_52_219 ();
 sg13g2_fill_2 FILLER_52_226 ();
 sg13g2_decap_4 FILLER_52_232 ();
 sg13g2_decap_8 FILLER_52_265 ();
 sg13g2_decap_8 FILLER_52_272 ();
 sg13g2_decap_4 FILLER_52_279 ();
 sg13g2_fill_1 FILLER_52_283 ();
 sg13g2_fill_2 FILLER_52_310 ();
 sg13g2_fill_1 FILLER_52_312 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_fill_2 FILLER_52_350 ();
 sg13g2_fill_1 FILLER_52_352 ();
 sg13g2_fill_1 FILLER_52_358 ();
 sg13g2_decap_8 FILLER_52_364 ();
 sg13g2_decap_8 FILLER_52_371 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_decap_4 FILLER_52_385 ();
 sg13g2_fill_1 FILLER_52_389 ();
 sg13g2_decap_4 FILLER_52_416 ();
 sg13g2_decap_8 FILLER_52_434 ();
 sg13g2_decap_4 FILLER_52_441 ();
 sg13g2_decap_4 FILLER_52_449 ();
 sg13g2_fill_1 FILLER_52_453 ();
 sg13g2_decap_4 FILLER_52_458 ();
 sg13g2_fill_2 FILLER_52_462 ();
 sg13g2_decap_8 FILLER_52_473 ();
 sg13g2_decap_8 FILLER_52_480 ();
 sg13g2_decap_8 FILLER_52_487 ();
 sg13g2_decap_8 FILLER_52_494 ();
 sg13g2_decap_8 FILLER_52_501 ();
 sg13g2_decap_4 FILLER_52_508 ();
 sg13g2_fill_1 FILLER_52_512 ();
 sg13g2_fill_2 FILLER_52_539 ();
 sg13g2_decap_8 FILLER_52_545 ();
 sg13g2_decap_8 FILLER_52_552 ();
 sg13g2_decap_8 FILLER_52_559 ();
 sg13g2_fill_2 FILLER_52_566 ();
 sg13g2_fill_1 FILLER_52_568 ();
 sg13g2_decap_8 FILLER_52_574 ();
 sg13g2_decap_8 FILLER_52_581 ();
 sg13g2_decap_8 FILLER_52_588 ();
 sg13g2_fill_1 FILLER_52_595 ();
 sg13g2_fill_1 FILLER_52_610 ();
 sg13g2_decap_4 FILLER_52_620 ();
 sg13g2_fill_2 FILLER_52_624 ();
 sg13g2_decap_8 FILLER_52_665 ();
 sg13g2_decap_8 FILLER_52_672 ();
 sg13g2_decap_8 FILLER_52_679 ();
 sg13g2_fill_2 FILLER_52_686 ();
 sg13g2_decap_8 FILLER_52_714 ();
 sg13g2_fill_1 FILLER_52_721 ();
 sg13g2_decap_8 FILLER_52_726 ();
 sg13g2_decap_8 FILLER_52_754 ();
 sg13g2_decap_8 FILLER_52_761 ();
 sg13g2_fill_1 FILLER_52_768 ();
 sg13g2_decap_4 FILLER_52_774 ();
 sg13g2_fill_1 FILLER_52_778 ();
 sg13g2_fill_2 FILLER_52_788 ();
 sg13g2_decap_8 FILLER_52_816 ();
 sg13g2_decap_4 FILLER_52_823 ();
 sg13g2_decap_8 FILLER_52_839 ();
 sg13g2_fill_1 FILLER_52_846 ();
 sg13g2_fill_2 FILLER_52_861 ();
 sg13g2_fill_2 FILLER_52_902 ();
 sg13g2_fill_1 FILLER_52_904 ();
 sg13g2_decap_4 FILLER_52_955 ();
 sg13g2_decap_8 FILLER_52_963 ();
 sg13g2_decap_8 FILLER_52_970 ();
 sg13g2_decap_4 FILLER_52_977 ();
 sg13g2_fill_1 FILLER_52_985 ();
 sg13g2_decap_4 FILLER_52_991 ();
 sg13g2_decap_8 FILLER_52_999 ();
 sg13g2_decap_8 FILLER_52_1006 ();
 sg13g2_decap_8 FILLER_52_1013 ();
 sg13g2_decap_8 FILLER_52_1020 ();
 sg13g2_decap_8 FILLER_52_1027 ();
 sg13g2_decap_8 FILLER_52_1038 ();
 sg13g2_decap_8 FILLER_52_1045 ();
 sg13g2_fill_1 FILLER_52_1052 ();
 sg13g2_decap_4 FILLER_52_1083 ();
 sg13g2_fill_1 FILLER_52_1087 ();
 sg13g2_decap_8 FILLER_52_1101 ();
 sg13g2_decap_8 FILLER_52_1113 ();
 sg13g2_fill_2 FILLER_52_1141 ();
 sg13g2_fill_2 FILLER_52_1169 ();
 sg13g2_decap_8 FILLER_52_1244 ();
 sg13g2_decap_8 FILLER_52_1251 ();
 sg13g2_decap_8 FILLER_52_1258 ();
 sg13g2_decap_4 FILLER_52_1265 ();
 sg13g2_fill_2 FILLER_52_1269 ();
 sg13g2_fill_2 FILLER_52_1276 ();
 sg13g2_fill_2 FILLER_52_1310 ();
 sg13g2_decap_8 FILLER_52_1317 ();
 sg13g2_decap_8 FILLER_52_1324 ();
 sg13g2_decap_8 FILLER_52_1331 ();
 sg13g2_fill_2 FILLER_52_1338 ();
 sg13g2_fill_1 FILLER_52_1340 ();
 sg13g2_fill_2 FILLER_52_1372 ();
 sg13g2_decap_8 FILLER_52_1400 ();
 sg13g2_decap_8 FILLER_52_1407 ();
 sg13g2_decap_8 FILLER_52_1414 ();
 sg13g2_decap_4 FILLER_52_1421 ();
 sg13g2_fill_1 FILLER_52_1425 ();
 sg13g2_fill_2 FILLER_52_1431 ();
 sg13g2_fill_1 FILLER_52_1433 ();
 sg13g2_fill_2 FILLER_52_1442 ();
 sg13g2_fill_1 FILLER_52_1444 ();
 sg13g2_decap_8 FILLER_52_1466 ();
 sg13g2_decap_4 FILLER_52_1473 ();
 sg13g2_decap_8 FILLER_52_1486 ();
 sg13g2_decap_8 FILLER_52_1493 ();
 sg13g2_decap_4 FILLER_52_1500 ();
 sg13g2_fill_2 FILLER_52_1509 ();
 sg13g2_decap_8 FILLER_52_1515 ();
 sg13g2_decap_8 FILLER_52_1522 ();
 sg13g2_fill_1 FILLER_52_1529 ();
 sg13g2_fill_2 FILLER_52_1535 ();
 sg13g2_decap_8 FILLER_52_1563 ();
 sg13g2_decap_8 FILLER_52_1570 ();
 sg13g2_decap_8 FILLER_52_1577 ();
 sg13g2_decap_8 FILLER_52_1584 ();
 sg13g2_decap_8 FILLER_52_1591 ();
 sg13g2_decap_8 FILLER_52_1598 ();
 sg13g2_decap_8 FILLER_52_1605 ();
 sg13g2_decap_8 FILLER_52_1612 ();
 sg13g2_decap_4 FILLER_52_1619 ();
 sg13g2_fill_2 FILLER_52_1623 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_4 FILLER_53_105 ();
 sg13g2_fill_2 FILLER_53_109 ();
 sg13g2_fill_2 FILLER_53_207 ();
 sg13g2_fill_1 FILLER_53_218 ();
 sg13g2_decap_4 FILLER_53_245 ();
 sg13g2_decap_8 FILLER_53_275 ();
 sg13g2_decap_4 FILLER_53_286 ();
 sg13g2_fill_2 FILLER_53_320 ();
 sg13g2_decap_8 FILLER_53_331 ();
 sg13g2_fill_1 FILLER_53_338 ();
 sg13g2_decap_4 FILLER_53_344 ();
 sg13g2_fill_1 FILLER_53_348 ();
 sg13g2_decap_4 FILLER_53_358 ();
 sg13g2_decap_8 FILLER_53_375 ();
 sg13g2_fill_1 FILLER_53_382 ();
 sg13g2_decap_4 FILLER_53_387 ();
 sg13g2_decap_4 FILLER_53_420 ();
 sg13g2_fill_1 FILLER_53_454 ();
 sg13g2_decap_8 FILLER_53_484 ();
 sg13g2_decap_8 FILLER_53_491 ();
 sg13g2_decap_8 FILLER_53_498 ();
 sg13g2_decap_4 FILLER_53_505 ();
 sg13g2_fill_1 FILLER_53_509 ();
 sg13g2_fill_1 FILLER_53_514 ();
 sg13g2_decap_4 FILLER_53_518 ();
 sg13g2_fill_1 FILLER_53_527 ();
 sg13g2_fill_1 FILLER_53_563 ();
 sg13g2_fill_1 FILLER_53_569 ();
 sg13g2_decap_4 FILLER_53_579 ();
 sg13g2_fill_2 FILLER_53_583 ();
 sg13g2_fill_2 FILLER_53_611 ();
 sg13g2_fill_1 FILLER_53_613 ();
 sg13g2_decap_8 FILLER_53_618 ();
 sg13g2_fill_2 FILLER_53_625 ();
 sg13g2_fill_1 FILLER_53_627 ();
 sg13g2_decap_8 FILLER_53_632 ();
 sg13g2_decap_8 FILLER_53_639 ();
 sg13g2_fill_1 FILLER_53_646 ();
 sg13g2_fill_2 FILLER_53_678 ();
 sg13g2_decap_8 FILLER_53_739 ();
 sg13g2_decap_8 FILLER_53_746 ();
 sg13g2_decap_4 FILLER_53_753 ();
 sg13g2_fill_2 FILLER_53_757 ();
 sg13g2_fill_1 FILLER_53_780 ();
 sg13g2_decap_8 FILLER_53_785 ();
 sg13g2_decap_4 FILLER_53_792 ();
 sg13g2_fill_1 FILLER_53_796 ();
 sg13g2_decap_8 FILLER_53_801 ();
 sg13g2_decap_8 FILLER_53_808 ();
 sg13g2_decap_8 FILLER_53_815 ();
 sg13g2_decap_8 FILLER_53_827 ();
 sg13g2_decap_4 FILLER_53_834 ();
 sg13g2_decap_8 FILLER_53_844 ();
 sg13g2_decap_8 FILLER_53_851 ();
 sg13g2_decap_8 FILLER_53_858 ();
 sg13g2_decap_8 FILLER_53_865 ();
 sg13g2_fill_2 FILLER_53_872 ();
 sg13g2_fill_1 FILLER_53_874 ();
 sg13g2_decap_4 FILLER_53_910 ();
 sg13g2_fill_1 FILLER_53_945 ();
 sg13g2_fill_1 FILLER_53_950 ();
 sg13g2_decap_8 FILLER_53_955 ();
 sg13g2_decap_8 FILLER_53_962 ();
 sg13g2_decap_4 FILLER_53_969 ();
 sg13g2_fill_2 FILLER_53_973 ();
 sg13g2_fill_1 FILLER_53_1001 ();
 sg13g2_fill_2 FILLER_53_1023 ();
 sg13g2_fill_1 FILLER_53_1025 ();
 sg13g2_decap_8 FILLER_53_1052 ();
 sg13g2_decap_8 FILLER_53_1059 ();
 sg13g2_decap_8 FILLER_53_1066 ();
 sg13g2_decap_8 FILLER_53_1073 ();
 sg13g2_decap_4 FILLER_53_1080 ();
 sg13g2_fill_2 FILLER_53_1084 ();
 sg13g2_decap_8 FILLER_53_1117 ();
 sg13g2_decap_8 FILLER_53_1124 ();
 sg13g2_decap_4 FILLER_53_1131 ();
 sg13g2_fill_1 FILLER_53_1135 ();
 sg13g2_decap_8 FILLER_53_1141 ();
 sg13g2_decap_8 FILLER_53_1148 ();
 sg13g2_decap_8 FILLER_53_1155 ();
 sg13g2_fill_2 FILLER_53_1162 ();
 sg13g2_fill_1 FILLER_53_1164 ();
 sg13g2_decap_8 FILLER_53_1170 ();
 sg13g2_decap_4 FILLER_53_1177 ();
 sg13g2_fill_1 FILLER_53_1181 ();
 sg13g2_decap_8 FILLER_53_1191 ();
 sg13g2_decap_8 FILLER_53_1198 ();
 sg13g2_decap_8 FILLER_53_1205 ();
 sg13g2_decap_8 FILLER_53_1212 ();
 sg13g2_decap_8 FILLER_53_1219 ();
 sg13g2_decap_8 FILLER_53_1226 ();
 sg13g2_decap_8 FILLER_53_1233 ();
 sg13g2_decap_8 FILLER_53_1240 ();
 sg13g2_decap_8 FILLER_53_1247 ();
 sg13g2_fill_2 FILLER_53_1254 ();
 sg13g2_fill_2 FILLER_53_1266 ();
 sg13g2_fill_1 FILLER_53_1268 ();
 sg13g2_decap_8 FILLER_53_1283 ();
 sg13g2_fill_1 FILLER_53_1290 ();
 sg13g2_fill_2 FILLER_53_1314 ();
 sg13g2_decap_8 FILLER_53_1330 ();
 sg13g2_decap_4 FILLER_53_1337 ();
 sg13g2_fill_1 FILLER_53_1341 ();
 sg13g2_decap_4 FILLER_53_1349 ();
 sg13g2_fill_2 FILLER_53_1357 ();
 sg13g2_decap_8 FILLER_53_1368 ();
 sg13g2_fill_1 FILLER_53_1378 ();
 sg13g2_decap_8 FILLER_53_1388 ();
 sg13g2_fill_2 FILLER_53_1395 ();
 sg13g2_fill_1 FILLER_53_1397 ();
 sg13g2_decap_8 FILLER_53_1407 ();
 sg13g2_decap_8 FILLER_53_1414 ();
 sg13g2_decap_8 FILLER_53_1421 ();
 sg13g2_fill_2 FILLER_53_1475 ();
 sg13g2_fill_1 FILLER_53_1503 ();
 sg13g2_decap_8 FILLER_53_1559 ();
 sg13g2_decap_8 FILLER_53_1566 ();
 sg13g2_decap_8 FILLER_53_1573 ();
 sg13g2_decap_8 FILLER_53_1580 ();
 sg13g2_decap_8 FILLER_53_1587 ();
 sg13g2_decap_8 FILLER_53_1594 ();
 sg13g2_decap_8 FILLER_53_1601 ();
 sg13g2_decap_8 FILLER_53_1608 ();
 sg13g2_decap_8 FILLER_53_1615 ();
 sg13g2_fill_2 FILLER_53_1622 ();
 sg13g2_fill_1 FILLER_53_1624 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_4 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_81 ();
 sg13g2_decap_8 FILLER_54_109 ();
 sg13g2_fill_1 FILLER_54_125 ();
 sg13g2_fill_2 FILLER_54_183 ();
 sg13g2_fill_1 FILLER_54_185 ();
 sg13g2_fill_2 FILLER_54_190 ();
 sg13g2_decap_8 FILLER_54_222 ();
 sg13g2_decap_8 FILLER_54_229 ();
 sg13g2_decap_4 FILLER_54_246 ();
 sg13g2_fill_2 FILLER_54_263 ();
 sg13g2_decap_8 FILLER_54_300 ();
 sg13g2_decap_8 FILLER_54_307 ();
 sg13g2_decap_8 FILLER_54_314 ();
 sg13g2_decap_8 FILLER_54_321 ();
 sg13g2_decap_8 FILLER_54_328 ();
 sg13g2_decap_8 FILLER_54_335 ();
 sg13g2_fill_1 FILLER_54_342 ();
 sg13g2_fill_1 FILLER_54_369 ();
 sg13g2_fill_2 FILLER_54_409 ();
 sg13g2_fill_1 FILLER_54_510 ();
 sg13g2_decap_8 FILLER_54_540 ();
 sg13g2_decap_8 FILLER_54_547 ();
 sg13g2_decap_8 FILLER_54_557 ();
 sg13g2_fill_2 FILLER_54_564 ();
 sg13g2_fill_1 FILLER_54_592 ();
 sg13g2_fill_1 FILLER_54_614 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_2 FILLER_54_656 ();
 sg13g2_decap_8 FILLER_54_662 ();
 sg13g2_decap_4 FILLER_54_669 ();
 sg13g2_fill_1 FILLER_54_677 ();
 sg13g2_decap_4 FILLER_54_725 ();
 sg13g2_decap_8 FILLER_54_750 ();
 sg13g2_fill_2 FILLER_54_757 ();
 sg13g2_fill_1 FILLER_54_759 ();
 sg13g2_fill_1 FILLER_54_781 ();
 sg13g2_fill_1 FILLER_54_787 ();
 sg13g2_fill_2 FILLER_54_830 ();
 sg13g2_fill_1 FILLER_54_832 ();
 sg13g2_decap_8 FILLER_54_844 ();
 sg13g2_decap_8 FILLER_54_851 ();
 sg13g2_decap_8 FILLER_54_858 ();
 sg13g2_decap_8 FILLER_54_865 ();
 sg13g2_decap_8 FILLER_54_872 ();
 sg13g2_fill_1 FILLER_54_879 ();
 sg13g2_decap_4 FILLER_54_910 ();
 sg13g2_fill_1 FILLER_54_923 ();
 sg13g2_decap_8 FILLER_54_936 ();
 sg13g2_fill_1 FILLER_54_969 ();
 sg13g2_fill_2 FILLER_54_979 ();
 sg13g2_fill_1 FILLER_54_981 ();
 sg13g2_decap_8 FILLER_54_986 ();
 sg13g2_decap_4 FILLER_54_993 ();
 sg13g2_fill_1 FILLER_54_1023 ();
 sg13g2_decap_8 FILLER_54_1034 ();
 sg13g2_decap_8 FILLER_54_1041 ();
 sg13g2_decap_8 FILLER_54_1048 ();
 sg13g2_fill_2 FILLER_54_1055 ();
 sg13g2_fill_1 FILLER_54_1090 ();
 sg13g2_fill_1 FILLER_54_1096 ();
 sg13g2_decap_8 FILLER_54_1102 ();
 sg13g2_decap_8 FILLER_54_1109 ();
 sg13g2_decap_8 FILLER_54_1116 ();
 sg13g2_decap_4 FILLER_54_1123 ();
 sg13g2_fill_2 FILLER_54_1148 ();
 sg13g2_decap_8 FILLER_54_1179 ();
 sg13g2_decap_4 FILLER_54_1186 ();
 sg13g2_decap_8 FILLER_54_1225 ();
 sg13g2_decap_8 FILLER_54_1232 ();
 sg13g2_fill_2 FILLER_54_1239 ();
 sg13g2_fill_2 FILLER_54_1262 ();
 sg13g2_fill_1 FILLER_54_1342 ();
 sg13g2_fill_2 FILLER_54_1368 ();
 sg13g2_fill_2 FILLER_54_1400 ();
 sg13g2_fill_1 FILLER_54_1402 ();
 sg13g2_decap_8 FILLER_54_1429 ();
 sg13g2_decap_8 FILLER_54_1436 ();
 sg13g2_decap_8 FILLER_54_1473 ();
 sg13g2_decap_4 FILLER_54_1480 ();
 sg13g2_fill_1 FILLER_54_1484 ();
 sg13g2_decap_4 FILLER_54_1489 ();
 sg13g2_fill_2 FILLER_54_1493 ();
 sg13g2_fill_1 FILLER_54_1500 ();
 sg13g2_fill_2 FILLER_54_1505 ();
 sg13g2_decap_8 FILLER_54_1511 ();
 sg13g2_decap_8 FILLER_54_1518 ();
 sg13g2_decap_4 FILLER_54_1525 ();
 sg13g2_fill_2 FILLER_54_1544 ();
 sg13g2_decap_8 FILLER_54_1550 ();
 sg13g2_decap_8 FILLER_54_1557 ();
 sg13g2_decap_8 FILLER_54_1564 ();
 sg13g2_decap_8 FILLER_54_1575 ();
 sg13g2_decap_8 FILLER_54_1582 ();
 sg13g2_decap_8 FILLER_54_1589 ();
 sg13g2_decap_8 FILLER_54_1596 ();
 sg13g2_decap_8 FILLER_54_1603 ();
 sg13g2_decap_8 FILLER_54_1610 ();
 sg13g2_decap_8 FILLER_54_1617 ();
 sg13g2_fill_1 FILLER_54_1624 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_4 FILLER_55_84 ();
 sg13g2_fill_2 FILLER_55_88 ();
 sg13g2_decap_8 FILLER_55_94 ();
 sg13g2_decap_4 FILLER_55_127 ();
 sg13g2_fill_2 FILLER_55_131 ();
 sg13g2_fill_1 FILLER_55_138 ();
 sg13g2_fill_2 FILLER_55_148 ();
 sg13g2_fill_1 FILLER_55_150 ();
 sg13g2_decap_8 FILLER_55_172 ();
 sg13g2_fill_2 FILLER_55_179 ();
 sg13g2_fill_1 FILLER_55_181 ();
 sg13g2_fill_1 FILLER_55_186 ();
 sg13g2_decap_8 FILLER_55_212 ();
 sg13g2_fill_2 FILLER_55_219 ();
 sg13g2_fill_1 FILLER_55_221 ();
 sg13g2_fill_2 FILLER_55_243 ();
 sg13g2_fill_1 FILLER_55_245 ();
 sg13g2_decap_8 FILLER_55_279 ();
 sg13g2_decap_8 FILLER_55_286 ();
 sg13g2_decap_4 FILLER_55_293 ();
 sg13g2_fill_1 FILLER_55_297 ();
 sg13g2_fill_2 FILLER_55_329 ();
 sg13g2_fill_1 FILLER_55_340 ();
 sg13g2_fill_1 FILLER_55_349 ();
 sg13g2_fill_2 FILLER_55_384 ();
 sg13g2_fill_1 FILLER_55_386 ();
 sg13g2_fill_2 FILLER_55_412 ();
 sg13g2_fill_2 FILLER_55_424 ();
 sg13g2_fill_1 FILLER_55_426 ();
 sg13g2_fill_1 FILLER_55_436 ();
 sg13g2_decap_4 FILLER_55_441 ();
 sg13g2_fill_1 FILLER_55_445 ();
 sg13g2_decap_8 FILLER_55_450 ();
 sg13g2_fill_2 FILLER_55_457 ();
 sg13g2_fill_1 FILLER_55_459 ();
 sg13g2_decap_8 FILLER_55_465 ();
 sg13g2_decap_8 FILLER_55_472 ();
 sg13g2_decap_4 FILLER_55_483 ();
 sg13g2_decap_8 FILLER_55_539 ();
 sg13g2_decap_4 FILLER_55_550 ();
 sg13g2_decap_8 FILLER_55_583 ();
 sg13g2_decap_8 FILLER_55_590 ();
 sg13g2_decap_8 FILLER_55_597 ();
 sg13g2_decap_8 FILLER_55_604 ();
 sg13g2_decap_8 FILLER_55_611 ();
 sg13g2_decap_8 FILLER_55_618 ();
 sg13g2_decap_8 FILLER_55_625 ();
 sg13g2_decap_8 FILLER_55_632 ();
 sg13g2_fill_2 FILLER_55_639 ();
 sg13g2_fill_1 FILLER_55_641 ();
 sg13g2_decap_8 FILLER_55_667 ();
 sg13g2_fill_1 FILLER_55_674 ();
 sg13g2_decap_8 FILLER_55_680 ();
 sg13g2_decap_8 FILLER_55_687 ();
 sg13g2_decap_8 FILLER_55_694 ();
 sg13g2_decap_8 FILLER_55_701 ();
 sg13g2_decap_4 FILLER_55_708 ();
 sg13g2_fill_1 FILLER_55_712 ();
 sg13g2_decap_8 FILLER_55_734 ();
 sg13g2_decap_4 FILLER_55_741 ();
 sg13g2_fill_1 FILLER_55_745 ();
 sg13g2_decap_8 FILLER_55_756 ();
 sg13g2_decap_8 FILLER_55_763 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_decap_8 FILLER_55_777 ();
 sg13g2_decap_4 FILLER_55_784 ();
 sg13g2_fill_2 FILLER_55_788 ();
 sg13g2_decap_4 FILLER_55_798 ();
 sg13g2_fill_2 FILLER_55_802 ();
 sg13g2_decap_8 FILLER_55_809 ();
 sg13g2_decap_8 FILLER_55_816 ();
 sg13g2_decap_8 FILLER_55_823 ();
 sg13g2_fill_2 FILLER_55_834 ();
 sg13g2_fill_1 FILLER_55_836 ();
 sg13g2_decap_8 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_55_868 ();
 sg13g2_decap_8 FILLER_55_875 ();
 sg13g2_decap_4 FILLER_55_882 ();
 sg13g2_fill_2 FILLER_55_886 ();
 sg13g2_decap_8 FILLER_55_898 ();
 sg13g2_decap_8 FILLER_55_905 ();
 sg13g2_fill_2 FILLER_55_912 ();
 sg13g2_decap_8 FILLER_55_918 ();
 sg13g2_fill_1 FILLER_55_925 ();
 sg13g2_decap_8 FILLER_55_1013 ();
 sg13g2_fill_2 FILLER_55_1049 ();
 sg13g2_fill_1 FILLER_55_1051 ();
 sg13g2_decap_8 FILLER_55_1087 ();
 sg13g2_decap_8 FILLER_55_1094 ();
 sg13g2_fill_2 FILLER_55_1101 ();
 sg13g2_decap_4 FILLER_55_1108 ();
 sg13g2_fill_1 FILLER_55_1112 ();
 sg13g2_fill_2 FILLER_55_1117 ();
 sg13g2_fill_1 FILLER_55_1119 ();
 sg13g2_fill_2 FILLER_55_1124 ();
 sg13g2_fill_1 FILLER_55_1126 ();
 sg13g2_fill_2 FILLER_55_1148 ();
 sg13g2_fill_1 FILLER_55_1150 ();
 sg13g2_fill_1 FILLER_55_1182 ();
 sg13g2_fill_1 FILLER_55_1223 ();
 sg13g2_decap_8 FILLER_55_1245 ();
 sg13g2_decap_8 FILLER_55_1252 ();
 sg13g2_decap_4 FILLER_55_1259 ();
 sg13g2_fill_2 FILLER_55_1263 ();
 sg13g2_fill_2 FILLER_55_1270 ();
 sg13g2_decap_4 FILLER_55_1276 ();
 sg13g2_fill_1 FILLER_55_1280 ();
 sg13g2_decap_8 FILLER_55_1357 ();
 sg13g2_fill_2 FILLER_55_1364 ();
 sg13g2_decap_4 FILLER_55_1392 ();
 sg13g2_fill_1 FILLER_55_1396 ();
 sg13g2_fill_2 FILLER_55_1411 ();
 sg13g2_decap_8 FILLER_55_1421 ();
 sg13g2_decap_8 FILLER_55_1428 ();
 sg13g2_decap_8 FILLER_55_1435 ();
 sg13g2_fill_1 FILLER_55_1442 ();
 sg13g2_decap_4 FILLER_55_1478 ();
 sg13g2_fill_1 FILLER_55_1482 ();
 sg13g2_decap_8 FILLER_55_1533 ();
 sg13g2_decap_4 FILLER_55_1540 ();
 sg13g2_fill_1 FILLER_55_1544 ();
 sg13g2_decap_4 FILLER_55_1549 ();
 sg13g2_fill_2 FILLER_55_1553 ();
 sg13g2_decap_8 FILLER_55_1580 ();
 sg13g2_decap_8 FILLER_55_1587 ();
 sg13g2_decap_8 FILLER_55_1594 ();
 sg13g2_decap_8 FILLER_55_1601 ();
 sg13g2_decap_8 FILLER_55_1608 ();
 sg13g2_decap_8 FILLER_55_1615 ();
 sg13g2_fill_2 FILLER_55_1622 ();
 sg13g2_fill_1 FILLER_55_1624 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_fill_2 FILLER_56_105 ();
 sg13g2_fill_1 FILLER_56_124 ();
 sg13g2_decap_8 FILLER_56_155 ();
 sg13g2_decap_8 FILLER_56_162 ();
 sg13g2_fill_1 FILLER_56_169 ();
 sg13g2_fill_2 FILLER_56_201 ();
 sg13g2_fill_1 FILLER_56_203 ();
 sg13g2_decap_4 FILLER_56_276 ();
 sg13g2_fill_2 FILLER_56_280 ();
 sg13g2_decap_8 FILLER_56_286 ();
 sg13g2_decap_4 FILLER_56_293 ();
 sg13g2_fill_1 FILLER_56_297 ();
 sg13g2_decap_4 FILLER_56_303 ();
 sg13g2_decap_8 FILLER_56_316 ();
 sg13g2_fill_2 FILLER_56_323 ();
 sg13g2_decap_4 FILLER_56_355 ();
 sg13g2_decap_4 FILLER_56_385 ();
 sg13g2_decap_4 FILLER_56_394 ();
 sg13g2_fill_2 FILLER_56_398 ();
 sg13g2_fill_1 FILLER_56_409 ();
 sg13g2_fill_2 FILLER_56_460 ();
 sg13g2_decap_8 FILLER_56_497 ();
 sg13g2_fill_2 FILLER_56_504 ();
 sg13g2_decap_8 FILLER_56_511 ();
 sg13g2_decap_8 FILLER_56_518 ();
 sg13g2_fill_2 FILLER_56_525 ();
 sg13g2_fill_1 FILLER_56_531 ();
 sg13g2_decap_4 FILLER_56_558 ();
 sg13g2_fill_1 FILLER_56_562 ();
 sg13g2_decap_8 FILLER_56_568 ();
 sg13g2_decap_8 FILLER_56_575 ();
 sg13g2_decap_8 FILLER_56_582 ();
 sg13g2_fill_2 FILLER_56_589 ();
 sg13g2_decap_4 FILLER_56_617 ();
 sg13g2_decap_4 FILLER_56_626 ();
 sg13g2_fill_2 FILLER_56_630 ();
 sg13g2_fill_2 FILLER_56_636 ();
 sg13g2_fill_1 FILLER_56_638 ();
 sg13g2_decap_4 FILLER_56_665 ();
 sg13g2_fill_2 FILLER_56_669 ();
 sg13g2_decap_4 FILLER_56_692 ();
 sg13g2_fill_2 FILLER_56_696 ();
 sg13g2_decap_8 FILLER_56_707 ();
 sg13g2_fill_2 FILLER_56_714 ();
 sg13g2_fill_1 FILLER_56_758 ();
 sg13g2_decap_8 FILLER_56_764 ();
 sg13g2_decap_8 FILLER_56_771 ();
 sg13g2_decap_4 FILLER_56_778 ();
 sg13g2_fill_2 FILLER_56_842 ();
 sg13g2_fill_1 FILLER_56_844 ();
 sg13g2_fill_1 FILLER_56_851 ();
 sg13g2_fill_2 FILLER_56_857 ();
 sg13g2_fill_2 FILLER_56_863 ();
 sg13g2_fill_2 FILLER_56_870 ();
 sg13g2_fill_2 FILLER_56_911 ();
 sg13g2_fill_1 FILLER_56_913 ();
 sg13g2_decap_4 FILLER_56_945 ();
 sg13g2_decap_4 FILLER_56_970 ();
 sg13g2_fill_2 FILLER_56_1000 ();
 sg13g2_fill_1 FILLER_56_1028 ();
 sg13g2_decap_8 FILLER_56_1055 ();
 sg13g2_fill_1 FILLER_56_1062 ();
 sg13g2_decap_8 FILLER_56_1067 ();
 sg13g2_decap_8 FILLER_56_1074 ();
 sg13g2_fill_1 FILLER_56_1081 ();
 sg13g2_fill_1 FILLER_56_1103 ();
 sg13g2_decap_8 FILLER_56_1130 ();
 sg13g2_decap_4 FILLER_56_1137 ();
 sg13g2_fill_2 FILLER_56_1141 ();
 sg13g2_decap_8 FILLER_56_1148 ();
 sg13g2_decap_8 FILLER_56_1155 ();
 sg13g2_fill_1 FILLER_56_1162 ();
 sg13g2_decap_8 FILLER_56_1167 ();
 sg13g2_decap_4 FILLER_56_1174 ();
 sg13g2_fill_1 FILLER_56_1187 ();
 sg13g2_fill_1 FILLER_56_1193 ();
 sg13g2_fill_1 FILLER_56_1198 ();
 sg13g2_decap_8 FILLER_56_1203 ();
 sg13g2_decap_8 FILLER_56_1210 ();
 sg13g2_fill_2 FILLER_56_1217 ();
 sg13g2_decap_8 FILLER_56_1240 ();
 sg13g2_decap_4 FILLER_56_1247 ();
 sg13g2_fill_1 FILLER_56_1251 ();
 sg13g2_decap_8 FILLER_56_1261 ();
 sg13g2_decap_8 FILLER_56_1268 ();
 sg13g2_fill_1 FILLER_56_1280 ();
 sg13g2_decap_8 FILLER_56_1285 ();
 sg13g2_fill_1 FILLER_56_1292 ();
 sg13g2_decap_8 FILLER_56_1344 ();
 sg13g2_decap_8 FILLER_56_1351 ();
 sg13g2_decap_8 FILLER_56_1358 ();
 sg13g2_decap_8 FILLER_56_1365 ();
 sg13g2_fill_1 FILLER_56_1372 ();
 sg13g2_decap_4 FILLER_56_1377 ();
 sg13g2_decap_8 FILLER_56_1385 ();
 sg13g2_fill_1 FILLER_56_1392 ();
 sg13g2_fill_1 FILLER_56_1403 ();
 sg13g2_decap_4 FILLER_56_1430 ();
 sg13g2_fill_1 FILLER_56_1434 ();
 sg13g2_fill_1 FILLER_56_1440 ();
 sg13g2_fill_1 FILLER_56_1445 ();
 sg13g2_fill_1 FILLER_56_1488 ();
 sg13g2_fill_1 FILLER_56_1524 ();
 sg13g2_fill_2 FILLER_56_1529 ();
 sg13g2_fill_1 FILLER_56_1531 ();
 sg13g2_decap_8 FILLER_56_1589 ();
 sg13g2_decap_8 FILLER_56_1596 ();
 sg13g2_decap_8 FILLER_56_1603 ();
 sg13g2_decap_8 FILLER_56_1610 ();
 sg13g2_decap_8 FILLER_56_1617 ();
 sg13g2_fill_1 FILLER_56_1624 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_fill_2 FILLER_57_105 ();
 sg13g2_fill_1 FILLER_57_107 ();
 sg13g2_decap_8 FILLER_57_143 ();
 sg13g2_decap_8 FILLER_57_150 ();
 sg13g2_decap_8 FILLER_57_157 ();
 sg13g2_decap_8 FILLER_57_164 ();
 sg13g2_decap_8 FILLER_57_171 ();
 sg13g2_decap_8 FILLER_57_178 ();
 sg13g2_decap_4 FILLER_57_185 ();
 sg13g2_fill_2 FILLER_57_189 ();
 sg13g2_fill_2 FILLER_57_199 ();
 sg13g2_decap_8 FILLER_57_222 ();
 sg13g2_decap_8 FILLER_57_229 ();
 sg13g2_decap_8 FILLER_57_236 ();
 sg13g2_decap_8 FILLER_57_243 ();
 sg13g2_decap_8 FILLER_57_250 ();
 sg13g2_decap_8 FILLER_57_257 ();
 sg13g2_fill_1 FILLER_57_264 ();
 sg13g2_decap_8 FILLER_57_300 ();
 sg13g2_decap_8 FILLER_57_311 ();
 sg13g2_decap_8 FILLER_57_318 ();
 sg13g2_fill_1 FILLER_57_325 ();
 sg13g2_fill_2 FILLER_57_381 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_fill_2 FILLER_57_399 ();
 sg13g2_fill_1 FILLER_57_401 ();
 sg13g2_fill_1 FILLER_57_428 ();
 sg13g2_decap_4 FILLER_57_489 ();
 sg13g2_fill_1 FILLER_57_493 ();
 sg13g2_fill_2 FILLER_57_498 ();
 sg13g2_fill_1 FILLER_57_500 ();
 sg13g2_decap_4 FILLER_57_552 ();
 sg13g2_decap_8 FILLER_57_577 ();
 sg13g2_decap_8 FILLER_57_584 ();
 sg13g2_decap_4 FILLER_57_591 ();
 sg13g2_decap_8 FILLER_57_646 ();
 sg13g2_decap_8 FILLER_57_653 ();
 sg13g2_fill_2 FILLER_57_660 ();
 sg13g2_decap_8 FILLER_57_688 ();
 sg13g2_decap_4 FILLER_57_695 ();
 sg13g2_decap_8 FILLER_57_725 ();
 sg13g2_decap_8 FILLER_57_732 ();
 sg13g2_decap_8 FILLER_57_739 ();
 sg13g2_decap_8 FILLER_57_746 ();
 sg13g2_decap_8 FILLER_57_753 ();
 sg13g2_decap_8 FILLER_57_781 ();
 sg13g2_decap_4 FILLER_57_788 ();
 sg13g2_fill_1 FILLER_57_792 ();
 sg13g2_decap_8 FILLER_57_818 ();
 sg13g2_fill_2 FILLER_57_825 ();
 sg13g2_decap_8 FILLER_57_852 ();
 sg13g2_decap_8 FILLER_57_859 ();
 sg13g2_decap_8 FILLER_57_866 ();
 sg13g2_decap_4 FILLER_57_873 ();
 sg13g2_fill_1 FILLER_57_877 ();
 sg13g2_decap_8 FILLER_57_882 ();
 sg13g2_decap_8 FILLER_57_889 ();
 sg13g2_fill_2 FILLER_57_896 ();
 sg13g2_decap_8 FILLER_57_928 ();
 sg13g2_decap_8 FILLER_57_935 ();
 sg13g2_decap_8 FILLER_57_942 ();
 sg13g2_decap_8 FILLER_57_949 ();
 sg13g2_decap_8 FILLER_57_956 ();
 sg13g2_fill_2 FILLER_57_963 ();
 sg13g2_fill_1 FILLER_57_965 ();
 sg13g2_decap_8 FILLER_57_971 ();
 sg13g2_decap_8 FILLER_57_978 ();
 sg13g2_decap_8 FILLER_57_985 ();
 sg13g2_decap_8 FILLER_57_992 ();
 sg13g2_fill_2 FILLER_57_999 ();
 sg13g2_fill_1 FILLER_57_1001 ();
 sg13g2_decap_8 FILLER_57_1006 ();
 sg13g2_decap_8 FILLER_57_1013 ();
 sg13g2_decap_8 FILLER_57_1023 ();
 sg13g2_decap_4 FILLER_57_1030 ();
 sg13g2_fill_1 FILLER_57_1034 ();
 sg13g2_decap_8 FILLER_57_1039 ();
 sg13g2_decap_8 FILLER_57_1046 ();
 sg13g2_decap_4 FILLER_57_1053 ();
 sg13g2_decap_8 FILLER_57_1062 ();
 sg13g2_decap_4 FILLER_57_1069 ();
 sg13g2_fill_2 FILLER_57_1073 ();
 sg13g2_decap_4 FILLER_57_1079 ();
 sg13g2_fill_1 FILLER_57_1083 ();
 sg13g2_decap_4 FILLER_57_1105 ();
 sg13g2_fill_1 FILLER_57_1109 ();
 sg13g2_decap_8 FILLER_57_1144 ();
 sg13g2_decap_4 FILLER_57_1151 ();
 sg13g2_fill_2 FILLER_57_1155 ();
 sg13g2_decap_8 FILLER_57_1162 ();
 sg13g2_fill_2 FILLER_57_1169 ();
 sg13g2_decap_4 FILLER_57_1202 ();
 sg13g2_fill_1 FILLER_57_1206 ();
 sg13g2_decap_4 FILLER_57_1212 ();
 sg13g2_fill_2 FILLER_57_1216 ();
 sg13g2_decap_8 FILLER_57_1222 ();
 sg13g2_fill_2 FILLER_57_1229 ();
 sg13g2_fill_1 FILLER_57_1231 ();
 sg13g2_fill_2 FILLER_57_1237 ();
 sg13g2_decap_4 FILLER_57_1300 ();
 sg13g2_fill_1 FILLER_57_1304 ();
 sg13g2_fill_1 FILLER_57_1336 ();
 sg13g2_decap_8 FILLER_57_1342 ();
 sg13g2_decap_8 FILLER_57_1349 ();
 sg13g2_fill_2 FILLER_57_1356 ();
 sg13g2_fill_2 FILLER_57_1392 ();
 sg13g2_fill_1 FILLER_57_1394 ();
 sg13g2_decap_8 FILLER_57_1421 ();
 sg13g2_decap_8 FILLER_57_1428 ();
 sg13g2_decap_4 FILLER_57_1440 ();
 sg13g2_decap_8 FILLER_57_1453 ();
 sg13g2_decap_8 FILLER_57_1460 ();
 sg13g2_decap_8 FILLER_57_1467 ();
 sg13g2_decap_8 FILLER_57_1474 ();
 sg13g2_decap_8 FILLER_57_1481 ();
 sg13g2_decap_8 FILLER_57_1488 ();
 sg13g2_fill_1 FILLER_57_1495 ();
 sg13g2_fill_1 FILLER_57_1500 ();
 sg13g2_decap_8 FILLER_57_1536 ();
 sg13g2_decap_8 FILLER_57_1593 ();
 sg13g2_decap_4 FILLER_57_1600 ();
 sg13g2_fill_2 FILLER_57_1604 ();
 sg13g2_decap_8 FILLER_57_1610 ();
 sg13g2_decap_8 FILLER_57_1617 ();
 sg13g2_fill_1 FILLER_57_1624 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_112 ();
 sg13g2_fill_2 FILLER_58_147 ();
 sg13g2_fill_1 FILLER_58_149 ();
 sg13g2_decap_8 FILLER_58_171 ();
 sg13g2_decap_4 FILLER_58_178 ();
 sg13g2_fill_1 FILLER_58_182 ();
 sg13g2_decap_4 FILLER_58_217 ();
 sg13g2_decap_8 FILLER_58_242 ();
 sg13g2_decap_8 FILLER_58_249 ();
 sg13g2_decap_8 FILLER_58_261 ();
 sg13g2_fill_2 FILLER_58_268 ();
 sg13g2_fill_1 FILLER_58_270 ();
 sg13g2_decap_8 FILLER_58_275 ();
 sg13g2_decap_8 FILLER_58_282 ();
 sg13g2_decap_4 FILLER_58_289 ();
 sg13g2_fill_1 FILLER_58_298 ();
 sg13g2_decap_8 FILLER_58_325 ();
 sg13g2_decap_8 FILLER_58_358 ();
 sg13g2_decap_8 FILLER_58_369 ();
 sg13g2_fill_2 FILLER_58_376 ();
 sg13g2_fill_2 FILLER_58_404 ();
 sg13g2_fill_1 FILLER_58_460 ();
 sg13g2_decap_8 FILLER_58_502 ();
 sg13g2_decap_4 FILLER_58_513 ();
 sg13g2_fill_2 FILLER_58_517 ();
 sg13g2_fill_2 FILLER_58_554 ();
 sg13g2_decap_8 FILLER_58_577 ();
 sg13g2_fill_1 FILLER_58_584 ();
 sg13g2_decap_8 FILLER_58_606 ();
 sg13g2_decap_8 FILLER_58_613 ();
 sg13g2_decap_8 FILLER_58_620 ();
 sg13g2_decap_4 FILLER_58_627 ();
 sg13g2_fill_2 FILLER_58_660 ();
 sg13g2_fill_2 FILLER_58_667 ();
 sg13g2_fill_1 FILLER_58_669 ();
 sg13g2_decap_4 FILLER_58_674 ();
 sg13g2_decap_8 FILLER_58_683 ();
 sg13g2_decap_4 FILLER_58_690 ();
 sg13g2_fill_1 FILLER_58_694 ();
 sg13g2_fill_1 FILLER_58_700 ();
 sg13g2_decap_8 FILLER_58_709 ();
 sg13g2_decap_8 FILLER_58_716 ();
 sg13g2_fill_1 FILLER_58_728 ();
 sg13g2_fill_2 FILLER_58_760 ();
 sg13g2_fill_1 FILLER_58_762 ();
 sg13g2_decap_8 FILLER_58_784 ();
 sg13g2_decap_4 FILLER_58_791 ();
 sg13g2_fill_2 FILLER_58_795 ();
 sg13g2_decap_8 FILLER_58_801 ();
 sg13g2_decap_4 FILLER_58_808 ();
 sg13g2_fill_2 FILLER_58_817 ();
 sg13g2_fill_1 FILLER_58_819 ();
 sg13g2_fill_2 FILLER_58_826 ();
 sg13g2_fill_1 FILLER_58_828 ();
 sg13g2_decap_8 FILLER_58_865 ();
 sg13g2_decap_8 FILLER_58_872 ();
 sg13g2_fill_2 FILLER_58_879 ();
 sg13g2_fill_1 FILLER_58_885 ();
 sg13g2_decap_8 FILLER_58_911 ();
 sg13g2_decap_4 FILLER_58_918 ();
 sg13g2_fill_2 FILLER_58_922 ();
 sg13g2_decap_8 FILLER_58_955 ();
 sg13g2_fill_2 FILLER_58_962 ();
 sg13g2_decap_8 FILLER_58_979 ();
 sg13g2_decap_8 FILLER_58_986 ();
 sg13g2_decap_8 FILLER_58_993 ();
 sg13g2_fill_1 FILLER_58_1000 ();
 sg13g2_decap_8 FILLER_58_1014 ();
 sg13g2_decap_8 FILLER_58_1021 ();
 sg13g2_decap_8 FILLER_58_1028 ();
 sg13g2_fill_1 FILLER_58_1039 ();
 sg13g2_decap_8 FILLER_58_1045 ();
 sg13g2_decap_4 FILLER_58_1052 ();
 sg13g2_fill_2 FILLER_58_1056 ();
 sg13g2_decap_8 FILLER_58_1084 ();
 sg13g2_decap_8 FILLER_58_1091 ();
 sg13g2_decap_8 FILLER_58_1098 ();
 sg13g2_decap_4 FILLER_58_1105 ();
 sg13g2_decap_8 FILLER_58_1142 ();
 sg13g2_decap_4 FILLER_58_1200 ();
 sg13g2_decap_8 FILLER_58_1235 ();
 sg13g2_decap_8 FILLER_58_1242 ();
 sg13g2_decap_8 FILLER_58_1249 ();
 sg13g2_decap_8 FILLER_58_1256 ();
 sg13g2_decap_8 FILLER_58_1263 ();
 sg13g2_decap_8 FILLER_58_1270 ();
 sg13g2_fill_2 FILLER_58_1277 ();
 sg13g2_fill_2 FILLER_58_1288 ();
 sg13g2_decap_4 FILLER_58_1294 ();
 sg13g2_fill_2 FILLER_58_1298 ();
 sg13g2_fill_2 FILLER_58_1372 ();
 sg13g2_decap_8 FILLER_58_1425 ();
 sg13g2_fill_1 FILLER_58_1432 ();
 sg13g2_fill_1 FILLER_58_1459 ();
 sg13g2_fill_1 FILLER_58_1491 ();
 sg13g2_decap_4 FILLER_58_1521 ();
 sg13g2_fill_2 FILLER_58_1525 ();
 sg13g2_fill_1 FILLER_58_1588 ();
 sg13g2_fill_1 FILLER_58_1624 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_4 FILLER_59_112 ();
 sg13g2_decap_4 FILLER_59_146 ();
 sg13g2_decap_8 FILLER_59_171 ();
 sg13g2_decap_8 FILLER_59_178 ();
 sg13g2_fill_2 FILLER_59_185 ();
 sg13g2_fill_1 FILLER_59_187 ();
 sg13g2_decap_8 FILLER_59_214 ();
 sg13g2_decap_8 FILLER_59_221 ();
 sg13g2_fill_2 FILLER_59_228 ();
 sg13g2_decap_4 FILLER_59_251 ();
 sg13g2_fill_1 FILLER_59_255 ();
 sg13g2_decap_4 FILLER_59_282 ();
 sg13g2_fill_1 FILLER_59_286 ();
 sg13g2_decap_8 FILLER_59_321 ();
 sg13g2_fill_2 FILLER_59_332 ();
 sg13g2_fill_1 FILLER_59_334 ();
 sg13g2_decap_8 FILLER_59_344 ();
 sg13g2_decap_4 FILLER_59_351 ();
 sg13g2_decap_4 FILLER_59_376 ();
 sg13g2_fill_2 FILLER_59_419 ();
 sg13g2_fill_1 FILLER_59_421 ();
 sg13g2_decap_8 FILLER_59_516 ();
 sg13g2_decap_8 FILLER_59_523 ();
 sg13g2_decap_4 FILLER_59_530 ();
 sg13g2_fill_1 FILLER_59_534 ();
 sg13g2_fill_1 FILLER_59_544 ();
 sg13g2_decap_8 FILLER_59_549 ();
 sg13g2_fill_1 FILLER_59_556 ();
 sg13g2_decap_8 FILLER_59_561 ();
 sg13g2_decap_8 FILLER_59_568 ();
 sg13g2_decap_4 FILLER_59_575 ();
 sg13g2_fill_2 FILLER_59_579 ();
 sg13g2_decap_8 FILLER_59_607 ();
 sg13g2_fill_1 FILLER_59_614 ();
 sg13g2_fill_1 FILLER_59_650 ();
 sg13g2_decap_4 FILLER_59_677 ();
 sg13g2_decap_8 FILLER_59_721 ();
 sg13g2_decap_8 FILLER_59_728 ();
 sg13g2_decap_8 FILLER_59_735 ();
 sg13g2_fill_2 FILLER_59_776 ();
 sg13g2_fill_1 FILLER_59_778 ();
 sg13g2_decap_4 FILLER_59_814 ();
 sg13g2_fill_1 FILLER_59_830 ();
 sg13g2_fill_2 FILLER_59_837 ();
 sg13g2_fill_2 FILLER_59_861 ();
 sg13g2_fill_1 FILLER_59_863 ();
 sg13g2_fill_1 FILLER_59_873 ();
 sg13g2_fill_1 FILLER_59_909 ();
 sg13g2_decap_4 FILLER_59_914 ();
 sg13g2_fill_1 FILLER_59_918 ();
 sg13g2_fill_2 FILLER_59_924 ();
 sg13g2_fill_1 FILLER_59_926 ();
 sg13g2_fill_2 FILLER_59_952 ();
 sg13g2_decap_8 FILLER_59_996 ();
 sg13g2_fill_1 FILLER_59_1064 ();
 sg13g2_decap_8 FILLER_59_1069 ();
 sg13g2_decap_8 FILLER_59_1076 ();
 sg13g2_decap_8 FILLER_59_1083 ();
 sg13g2_decap_8 FILLER_59_1090 ();
 sg13g2_decap_8 FILLER_59_1128 ();
 sg13g2_decap_8 FILLER_59_1135 ();
 sg13g2_decap_8 FILLER_59_1142 ();
 sg13g2_decap_8 FILLER_59_1149 ();
 sg13g2_decap_8 FILLER_59_1164 ();
 sg13g2_fill_2 FILLER_59_1171 ();
 sg13g2_decap_4 FILLER_59_1211 ();
 sg13g2_fill_2 FILLER_59_1215 ();
 sg13g2_decap_8 FILLER_59_1221 ();
 sg13g2_decap_8 FILLER_59_1228 ();
 sg13g2_decap_8 FILLER_59_1235 ();
 sg13g2_decap_8 FILLER_59_1242 ();
 sg13g2_decap_8 FILLER_59_1249 ();
 sg13g2_decap_8 FILLER_59_1256 ();
 sg13g2_decap_8 FILLER_59_1263 ();
 sg13g2_decap_8 FILLER_59_1270 ();
 sg13g2_fill_1 FILLER_59_1277 ();
 sg13g2_fill_1 FILLER_59_1314 ();
 sg13g2_fill_1 FILLER_59_1345 ();
 sg13g2_fill_1 FILLER_59_1376 ();
 sg13g2_decap_4 FILLER_59_1437 ();
 sg13g2_fill_1 FILLER_59_1441 ();
 sg13g2_decap_8 FILLER_59_1446 ();
 sg13g2_fill_1 FILLER_59_1453 ();
 sg13g2_decap_8 FILLER_59_1485 ();
 sg13g2_decap_4 FILLER_59_1492 ();
 sg13g2_fill_1 FILLER_59_1522 ();
 sg13g2_decap_8 FILLER_59_1528 ();
 sg13g2_decap_4 FILLER_59_1535 ();
 sg13g2_decap_8 FILLER_59_1585 ();
 sg13g2_decap_4 FILLER_59_1592 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_fill_2 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_97 ();
 sg13g2_decap_4 FILLER_60_104 ();
 sg13g2_fill_2 FILLER_60_108 ();
 sg13g2_fill_2 FILLER_60_115 ();
 sg13g2_decap_8 FILLER_60_155 ();
 sg13g2_fill_2 FILLER_60_162 ();
 sg13g2_fill_1 FILLER_60_164 ();
 sg13g2_decap_8 FILLER_60_200 ();
 sg13g2_fill_1 FILLER_60_207 ();
 sg13g2_fill_2 FILLER_60_229 ();
 sg13g2_fill_1 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_237 ();
 sg13g2_decap_8 FILLER_60_244 ();
 sg13g2_decap_8 FILLER_60_251 ();
 sg13g2_decap_4 FILLER_60_258 ();
 sg13g2_fill_2 FILLER_60_262 ();
 sg13g2_decap_8 FILLER_60_268 ();
 sg13g2_decap_8 FILLER_60_275 ();
 sg13g2_fill_1 FILLER_60_282 ();
 sg13g2_decap_4 FILLER_60_318 ();
 sg13g2_fill_2 FILLER_60_348 ();
 sg13g2_fill_1 FILLER_60_355 ();
 sg13g2_decap_8 FILLER_60_377 ();
 sg13g2_fill_1 FILLER_60_431 ();
 sg13g2_fill_1 FILLER_60_453 ();
 sg13g2_decap_8 FILLER_60_515 ();
 sg13g2_decap_8 FILLER_60_522 ();
 sg13g2_decap_8 FILLER_60_529 ();
 sg13g2_fill_1 FILLER_60_536 ();
 sg13g2_fill_2 FILLER_60_542 ();
 sg13g2_fill_1 FILLER_60_544 ();
 sg13g2_decap_8 FILLER_60_581 ();
 sg13g2_decap_8 FILLER_60_588 ();
 sg13g2_decap_8 FILLER_60_595 ();
 sg13g2_decap_8 FILLER_60_602 ();
 sg13g2_decap_8 FILLER_60_609 ();
 sg13g2_decap_8 FILLER_60_616 ();
 sg13g2_decap_8 FILLER_60_623 ();
 sg13g2_decap_4 FILLER_60_630 ();
 sg13g2_fill_1 FILLER_60_634 ();
 sg13g2_decap_8 FILLER_60_638 ();
 sg13g2_decap_8 FILLER_60_645 ();
 sg13g2_decap_4 FILLER_60_652 ();
 sg13g2_fill_1 FILLER_60_656 ();
 sg13g2_decap_4 FILLER_60_661 ();
 sg13g2_fill_1 FILLER_60_665 ();
 sg13g2_decap_4 FILLER_60_670 ();
 sg13g2_decap_4 FILLER_60_678 ();
 sg13g2_fill_2 FILLER_60_682 ();
 sg13g2_fill_2 FILLER_60_731 ();
 sg13g2_fill_1 FILLER_60_733 ();
 sg13g2_decap_8 FILLER_60_769 ();
 sg13g2_decap_8 FILLER_60_780 ();
 sg13g2_decap_8 FILLER_60_787 ();
 sg13g2_decap_8 FILLER_60_794 ();
 sg13g2_decap_8 FILLER_60_805 ();
 sg13g2_decap_4 FILLER_60_812 ();
 sg13g2_fill_1 FILLER_60_816 ();
 sg13g2_decap_8 FILLER_60_828 ();
 sg13g2_fill_2 FILLER_60_835 ();
 sg13g2_fill_2 FILLER_60_846 ();
 sg13g2_fill_1 FILLER_60_848 ();
 sg13g2_fill_2 FILLER_60_859 ();
 sg13g2_decap_8 FILLER_60_886 ();
 sg13g2_fill_2 FILLER_60_893 ();
 sg13g2_fill_1 FILLER_60_895 ();
 sg13g2_decap_4 FILLER_60_901 ();
 sg13g2_fill_1 FILLER_60_905 ();
 sg13g2_decap_8 FILLER_60_932 ();
 sg13g2_decap_8 FILLER_60_939 ();
 sg13g2_decap_8 FILLER_60_946 ();
 sg13g2_decap_8 FILLER_60_953 ();
 sg13g2_decap_8 FILLER_60_960 ();
 sg13g2_decap_8 FILLER_60_967 ();
 sg13g2_decap_8 FILLER_60_974 ();
 sg13g2_decap_8 FILLER_60_981 ();
 sg13g2_fill_1 FILLER_60_988 ();
 sg13g2_decap_8 FILLER_60_994 ();
 sg13g2_decap_8 FILLER_60_1001 ();
 sg13g2_decap_8 FILLER_60_1008 ();
 sg13g2_fill_2 FILLER_60_1015 ();
 sg13g2_fill_1 FILLER_60_1017 ();
 sg13g2_decap_8 FILLER_60_1067 ();
 sg13g2_decap_4 FILLER_60_1074 ();
 sg13g2_fill_2 FILLER_60_1078 ();
 sg13g2_decap_4 FILLER_60_1084 ();
 sg13g2_fill_1 FILLER_60_1088 ();
 sg13g2_decap_8 FILLER_60_1124 ();
 sg13g2_fill_2 FILLER_60_1131 ();
 sg13g2_fill_1 FILLER_60_1133 ();
 sg13g2_decap_8 FILLER_60_1144 ();
 sg13g2_decap_8 FILLER_60_1151 ();
 sg13g2_decap_8 FILLER_60_1158 ();
 sg13g2_decap_8 FILLER_60_1165 ();
 sg13g2_decap_4 FILLER_60_1172 ();
 sg13g2_fill_1 FILLER_60_1176 ();
 sg13g2_decap_4 FILLER_60_1200 ();
 sg13g2_fill_2 FILLER_60_1204 ();
 sg13g2_fill_2 FILLER_60_1248 ();
 sg13g2_fill_1 FILLER_60_1250 ();
 sg13g2_fill_2 FILLER_60_1260 ();
 sg13g2_fill_1 FILLER_60_1262 ();
 sg13g2_decap_8 FILLER_60_1267 ();
 sg13g2_decap_8 FILLER_60_1274 ();
 sg13g2_decap_8 FILLER_60_1281 ();
 sg13g2_fill_1 FILLER_60_1288 ();
 sg13g2_decap_8 FILLER_60_1293 ();
 sg13g2_fill_1 FILLER_60_1300 ();
 sg13g2_decap_8 FILLER_60_1331 ();
 sg13g2_decap_8 FILLER_60_1338 ();
 sg13g2_decap_8 FILLER_60_1345 ();
 sg13g2_decap_8 FILLER_60_1352 ();
 sg13g2_decap_4 FILLER_60_1359 ();
 sg13g2_fill_2 FILLER_60_1363 ();
 sg13g2_fill_1 FILLER_60_1369 ();
 sg13g2_decap_8 FILLER_60_1374 ();
 sg13g2_decap_8 FILLER_60_1441 ();
 sg13g2_decap_8 FILLER_60_1448 ();
 sg13g2_decap_8 FILLER_60_1455 ();
 sg13g2_decap_8 FILLER_60_1462 ();
 sg13g2_decap_8 FILLER_60_1469 ();
 sg13g2_decap_8 FILLER_60_1476 ();
 sg13g2_decap_8 FILLER_60_1483 ();
 sg13g2_fill_1 FILLER_60_1490 ();
 sg13g2_fill_1 FILLER_60_1500 ();
 sg13g2_fill_2 FILLER_60_1526 ();
 sg13g2_fill_1 FILLER_60_1585 ();
 sg13g2_decap_4 FILLER_60_1595 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_fill_2 FILLER_61_84 ();
 sg13g2_fill_1 FILLER_61_112 ();
 sg13g2_fill_2 FILLER_61_139 ();
 sg13g2_fill_1 FILLER_61_141 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_fill_2 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_181 ();
 sg13g2_decap_8 FILLER_61_188 ();
 sg13g2_decap_8 FILLER_61_195 ();
 sg13g2_decap_4 FILLER_61_202 ();
 sg13g2_fill_2 FILLER_61_206 ();
 sg13g2_decap_8 FILLER_61_229 ();
 sg13g2_decap_4 FILLER_61_236 ();
 sg13g2_fill_2 FILLER_61_240 ();
 sg13g2_fill_1 FILLER_61_246 ();
 sg13g2_fill_2 FILLER_61_252 ();
 sg13g2_fill_2 FILLER_61_258 ();
 sg13g2_fill_1 FILLER_61_265 ();
 sg13g2_decap_8 FILLER_61_274 ();
 sg13g2_decap_8 FILLER_61_281 ();
 sg13g2_decap_4 FILLER_61_288 ();
 sg13g2_fill_2 FILLER_61_292 ();
 sg13g2_decap_8 FILLER_61_298 ();
 sg13g2_decap_8 FILLER_61_305 ();
 sg13g2_decap_8 FILLER_61_312 ();
 sg13g2_decap_8 FILLER_61_319 ();
 sg13g2_decap_8 FILLER_61_326 ();
 sg13g2_decap_8 FILLER_61_333 ();
 sg13g2_decap_8 FILLER_61_344 ();
 sg13g2_decap_8 FILLER_61_351 ();
 sg13g2_decap_4 FILLER_61_358 ();
 sg13g2_decap_8 FILLER_61_366 ();
 sg13g2_decap_8 FILLER_61_373 ();
 sg13g2_decap_8 FILLER_61_380 ();
 sg13g2_decap_8 FILLER_61_387 ();
 sg13g2_fill_1 FILLER_61_394 ();
 sg13g2_fill_2 FILLER_61_420 ();
 sg13g2_decap_8 FILLER_61_436 ();
 sg13g2_fill_2 FILLER_61_464 ();
 sg13g2_fill_1 FILLER_61_466 ();
 sg13g2_decap_8 FILLER_61_496 ();
 sg13g2_fill_2 FILLER_61_503 ();
 sg13g2_decap_8 FILLER_61_510 ();
 sg13g2_decap_8 FILLER_61_517 ();
 sg13g2_decap_8 FILLER_61_524 ();
 sg13g2_decap_4 FILLER_61_531 ();
 sg13g2_fill_1 FILLER_61_535 ();
 sg13g2_decap_8 FILLER_61_541 ();
 sg13g2_decap_8 FILLER_61_548 ();
 sg13g2_decap_4 FILLER_61_555 ();
 sg13g2_fill_1 FILLER_61_559 ();
 sg13g2_decap_8 FILLER_61_589 ();
 sg13g2_decap_4 FILLER_61_596 ();
 sg13g2_decap_8 FILLER_61_605 ();
 sg13g2_decap_8 FILLER_61_612 ();
 sg13g2_fill_2 FILLER_61_619 ();
 sg13g2_fill_1 FILLER_61_621 ();
 sg13g2_decap_4 FILLER_61_631 ();
 sg13g2_decap_8 FILLER_61_639 ();
 sg13g2_decap_8 FILLER_61_646 ();
 sg13g2_fill_2 FILLER_61_653 ();
 sg13g2_fill_1 FILLER_61_690 ();
 sg13g2_decap_4 FILLER_61_695 ();
 sg13g2_fill_1 FILLER_61_699 ();
 sg13g2_decap_4 FILLER_61_705 ();
 sg13g2_fill_1 FILLER_61_709 ();
 sg13g2_decap_8 FILLER_61_731 ();
 sg13g2_decap_8 FILLER_61_738 ();
 sg13g2_fill_2 FILLER_61_745 ();
 sg13g2_fill_2 FILLER_61_752 ();
 sg13g2_fill_1 FILLER_61_754 ();
 sg13g2_decap_8 FILLER_61_819 ();
 sg13g2_decap_8 FILLER_61_830 ();
 sg13g2_decap_8 FILLER_61_837 ();
 sg13g2_decap_8 FILLER_61_844 ();
 sg13g2_decap_8 FILLER_61_851 ();
 sg13g2_decap_8 FILLER_61_858 ();
 sg13g2_decap_8 FILLER_61_865 ();
 sg13g2_decap_8 FILLER_61_872 ();
 sg13g2_decap_8 FILLER_61_879 ();
 sg13g2_decap_4 FILLER_61_886 ();
 sg13g2_fill_2 FILLER_61_890 ();
 sg13g2_decap_4 FILLER_61_897 ();
 sg13g2_decap_8 FILLER_61_905 ();
 sg13g2_fill_1 FILLER_61_912 ();
 sg13g2_decap_4 FILLER_61_960 ();
 sg13g2_decap_8 FILLER_61_990 ();
 sg13g2_decap_8 FILLER_61_997 ();
 sg13g2_decap_8 FILLER_61_1004 ();
 sg13g2_decap_8 FILLER_61_1011 ();
 sg13g2_fill_2 FILLER_61_1018 ();
 sg13g2_decap_4 FILLER_61_1035 ();
 sg13g2_decap_4 FILLER_61_1043 ();
 sg13g2_fill_1 FILLER_61_1047 ();
 sg13g2_fill_2 FILLER_61_1069 ();
 sg13g2_decap_8 FILLER_61_1118 ();
 sg13g2_decap_8 FILLER_61_1125 ();
 sg13g2_fill_2 FILLER_61_1132 ();
 sg13g2_fill_1 FILLER_61_1134 ();
 sg13g2_fill_1 FILLER_61_1156 ();
 sg13g2_decap_8 FILLER_61_1234 ();
 sg13g2_decap_8 FILLER_61_1241 ();
 sg13g2_fill_2 FILLER_61_1248 ();
 sg13g2_decap_4 FILLER_61_1281 ();
 sg13g2_fill_2 FILLER_61_1356 ();
 sg13g2_fill_2 FILLER_61_1384 ();
 sg13g2_fill_1 FILLER_61_1391 ();
 sg13g2_fill_2 FILLER_61_1426 ();
 sg13g2_fill_1 FILLER_61_1437 ();
 sg13g2_decap_4 FILLER_61_1463 ();
 sg13g2_fill_2 FILLER_61_1467 ();
 sg13g2_decap_8 FILLER_61_1474 ();
 sg13g2_decap_8 FILLER_61_1481 ();
 sg13g2_decap_8 FILLER_61_1488 ();
 sg13g2_decap_4 FILLER_61_1495 ();
 sg13g2_fill_2 FILLER_61_1554 ();
 sg13g2_fill_1 FILLER_61_1556 ();
 sg13g2_decap_8 FILLER_61_1592 ();
 sg13g2_decap_8 FILLER_61_1599 ();
 sg13g2_decap_8 FILLER_61_1606 ();
 sg13g2_decap_8 FILLER_61_1613 ();
 sg13g2_decap_4 FILLER_61_1620 ();
 sg13g2_fill_1 FILLER_61_1624 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_fill_1 FILLER_62_112 ();
 sg13g2_decap_4 FILLER_62_117 ();
 sg13g2_decap_4 FILLER_62_124 ();
 sg13g2_decap_8 FILLER_62_137 ();
 sg13g2_fill_1 FILLER_62_144 ();
 sg13g2_decap_8 FILLER_62_149 ();
 sg13g2_decap_8 FILLER_62_156 ();
 sg13g2_decap_8 FILLER_62_163 ();
 sg13g2_decap_8 FILLER_62_170 ();
 sg13g2_decap_8 FILLER_62_177 ();
 sg13g2_decap_8 FILLER_62_184 ();
 sg13g2_decap_4 FILLER_62_191 ();
 sg13g2_fill_1 FILLER_62_195 ();
 sg13g2_decap_4 FILLER_62_200 ();
 sg13g2_fill_1 FILLER_62_209 ();
 sg13g2_fill_2 FILLER_62_214 ();
 sg13g2_fill_1 FILLER_62_216 ();
 sg13g2_fill_2 FILLER_62_222 ();
 sg13g2_fill_2 FILLER_62_228 ();
 sg13g2_fill_1 FILLER_62_233 ();
 sg13g2_decap_8 FILLER_62_288 ();
 sg13g2_decap_8 FILLER_62_295 ();
 sg13g2_fill_1 FILLER_62_302 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_fill_2 FILLER_62_353 ();
 sg13g2_decap_8 FILLER_62_381 ();
 sg13g2_decap_8 FILLER_62_388 ();
 sg13g2_decap_8 FILLER_62_395 ();
 sg13g2_fill_2 FILLER_62_402 ();
 sg13g2_fill_1 FILLER_62_409 ();
 sg13g2_decap_4 FILLER_62_439 ();
 sg13g2_fill_2 FILLER_62_443 ();
 sg13g2_decap_4 FILLER_62_450 ();
 sg13g2_fill_2 FILLER_62_454 ();
 sg13g2_decap_4 FILLER_62_517 ();
 sg13g2_decap_4 FILLER_62_547 ();
 sg13g2_decap_4 FILLER_62_559 ();
 sg13g2_fill_2 FILLER_62_563 ();
 sg13g2_fill_1 FILLER_62_596 ();
 sg13g2_fill_2 FILLER_62_623 ();
 sg13g2_fill_1 FILLER_62_625 ();
 sg13g2_fill_2 FILLER_62_657 ();
 sg13g2_fill_1 FILLER_62_659 ();
 sg13g2_fill_2 FILLER_62_686 ();
 sg13g2_decap_8 FILLER_62_702 ();
 sg13g2_decap_4 FILLER_62_709 ();
 sg13g2_fill_2 FILLER_62_713 ();
 sg13g2_decap_8 FILLER_62_720 ();
 sg13g2_decap_4 FILLER_62_727 ();
 sg13g2_fill_2 FILLER_62_736 ();
 sg13g2_decap_8 FILLER_62_743 ();
 sg13g2_fill_1 FILLER_62_750 ();
 sg13g2_fill_2 FILLER_62_756 ();
 sg13g2_fill_2 FILLER_62_783 ();
 sg13g2_fill_1 FILLER_62_789 ();
 sg13g2_decap_8 FILLER_62_794 ();
 sg13g2_decap_8 FILLER_62_801 ();
 sg13g2_decap_8 FILLER_62_808 ();
 sg13g2_decap_4 FILLER_62_815 ();
 sg13g2_decap_4 FILLER_62_850 ();
 sg13g2_fill_1 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_860 ();
 sg13g2_decap_8 FILLER_62_865 ();
 sg13g2_decap_8 FILLER_62_872 ();
 sg13g2_fill_1 FILLER_62_939 ();
 sg13g2_decap_4 FILLER_62_966 ();
 sg13g2_fill_1 FILLER_62_970 ();
 sg13g2_decap_4 FILLER_62_992 ();
 sg13g2_fill_2 FILLER_62_996 ();
 sg13g2_fill_2 FILLER_62_1003 ();
 sg13g2_decap_8 FILLER_62_1009 ();
 sg13g2_decap_4 FILLER_62_1016 ();
 sg13g2_fill_2 FILLER_62_1020 ();
 sg13g2_decap_8 FILLER_62_1053 ();
 sg13g2_decap_8 FILLER_62_1060 ();
 sg13g2_decap_8 FILLER_62_1067 ();
 sg13g2_fill_1 FILLER_62_1078 ();
 sg13g2_fill_2 FILLER_62_1084 ();
 sg13g2_decap_8 FILLER_62_1111 ();
 sg13g2_decap_8 FILLER_62_1118 ();
 sg13g2_decap_8 FILLER_62_1125 ();
 sg13g2_fill_2 FILLER_62_1132 ();
 sg13g2_decap_8 FILLER_62_1155 ();
 sg13g2_fill_2 FILLER_62_1162 ();
 sg13g2_decap_8 FILLER_62_1168 ();
 sg13g2_decap_8 FILLER_62_1175 ();
 sg13g2_fill_1 FILLER_62_1182 ();
 sg13g2_decap_8 FILLER_62_1213 ();
 sg13g2_decap_8 FILLER_62_1220 ();
 sg13g2_decap_8 FILLER_62_1227 ();
 sg13g2_fill_1 FILLER_62_1234 ();
 sg13g2_decap_8 FILLER_62_1240 ();
 sg13g2_fill_2 FILLER_62_1247 ();
 sg13g2_fill_2 FILLER_62_1254 ();
 sg13g2_fill_1 FILLER_62_1256 ();
 sg13g2_fill_1 FILLER_62_1304 ();
 sg13g2_fill_2 FILLER_62_1352 ();
 sg13g2_decap_4 FILLER_62_1403 ();
 sg13g2_fill_1 FILLER_62_1407 ();
 sg13g2_fill_2 FILLER_62_1460 ();
 sg13g2_fill_1 FILLER_62_1462 ();
 sg13g2_fill_2 FILLER_62_1494 ();
 sg13g2_fill_2 FILLER_62_1522 ();
 sg13g2_fill_1 FILLER_62_1524 ();
 sg13g2_fill_1 FILLER_62_1546 ();
 sg13g2_fill_1 FILLER_62_1568 ();
 sg13g2_decap_8 FILLER_62_1595 ();
 sg13g2_decap_4 FILLER_62_1602 ();
 sg13g2_fill_2 FILLER_62_1606 ();
 sg13g2_decap_8 FILLER_62_1612 ();
 sg13g2_decap_4 FILLER_62_1619 ();
 sg13g2_fill_2 FILLER_62_1623 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_fill_2 FILLER_63_109 ();
 sg13g2_fill_1 FILLER_63_111 ();
 sg13g2_decap_8 FILLER_63_117 ();
 sg13g2_decap_8 FILLER_63_124 ();
 sg13g2_fill_1 FILLER_63_135 ();
 sg13g2_decap_4 FILLER_63_145 ();
 sg13g2_fill_1 FILLER_63_149 ();
 sg13g2_decap_4 FILLER_63_171 ();
 sg13g2_fill_2 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_181 ();
 sg13g2_fill_2 FILLER_63_188 ();
 sg13g2_decap_8 FILLER_63_242 ();
 sg13g2_decap_8 FILLER_63_249 ();
 sg13g2_decap_4 FILLER_63_256 ();
 sg13g2_fill_2 FILLER_63_290 ();
 sg13g2_fill_2 FILLER_63_297 ();
 sg13g2_decap_4 FILLER_63_303 ();
 sg13g2_fill_2 FILLER_63_307 ();
 sg13g2_decap_4 FILLER_63_330 ();
 sg13g2_decap_4 FILLER_63_338 ();
 sg13g2_fill_1 FILLER_63_342 ();
 sg13g2_decap_4 FILLER_63_352 ();
 sg13g2_decap_4 FILLER_63_365 ();
 sg13g2_decap_8 FILLER_63_374 ();
 sg13g2_decap_8 FILLER_63_381 ();
 sg13g2_decap_8 FILLER_63_388 ();
 sg13g2_decap_4 FILLER_63_395 ();
 sg13g2_fill_1 FILLER_63_399 ();
 sg13g2_decap_4 FILLER_63_404 ();
 sg13g2_decap_8 FILLER_63_439 ();
 sg13g2_decap_8 FILLER_63_446 ();
 sg13g2_decap_8 FILLER_63_453 ();
 sg13g2_decap_4 FILLER_63_460 ();
 sg13g2_fill_1 FILLER_63_464 ();
 sg13g2_fill_1 FILLER_63_469 ();
 sg13g2_decap_8 FILLER_63_491 ();
 sg13g2_decap_4 FILLER_63_498 ();
 sg13g2_fill_2 FILLER_63_502 ();
 sg13g2_decap_8 FILLER_63_508 ();
 sg13g2_decap_8 FILLER_63_515 ();
 sg13g2_fill_2 FILLER_63_522 ();
 sg13g2_fill_1 FILLER_63_524 ();
 sg13g2_decap_4 FILLER_63_572 ();
 sg13g2_fill_2 FILLER_63_576 ();
 sg13g2_decap_8 FILLER_63_582 ();
 sg13g2_decap_8 FILLER_63_589 ();
 sg13g2_decap_4 FILLER_63_596 ();
 sg13g2_decap_4 FILLER_63_608 ();
 sg13g2_fill_1 FILLER_63_612 ();
 sg13g2_fill_2 FILLER_63_652 ();
 sg13g2_fill_1 FILLER_63_654 ();
 sg13g2_decap_8 FILLER_63_659 ();
 sg13g2_decap_8 FILLER_63_666 ();
 sg13g2_decap_8 FILLER_63_673 ();
 sg13g2_decap_4 FILLER_63_680 ();
 sg13g2_decap_4 FILLER_63_714 ();
 sg13g2_fill_2 FILLER_63_718 ();
 sg13g2_fill_2 FILLER_63_767 ();
 sg13g2_fill_1 FILLER_63_769 ();
 sg13g2_decap_8 FILLER_63_809 ();
 sg13g2_decap_8 FILLER_63_816 ();
 sg13g2_fill_1 FILLER_63_852 ();
 sg13g2_fill_2 FILLER_63_879 ();
 sg13g2_fill_1 FILLER_63_881 ();
 sg13g2_fill_2 FILLER_63_907 ();
 sg13g2_fill_1 FILLER_63_909 ();
 sg13g2_decap_4 FILLER_63_919 ();
 sg13g2_fill_1 FILLER_63_923 ();
 sg13g2_fill_1 FILLER_63_929 ();
 sg13g2_decap_4 FILLER_63_942 ();
 sg13g2_fill_2 FILLER_63_946 ();
 sg13g2_decap_8 FILLER_63_951 ();
 sg13g2_decap_4 FILLER_63_958 ();
 sg13g2_fill_1 FILLER_63_962 ();
 sg13g2_decap_8 FILLER_63_967 ();
 sg13g2_decap_8 FILLER_63_974 ();
 sg13g2_decap_8 FILLER_63_981 ();
 sg13g2_decap_4 FILLER_63_988 ();
 sg13g2_decap_4 FILLER_63_1023 ();
 sg13g2_fill_1 FILLER_63_1027 ();
 sg13g2_decap_8 FILLER_63_1032 ();
 sg13g2_decap_8 FILLER_63_1039 ();
 sg13g2_decap_8 FILLER_63_1046 ();
 sg13g2_decap_8 FILLER_63_1053 ();
 sg13g2_decap_4 FILLER_63_1060 ();
 sg13g2_fill_2 FILLER_63_1064 ();
 sg13g2_decap_8 FILLER_63_1099 ();
 sg13g2_decap_4 FILLER_63_1106 ();
 sg13g2_fill_2 FILLER_63_1110 ();
 sg13g2_decap_4 FILLER_63_1117 ();
 sg13g2_fill_1 FILLER_63_1121 ();
 sg13g2_decap_8 FILLER_63_1160 ();
 sg13g2_decap_8 FILLER_63_1167 ();
 sg13g2_decap_8 FILLER_63_1174 ();
 sg13g2_decap_8 FILLER_63_1181 ();
 sg13g2_fill_2 FILLER_63_1188 ();
 sg13g2_decap_8 FILLER_63_1194 ();
 sg13g2_decap_8 FILLER_63_1201 ();
 sg13g2_decap_8 FILLER_63_1208 ();
 sg13g2_fill_2 FILLER_63_1228 ();
 sg13g2_fill_1 FILLER_63_1230 ();
 sg13g2_decap_8 FILLER_63_1257 ();
 sg13g2_decap_4 FILLER_63_1264 ();
 sg13g2_fill_1 FILLER_63_1268 ();
 sg13g2_decap_8 FILLER_63_1303 ();
 sg13g2_decap_8 FILLER_63_1310 ();
 sg13g2_decap_4 FILLER_63_1317 ();
 sg13g2_fill_2 FILLER_63_1321 ();
 sg13g2_decap_8 FILLER_63_1344 ();
 sg13g2_decap_8 FILLER_63_1351 ();
 sg13g2_decap_4 FILLER_63_1358 ();
 sg13g2_fill_2 FILLER_63_1380 ();
 sg13g2_decap_8 FILLER_63_1430 ();
 sg13g2_decap_8 FILLER_63_1437 ();
 sg13g2_decap_8 FILLER_63_1444 ();
 sg13g2_decap_8 FILLER_63_1461 ();
 sg13g2_fill_2 FILLER_63_1468 ();
 sg13g2_fill_1 FILLER_63_1470 ();
 sg13g2_decap_8 FILLER_63_1480 ();
 sg13g2_fill_2 FILLER_63_1487 ();
 sg13g2_decap_8 FILLER_63_1528 ();
 sg13g2_decap_8 FILLER_63_1535 ();
 sg13g2_fill_2 FILLER_63_1542 ();
 sg13g2_decap_8 FILLER_63_1549 ();
 sg13g2_fill_1 FILLER_63_1556 ();
 sg13g2_fill_2 FILLER_63_1567 ();
 sg13g2_decap_4 FILLER_63_1573 ();
 sg13g2_decap_4 FILLER_63_1581 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_4 FILLER_64_91 ();
 sg13g2_fill_2 FILLER_64_95 ();
 sg13g2_fill_1 FILLER_64_149 ();
 sg13g2_fill_2 FILLER_64_202 ();
 sg13g2_fill_1 FILLER_64_204 ();
 sg13g2_decap_4 FILLER_64_276 ();
 sg13g2_fill_2 FILLER_64_327 ();
 sg13g2_fill_2 FILLER_64_387 ();
 sg13g2_fill_2 FILLER_64_420 ();
 sg13g2_fill_2 FILLER_64_431 ();
 sg13g2_fill_1 FILLER_64_433 ();
 sg13g2_decap_4 FILLER_64_439 ();
 sg13g2_fill_1 FILLER_64_443 ();
 sg13g2_fill_1 FILLER_64_491 ();
 sg13g2_fill_1 FILLER_64_523 ();
 sg13g2_decap_8 FILLER_64_528 ();
 sg13g2_decap_8 FILLER_64_535 ();
 sg13g2_decap_8 FILLER_64_542 ();
 sg13g2_decap_8 FILLER_64_549 ();
 sg13g2_decap_8 FILLER_64_561 ();
 sg13g2_fill_2 FILLER_64_568 ();
 sg13g2_decap_8 FILLER_64_574 ();
 sg13g2_fill_2 FILLER_64_581 ();
 sg13g2_fill_2 FILLER_64_639 ();
 sg13g2_fill_1 FILLER_64_641 ();
 sg13g2_decap_8 FILLER_64_673 ();
 sg13g2_decap_8 FILLER_64_680 ();
 sg13g2_fill_2 FILLER_64_687 ();
 sg13g2_decap_8 FILLER_64_693 ();
 sg13g2_fill_2 FILLER_64_700 ();
 sg13g2_decap_8 FILLER_64_809 ();
 sg13g2_decap_8 FILLER_64_816 ();
 sg13g2_fill_2 FILLER_64_823 ();
 sg13g2_fill_1 FILLER_64_825 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_decap_8 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_950 ();
 sg13g2_fill_2 FILLER_64_994 ();
 sg13g2_decap_8 FILLER_64_1000 ();
 sg13g2_decap_8 FILLER_64_1007 ();
 sg13g2_decap_8 FILLER_64_1014 ();
 sg13g2_decap_8 FILLER_64_1021 ();
 sg13g2_decap_8 FILLER_64_1028 ();
 sg13g2_fill_1 FILLER_64_1035 ();
 sg13g2_decap_4 FILLER_64_1041 ();
 sg13g2_fill_1 FILLER_64_1045 ();
 sg13g2_decap_8 FILLER_64_1054 ();
 sg13g2_decap_4 FILLER_64_1061 ();
 sg13g2_fill_2 FILLER_64_1065 ();
 sg13g2_decap_8 FILLER_64_1093 ();
 sg13g2_decap_8 FILLER_64_1100 ();
 sg13g2_decap_4 FILLER_64_1107 ();
 sg13g2_fill_1 FILLER_64_1167 ();
 sg13g2_decap_4 FILLER_64_1172 ();
 sg13g2_fill_1 FILLER_64_1176 ();
 sg13g2_decap_8 FILLER_64_1186 ();
 sg13g2_decap_4 FILLER_64_1193 ();
 sg13g2_fill_1 FILLER_64_1197 ();
 sg13g2_decap_4 FILLER_64_1203 ();
 sg13g2_decap_4 FILLER_64_1233 ();
 sg13g2_fill_1 FILLER_64_1241 ();
 sg13g2_decap_4 FILLER_64_1247 ();
 sg13g2_fill_1 FILLER_64_1251 ();
 sg13g2_fill_2 FILLER_64_1256 ();
 sg13g2_decap_8 FILLER_64_1309 ();
 sg13g2_decap_8 FILLER_64_1316 ();
 sg13g2_decap_8 FILLER_64_1323 ();
 sg13g2_decap_4 FILLER_64_1330 ();
 sg13g2_fill_2 FILLER_64_1355 ();
 sg13g2_fill_1 FILLER_64_1357 ();
 sg13g2_fill_1 FILLER_64_1418 ();
 sg13g2_decap_8 FILLER_64_1423 ();
 sg13g2_decap_8 FILLER_64_1448 ();
 sg13g2_decap_8 FILLER_64_1455 ();
 sg13g2_decap_8 FILLER_64_1462 ();
 sg13g2_decap_8 FILLER_64_1469 ();
 sg13g2_decap_8 FILLER_64_1476 ();
 sg13g2_decap_8 FILLER_64_1483 ();
 sg13g2_decap_4 FILLER_64_1490 ();
 sg13g2_fill_2 FILLER_64_1498 ();
 sg13g2_fill_1 FILLER_64_1500 ();
 sg13g2_decap_4 FILLER_64_1506 ();
 sg13g2_fill_1 FILLER_64_1510 ();
 sg13g2_fill_2 FILLER_64_1516 ();
 sg13g2_fill_1 FILLER_64_1518 ();
 sg13g2_fill_2 FILLER_64_1523 ();
 sg13g2_fill_1 FILLER_64_1525 ();
 sg13g2_decap_8 FILLER_64_1531 ();
 sg13g2_decap_8 FILLER_64_1538 ();
 sg13g2_decap_8 FILLER_64_1545 ();
 sg13g2_decap_8 FILLER_64_1552 ();
 sg13g2_decap_8 FILLER_64_1559 ();
 sg13g2_fill_1 FILLER_64_1566 ();
 sg13g2_fill_1 FILLER_64_1588 ();
 sg13g2_decap_8 FILLER_64_1618 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_4 FILLER_65_98 ();
 sg13g2_fill_2 FILLER_65_102 ();
 sg13g2_fill_2 FILLER_65_133 ();
 sg13g2_fill_1 FILLER_65_135 ();
 sg13g2_decap_4 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_145 ();
 sg13g2_decap_8 FILLER_65_171 ();
 sg13g2_decap_8 FILLER_65_178 ();
 sg13g2_decap_8 FILLER_65_214 ();
 sg13g2_decap_4 FILLER_65_221 ();
 sg13g2_fill_1 FILLER_65_225 ();
 sg13g2_decap_4 FILLER_65_247 ();
 sg13g2_fill_2 FILLER_65_251 ();
 sg13g2_decap_8 FILLER_65_279 ();
 sg13g2_decap_8 FILLER_65_286 ();
 sg13g2_fill_2 FILLER_65_293 ();
 sg13g2_fill_1 FILLER_65_300 ();
 sg13g2_decap_4 FILLER_65_305 ();
 sg13g2_fill_1 FILLER_65_309 ();
 sg13g2_decap_8 FILLER_65_315 ();
 sg13g2_decap_8 FILLER_65_322 ();
 sg13g2_fill_2 FILLER_65_334 ();
 sg13g2_fill_1 FILLER_65_336 ();
 sg13g2_decap_8 FILLER_65_363 ();
 sg13g2_fill_1 FILLER_65_374 ();
 sg13g2_fill_2 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_403 ();
 sg13g2_decap_8 FILLER_65_443 ();
 sg13g2_fill_2 FILLER_65_450 ();
 sg13g2_decap_4 FILLER_65_456 ();
 sg13g2_fill_2 FILLER_65_460 ();
 sg13g2_decap_8 FILLER_65_472 ();
 sg13g2_decap_8 FILLER_65_479 ();
 sg13g2_decap_8 FILLER_65_486 ();
 sg13g2_decap_8 FILLER_65_493 ();
 sg13g2_decap_8 FILLER_65_500 ();
 sg13g2_decap_8 FILLER_65_507 ();
 sg13g2_decap_8 FILLER_65_514 ();
 sg13g2_fill_1 FILLER_65_521 ();
 sg13g2_fill_1 FILLER_65_527 ();
 sg13g2_decap_8 FILLER_65_536 ();
 sg13g2_fill_2 FILLER_65_543 ();
 sg13g2_fill_2 FILLER_65_550 ();
 sg13g2_fill_1 FILLER_65_552 ();
 sg13g2_fill_2 FILLER_65_584 ();
 sg13g2_fill_1 FILLER_65_586 ();
 sg13g2_decap_8 FILLER_65_608 ();
 sg13g2_decap_8 FILLER_65_615 ();
 sg13g2_decap_8 FILLER_65_622 ();
 sg13g2_decap_8 FILLER_65_629 ();
 sg13g2_decap_8 FILLER_65_636 ();
 sg13g2_decap_8 FILLER_65_643 ();
 sg13g2_decap_4 FILLER_65_650 ();
 sg13g2_decap_8 FILLER_65_658 ();
 sg13g2_decap_8 FILLER_65_665 ();
 sg13g2_decap_8 FILLER_65_672 ();
 sg13g2_fill_2 FILLER_65_679 ();
 sg13g2_fill_1 FILLER_65_715 ();
 sg13g2_decap_4 FILLER_65_723 ();
 sg13g2_fill_2 FILLER_65_727 ();
 sg13g2_fill_2 FILLER_65_778 ();
 sg13g2_fill_2 FILLER_65_785 ();
 sg13g2_decap_8 FILLER_65_822 ();
 sg13g2_decap_8 FILLER_65_829 ();
 sg13g2_decap_8 FILLER_65_836 ();
 sg13g2_decap_4 FILLER_65_843 ();
 sg13g2_decap_4 FILLER_65_911 ();
 sg13g2_fill_1 FILLER_65_915 ();
 sg13g2_fill_2 FILLER_65_950 ();
 sg13g2_decap_4 FILLER_65_978 ();
 sg13g2_decap_4 FILLER_65_1008 ();
 sg13g2_decap_4 FILLER_65_1017 ();
 sg13g2_decap_8 FILLER_65_1025 ();
 sg13g2_fill_2 FILLER_65_1037 ();
 sg13g2_decap_4 FILLER_65_1065 ();
 sg13g2_fill_1 FILLER_65_1069 ();
 sg13g2_decap_4 FILLER_65_1075 ();
 sg13g2_fill_1 FILLER_65_1079 ();
 sg13g2_decap_8 FILLER_65_1098 ();
 sg13g2_decap_8 FILLER_65_1105 ();
 sg13g2_decap_4 FILLER_65_1112 ();
 sg13g2_fill_1 FILLER_65_1116 ();
 sg13g2_decap_4 FILLER_65_1126 ();
 sg13g2_fill_1 FILLER_65_1130 ();
 sg13g2_decap_8 FILLER_65_1134 ();
 sg13g2_decap_8 FILLER_65_1141 ();
 sg13g2_decap_8 FILLER_65_1148 ();
 sg13g2_decap_8 FILLER_65_1155 ();
 sg13g2_decap_8 FILLER_65_1214 ();
 sg13g2_fill_2 FILLER_65_1221 ();
 sg13g2_fill_1 FILLER_65_1223 ();
 sg13g2_fill_2 FILLER_65_1249 ();
 sg13g2_decap_8 FILLER_65_1255 ();
 sg13g2_decap_8 FILLER_65_1262 ();
 sg13g2_decap_8 FILLER_65_1269 ();
 sg13g2_decap_4 FILLER_65_1276 ();
 sg13g2_fill_1 FILLER_65_1280 ();
 sg13g2_decap_8 FILLER_65_1295 ();
 sg13g2_decap_4 FILLER_65_1302 ();
 sg13g2_fill_2 FILLER_65_1306 ();
 sg13g2_decap_4 FILLER_65_1329 ();
 sg13g2_decap_8 FILLER_65_1354 ();
 sg13g2_fill_1 FILLER_65_1361 ();
 sg13g2_decap_8 FILLER_65_1366 ();
 sg13g2_decap_8 FILLER_65_1373 ();
 sg13g2_decap_8 FILLER_65_1380 ();
 sg13g2_decap_8 FILLER_65_1387 ();
 sg13g2_decap_4 FILLER_65_1394 ();
 sg13g2_fill_2 FILLER_65_1398 ();
 sg13g2_fill_1 FILLER_65_1405 ();
 sg13g2_decap_8 FILLER_65_1463 ();
 sg13g2_fill_2 FILLER_65_1470 ();
 sg13g2_fill_1 FILLER_65_1472 ();
 sg13g2_fill_1 FILLER_65_1478 ();
 sg13g2_fill_1 FILLER_65_1484 ();
 sg13g2_decap_4 FILLER_65_1537 ();
 sg13g2_fill_1 FILLER_65_1550 ();
 sg13g2_decap_8 FILLER_65_1555 ();
 sg13g2_decap_4 FILLER_65_1562 ();
 sg13g2_fill_2 FILLER_65_1566 ();
 sg13g2_fill_2 FILLER_65_1589 ();
 sg13g2_fill_1 FILLER_65_1591 ();
 sg13g2_fill_2 FILLER_65_1622 ();
 sg13g2_fill_1 FILLER_65_1624 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_4 FILLER_66_105 ();
 sg13g2_fill_1 FILLER_66_109 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_4 FILLER_66_175 ();
 sg13g2_fill_2 FILLER_66_179 ();
 sg13g2_decap_4 FILLER_66_185 ();
 sg13g2_fill_1 FILLER_66_194 ();
 sg13g2_fill_1 FILLER_66_204 ();
 sg13g2_fill_1 FILLER_66_226 ();
 sg13g2_decap_8 FILLER_66_253 ();
 sg13g2_decap_8 FILLER_66_260 ();
 sg13g2_decap_8 FILLER_66_267 ();
 sg13g2_decap_8 FILLER_66_274 ();
 sg13g2_decap_8 FILLER_66_281 ();
 sg13g2_decap_4 FILLER_66_314 ();
 sg13g2_fill_1 FILLER_66_318 ();
 sg13g2_fill_1 FILLER_66_362 ();
 sg13g2_decap_8 FILLER_66_384 ();
 sg13g2_decap_4 FILLER_66_420 ();
 sg13g2_fill_1 FILLER_66_424 ();
 sg13g2_decap_8 FILLER_66_446 ();
 sg13g2_decap_8 FILLER_66_453 ();
 sg13g2_fill_2 FILLER_66_460 ();
 sg13g2_fill_1 FILLER_66_462 ();
 sg13g2_decap_8 FILLER_66_468 ();
 sg13g2_decap_8 FILLER_66_475 ();
 sg13g2_decap_8 FILLER_66_482 ();
 sg13g2_decap_8 FILLER_66_493 ();
 sg13g2_fill_2 FILLER_66_500 ();
 sg13g2_decap_8 FILLER_66_506 ();
 sg13g2_fill_2 FILLER_66_513 ();
 sg13g2_fill_1 FILLER_66_515 ();
 sg13g2_decap_8 FILLER_66_547 ();
 sg13g2_decap_8 FILLER_66_554 ();
 sg13g2_fill_2 FILLER_66_561 ();
 sg13g2_fill_1 FILLER_66_563 ();
 sg13g2_decap_8 FILLER_66_568 ();
 sg13g2_decap_8 FILLER_66_575 ();
 sg13g2_decap_8 FILLER_66_582 ();
 sg13g2_decap_8 FILLER_66_589 ();
 sg13g2_decap_8 FILLER_66_596 ();
 sg13g2_decap_8 FILLER_66_603 ();
 sg13g2_decap_4 FILLER_66_610 ();
 sg13g2_fill_1 FILLER_66_645 ();
 sg13g2_fill_1 FILLER_66_667 ();
 sg13g2_fill_2 FILLER_66_694 ();
 sg13g2_fill_1 FILLER_66_696 ();
 sg13g2_fill_1 FILLER_66_772 ();
 sg13g2_fill_2 FILLER_66_799 ();
 sg13g2_fill_1 FILLER_66_801 ();
 sg13g2_fill_1 FILLER_66_822 ();
 sg13g2_decap_8 FILLER_66_832 ();
 sg13g2_fill_2 FILLER_66_839 ();
 sg13g2_fill_1 FILLER_66_867 ();
 sg13g2_fill_2 FILLER_66_893 ();
 sg13g2_fill_1 FILLER_66_895 ();
 sg13g2_fill_1 FILLER_66_957 ();
 sg13g2_decap_8 FILLER_66_996 ();
 sg13g2_decap_8 FILLER_66_1003 ();
 sg13g2_fill_1 FILLER_66_1010 ();
 sg13g2_decap_8 FILLER_66_1040 ();
 sg13g2_decap_8 FILLER_66_1082 ();
 sg13g2_fill_1 FILLER_66_1089 ();
 sg13g2_decap_4 FILLER_66_1116 ();
 sg13g2_fill_1 FILLER_66_1125 ();
 sg13g2_decap_4 FILLER_66_1134 ();
 sg13g2_fill_2 FILLER_66_1138 ();
 sg13g2_decap_4 FILLER_66_1145 ();
 sg13g2_fill_2 FILLER_66_1149 ();
 sg13g2_decap_4 FILLER_66_1155 ();
 sg13g2_fill_2 FILLER_66_1159 ();
 sg13g2_decap_8 FILLER_66_1186 ();
 sg13g2_decap_4 FILLER_66_1206 ();
 sg13g2_fill_2 FILLER_66_1210 ();
 sg13g2_decap_8 FILLER_66_1237 ();
 sg13g2_fill_1 FILLER_66_1244 ();
 sg13g2_decap_4 FILLER_66_1271 ();
 sg13g2_fill_1 FILLER_66_1275 ();
 sg13g2_decap_8 FILLER_66_1285 ();
 sg13g2_decap_8 FILLER_66_1292 ();
 sg13g2_decap_8 FILLER_66_1299 ();
 sg13g2_decap_8 FILLER_66_1306 ();
 sg13g2_decap_8 FILLER_66_1313 ();
 sg13g2_decap_8 FILLER_66_1320 ();
 sg13g2_decap_8 FILLER_66_1327 ();
 sg13g2_decap_8 FILLER_66_1334 ();
 sg13g2_fill_2 FILLER_66_1341 ();
 sg13g2_fill_1 FILLER_66_1343 ();
 sg13g2_decap_4 FILLER_66_1354 ();
 sg13g2_fill_2 FILLER_66_1367 ();
 sg13g2_decap_8 FILLER_66_1395 ();
 sg13g2_decap_8 FILLER_66_1402 ();
 sg13g2_decap_8 FILLER_66_1409 ();
 sg13g2_decap_8 FILLER_66_1416 ();
 sg13g2_decap_8 FILLER_66_1423 ();
 sg13g2_decap_8 FILLER_66_1430 ();
 sg13g2_fill_2 FILLER_66_1437 ();
 sg13g2_fill_1 FILLER_66_1439 ();
 sg13g2_decap_8 FILLER_66_1444 ();
 sg13g2_fill_2 FILLER_66_1451 ();
 sg13g2_fill_1 FILLER_66_1453 ();
 sg13g2_decap_8 FILLER_66_1468 ();
 sg13g2_decap_8 FILLER_66_1475 ();
 sg13g2_fill_1 FILLER_66_1482 ();
 sg13g2_decap_8 FILLER_66_1492 ();
 sg13g2_decap_8 FILLER_66_1499 ();
 sg13g2_decap_8 FILLER_66_1506 ();
 sg13g2_fill_2 FILLER_66_1513 ();
 sg13g2_decap_8 FILLER_66_1519 ();
 sg13g2_fill_2 FILLER_66_1531 ();
 sg13g2_decap_4 FILLER_66_1538 ();
 sg13g2_fill_1 FILLER_66_1542 ();
 sg13g2_decap_4 FILLER_66_1569 ();
 sg13g2_fill_1 FILLER_66_1573 ();
 sg13g2_decap_4 FILLER_66_1583 ();
 sg13g2_fill_1 FILLER_66_1587 ();
 sg13g2_fill_2 FILLER_66_1592 ();
 sg13g2_decap_8 FILLER_66_1599 ();
 sg13g2_decap_8 FILLER_66_1606 ();
 sg13g2_decap_8 FILLER_66_1613 ();
 sg13g2_decap_4 FILLER_66_1620 ();
 sg13g2_fill_1 FILLER_66_1624 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_4 FILLER_67_112 ();
 sg13g2_fill_1 FILLER_67_124 ();
 sg13g2_fill_2 FILLER_67_172 ();
 sg13g2_decap_8 FILLER_67_200 ();
 sg13g2_decap_8 FILLER_67_207 ();
 sg13g2_decap_8 FILLER_67_214 ();
 sg13g2_decap_8 FILLER_67_221 ();
 sg13g2_decap_8 FILLER_67_228 ();
 sg13g2_decap_8 FILLER_67_235 ();
 sg13g2_decap_8 FILLER_67_242 ();
 sg13g2_decap_8 FILLER_67_249 ();
 sg13g2_decap_4 FILLER_67_256 ();
 sg13g2_fill_1 FILLER_67_260 ();
 sg13g2_decap_4 FILLER_67_282 ();
 sg13g2_fill_2 FILLER_67_286 ();
 sg13g2_fill_2 FILLER_67_293 ();
 sg13g2_decap_8 FILLER_67_303 ();
 sg13g2_fill_2 FILLER_67_315 ();
 sg13g2_fill_2 FILLER_67_343 ();
 sg13g2_decap_4 FILLER_67_387 ();
 sg13g2_fill_1 FILLER_67_391 ();
 sg13g2_decap_8 FILLER_67_423 ();
 sg13g2_fill_2 FILLER_67_430 ();
 sg13g2_fill_1 FILLER_67_488 ();
 sg13g2_decap_8 FILLER_67_520 ();
 sg13g2_decap_8 FILLER_67_527 ();
 sg13g2_decap_4 FILLER_67_534 ();
 sg13g2_fill_2 FILLER_67_569 ();
 sg13g2_decap_4 FILLER_67_592 ();
 sg13g2_fill_1 FILLER_67_596 ();
 sg13g2_decap_8 FILLER_67_628 ();
 sg13g2_decap_8 FILLER_67_635 ();
 sg13g2_decap_4 FILLER_67_642 ();
 sg13g2_fill_1 FILLER_67_667 ();
 sg13g2_fill_2 FILLER_67_673 ();
 sg13g2_fill_1 FILLER_67_675 ();
 sg13g2_fill_2 FILLER_67_680 ();
 sg13g2_decap_4 FILLER_67_734 ();
 sg13g2_fill_2 FILLER_67_738 ();
 sg13g2_fill_2 FILLER_67_776 ();
 sg13g2_fill_2 FILLER_67_782 ();
 sg13g2_fill_1 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_825 ();
 sg13g2_fill_2 FILLER_67_832 ();
 sg13g2_fill_1 FILLER_67_834 ();
 sg13g2_decap_4 FILLER_67_886 ();
 sg13g2_fill_1 FILLER_67_890 ();
 sg13g2_decap_4 FILLER_67_896 ();
 sg13g2_decap_4 FILLER_67_908 ();
 sg13g2_fill_1 FILLER_67_912 ();
 sg13g2_fill_2 FILLER_67_1040 ();
 sg13g2_fill_1 FILLER_67_1042 ();
 sg13g2_decap_8 FILLER_67_1047 ();
 sg13g2_decap_8 FILLER_67_1054 ();
 sg13g2_decap_4 FILLER_67_1061 ();
 sg13g2_decap_8 FILLER_67_1091 ();
 sg13g2_fill_2 FILLER_67_1102 ();
 sg13g2_decap_8 FILLER_67_1109 ();
 sg13g2_fill_1 FILLER_67_1116 ();
 sg13g2_fill_2 FILLER_67_1169 ();
 sg13g2_decap_8 FILLER_67_1180 ();
 sg13g2_decap_4 FILLER_67_1187 ();
 sg13g2_fill_2 FILLER_67_1191 ();
 sg13g2_fill_2 FILLER_67_1239 ();
 sg13g2_fill_1 FILLER_67_1241 ();
 sg13g2_decap_8 FILLER_67_1251 ();
 sg13g2_fill_2 FILLER_67_1258 ();
 sg13g2_decap_4 FILLER_67_1264 ();
 sg13g2_decap_8 FILLER_67_1272 ();
 sg13g2_decap_8 FILLER_67_1305 ();
 sg13g2_decap_8 FILLER_67_1317 ();
 sg13g2_fill_2 FILLER_67_1324 ();
 sg13g2_decap_8 FILLER_67_1331 ();
 sg13g2_fill_2 FILLER_67_1338 ();
 sg13g2_fill_1 FILLER_67_1340 ();
 sg13g2_decap_8 FILLER_67_1354 ();
 sg13g2_decap_8 FILLER_67_1361 ();
 sg13g2_decap_4 FILLER_67_1368 ();
 sg13g2_fill_1 FILLER_67_1372 ();
 sg13g2_decap_8 FILLER_67_1402 ();
 sg13g2_decap_8 FILLER_67_1409 ();
 sg13g2_decap_8 FILLER_67_1416 ();
 sg13g2_decap_8 FILLER_67_1428 ();
 sg13g2_decap_8 FILLER_67_1435 ();
 sg13g2_fill_2 FILLER_67_1442 ();
 sg13g2_decap_8 FILLER_67_1485 ();
 sg13g2_fill_2 FILLER_67_1492 ();
 sg13g2_fill_1 FILLER_67_1494 ();
 sg13g2_fill_2 FILLER_67_1508 ();
 sg13g2_decap_4 FILLER_67_1514 ();
 sg13g2_fill_2 FILLER_67_1547 ();
 sg13g2_fill_2 FILLER_67_1578 ();
 sg13g2_fill_2 FILLER_67_1606 ();
 sg13g2_decap_8 FILLER_67_1612 ();
 sg13g2_decap_4 FILLER_67_1619 ();
 sg13g2_fill_2 FILLER_67_1623 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_4 FILLER_68_133 ();
 sg13g2_fill_1 FILLER_68_137 ();
 sg13g2_decap_8 FILLER_68_142 ();
 sg13g2_decap_4 FILLER_68_149 ();
 sg13g2_fill_2 FILLER_68_153 ();
 sg13g2_decap_8 FILLER_68_164 ();
 sg13g2_decap_4 FILLER_68_171 ();
 sg13g2_fill_1 FILLER_68_175 ();
 sg13g2_fill_2 FILLER_68_210 ();
 sg13g2_fill_1 FILLER_68_212 ();
 sg13g2_fill_1 FILLER_68_222 ();
 sg13g2_decap_8 FILLER_68_227 ();
 sg13g2_decap_8 FILLER_68_234 ();
 sg13g2_decap_8 FILLER_68_241 ();
 sg13g2_decap_8 FILLER_68_340 ();
 sg13g2_decap_8 FILLER_68_347 ();
 sg13g2_fill_2 FILLER_68_354 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_decap_4 FILLER_68_416 ();
 sg13g2_fill_1 FILLER_68_420 ();
 sg13g2_decap_8 FILLER_68_442 ();
 sg13g2_decap_8 FILLER_68_449 ();
 sg13g2_decap_4 FILLER_68_456 ();
 sg13g2_decap_8 FILLER_68_464 ();
 sg13g2_decap_8 FILLER_68_471 ();
 sg13g2_fill_1 FILLER_68_499 ();
 sg13g2_fill_1 FILLER_68_515 ();
 sg13g2_fill_1 FILLER_68_525 ();
 sg13g2_decap_4 FILLER_68_530 ();
 sg13g2_decap_8 FILLER_68_539 ();
 sg13g2_fill_2 FILLER_68_546 ();
 sg13g2_fill_1 FILLER_68_548 ();
 sg13g2_decap_4 FILLER_68_553 ();
 sg13g2_decap_4 FILLER_68_566 ();
 sg13g2_decap_8 FILLER_68_612 ();
 sg13g2_decap_8 FILLER_68_619 ();
 sg13g2_decap_8 FILLER_68_626 ();
 sg13g2_decap_8 FILLER_68_633 ();
 sg13g2_decap_8 FILLER_68_640 ();
 sg13g2_fill_2 FILLER_68_647 ();
 sg13g2_decap_8 FILLER_68_653 ();
 sg13g2_decap_4 FILLER_68_660 ();
 sg13g2_fill_1 FILLER_68_664 ();
 sg13g2_decap_8 FILLER_68_733 ();
 sg13g2_decap_8 FILLER_68_740 ();
 sg13g2_decap_8 FILLER_68_751 ();
 sg13g2_fill_1 FILLER_68_758 ();
 sg13g2_fill_2 FILLER_68_778 ();
 sg13g2_fill_1 FILLER_68_780 ();
 sg13g2_decap_8 FILLER_68_807 ();
 sg13g2_decap_8 FILLER_68_814 ();
 sg13g2_decap_4 FILLER_68_821 ();
 sg13g2_fill_1 FILLER_68_825 ();
 sg13g2_decap_8 FILLER_68_830 ();
 sg13g2_decap_8 FILLER_68_837 ();
 sg13g2_decap_8 FILLER_68_844 ();
 sg13g2_fill_1 FILLER_68_851 ();
 sg13g2_fill_2 FILLER_68_856 ();
 sg13g2_fill_1 FILLER_68_858 ();
 sg13g2_decap_4 FILLER_68_868 ();
 sg13g2_fill_1 FILLER_68_872 ();
 sg13g2_fill_1 FILLER_68_878 ();
 sg13g2_fill_2 FILLER_68_884 ();
 sg13g2_fill_1 FILLER_68_886 ();
 sg13g2_fill_2 FILLER_68_892 ();
 sg13g2_decap_4 FILLER_68_901 ();
 sg13g2_fill_2 FILLER_68_905 ();
 sg13g2_decap_8 FILLER_68_916 ();
 sg13g2_fill_2 FILLER_68_923 ();
 sg13g2_decap_8 FILLER_68_933 ();
 sg13g2_decap_4 FILLER_68_966 ();
 sg13g2_fill_2 FILLER_68_970 ();
 sg13g2_decap_8 FILLER_68_976 ();
 sg13g2_decap_8 FILLER_68_983 ();
 sg13g2_decap_4 FILLER_68_990 ();
 sg13g2_fill_2 FILLER_68_994 ();
 sg13g2_decap_4 FILLER_68_1000 ();
 sg13g2_fill_1 FILLER_68_1004 ();
 sg13g2_decap_4 FILLER_68_1031 ();
 sg13g2_fill_2 FILLER_68_1035 ();
 sg13g2_decap_8 FILLER_68_1063 ();
 sg13g2_decap_8 FILLER_68_1074 ();
 sg13g2_decap_4 FILLER_68_1081 ();
 sg13g2_decap_8 FILLER_68_1089 ();
 sg13g2_decap_4 FILLER_68_1096 ();
 sg13g2_fill_1 FILLER_68_1100 ();
 sg13g2_decap_8 FILLER_68_1132 ();
 sg13g2_fill_2 FILLER_68_1139 ();
 sg13g2_fill_1 FILLER_68_1141 ();
 sg13g2_decap_8 FILLER_68_1146 ();
 sg13g2_decap_8 FILLER_68_1153 ();
 sg13g2_fill_2 FILLER_68_1160 ();
 sg13g2_fill_1 FILLER_68_1162 ();
 sg13g2_decap_8 FILLER_68_1215 ();
 sg13g2_fill_2 FILLER_68_1222 ();
 sg13g2_decap_4 FILLER_68_1228 ();
 sg13g2_decap_8 FILLER_68_1241 ();
 sg13g2_fill_1 FILLER_68_1248 ();
 sg13g2_decap_8 FILLER_68_1279 ();
 sg13g2_fill_2 FILLER_68_1290 ();
 sg13g2_fill_1 FILLER_68_1292 ();
 sg13g2_decap_8 FILLER_68_1314 ();
 sg13g2_fill_1 FILLER_68_1321 ();
 sg13g2_decap_4 FILLER_68_1348 ();
 sg13g2_fill_2 FILLER_68_1352 ();
 sg13g2_decap_8 FILLER_68_1380 ();
 sg13g2_decap_8 FILLER_68_1387 ();
 sg13g2_fill_1 FILLER_68_1420 ();
 sg13g2_decap_4 FILLER_68_1426 ();
 sg13g2_decap_4 FILLER_68_1438 ();
 sg13g2_fill_1 FILLER_68_1442 ();
 sg13g2_fill_1 FILLER_68_1552 ();
 sg13g2_decap_8 FILLER_68_1579 ();
 sg13g2_decap_8 FILLER_68_1586 ();
 sg13g2_decap_4 FILLER_68_1593 ();
 sg13g2_fill_2 FILLER_68_1622 ();
 sg13g2_fill_1 FILLER_68_1624 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_fill_2 FILLER_69_126 ();
 sg13g2_fill_1 FILLER_69_128 ();
 sg13g2_decap_8 FILLER_69_155 ();
 sg13g2_fill_1 FILLER_69_162 ();
 sg13g2_decap_8 FILLER_69_168 ();
 sg13g2_fill_1 FILLER_69_175 ();
 sg13g2_fill_2 FILLER_69_183 ();
 sg13g2_decap_4 FILLER_69_211 ();
 sg13g2_fill_1 FILLER_69_215 ();
 sg13g2_fill_1 FILLER_69_242 ();
 sg13g2_decap_8 FILLER_69_269 ();
 sg13g2_decap_8 FILLER_69_276 ();
 sg13g2_decap_4 FILLER_69_283 ();
 sg13g2_fill_1 FILLER_69_313 ();
 sg13g2_fill_1 FILLER_69_321 ();
 sg13g2_fill_1 FILLER_69_326 ();
 sg13g2_decap_8 FILLER_69_331 ();
 sg13g2_decap_8 FILLER_69_367 ();
 sg13g2_decap_8 FILLER_69_374 ();
 sg13g2_decap_8 FILLER_69_381 ();
 sg13g2_fill_1 FILLER_69_388 ();
 sg13g2_decap_8 FILLER_69_453 ();
 sg13g2_decap_8 FILLER_69_460 ();
 sg13g2_decap_4 FILLER_69_467 ();
 sg13g2_fill_2 FILLER_69_471 ();
 sg13g2_fill_1 FILLER_69_483 ();
 sg13g2_fill_1 FILLER_69_516 ();
 sg13g2_decap_4 FILLER_69_543 ();
 sg13g2_decap_8 FILLER_69_579 ();
 sg13g2_decap_8 FILLER_69_586 ();
 sg13g2_decap_8 FILLER_69_593 ();
 sg13g2_decap_4 FILLER_69_621 ();
 sg13g2_fill_2 FILLER_69_625 ();
 sg13g2_decap_4 FILLER_69_670 ();
 sg13g2_fill_1 FILLER_69_707 ();
 sg13g2_fill_1 FILLER_69_734 ();
 sg13g2_fill_1 FILLER_69_740 ();
 sg13g2_fill_1 FILLER_69_747 ();
 sg13g2_fill_1 FILLER_69_752 ();
 sg13g2_fill_1 FILLER_69_813 ();
 sg13g2_decap_8 FILLER_69_848 ();
 sg13g2_decap_4 FILLER_69_855 ();
 sg13g2_fill_2 FILLER_69_864 ();
 sg13g2_fill_2 FILLER_69_874 ();
 sg13g2_fill_2 FILLER_69_881 ();
 sg13g2_decap_4 FILLER_69_888 ();
 sg13g2_decap_4 FILLER_69_897 ();
 sg13g2_decap_8 FILLER_69_906 ();
 sg13g2_decap_4 FILLER_69_916 ();
 sg13g2_fill_1 FILLER_69_920 ();
 sg13g2_decap_8 FILLER_69_951 ();
 sg13g2_decap_8 FILLER_69_958 ();
 sg13g2_decap_8 FILLER_69_965 ();
 sg13g2_decap_8 FILLER_69_972 ();
 sg13g2_fill_2 FILLER_69_979 ();
 sg13g2_fill_1 FILLER_69_985 ();
 sg13g2_fill_2 FILLER_69_1011 ();
 sg13g2_fill_2 FILLER_69_1017 ();
 sg13g2_fill_1 FILLER_69_1019 ();
 sg13g2_decap_8 FILLER_69_1024 ();
 sg13g2_decap_8 FILLER_69_1031 ();
 sg13g2_decap_4 FILLER_69_1038 ();
 sg13g2_decap_8 FILLER_69_1046 ();
 sg13g2_decap_8 FILLER_69_1053 ();
 sg13g2_decap_8 FILLER_69_1060 ();
 sg13g2_fill_1 FILLER_69_1067 ();
 sg13g2_decap_4 FILLER_69_1072 ();
 sg13g2_fill_1 FILLER_69_1076 ();
 sg13g2_fill_1 FILLER_69_1103 ();
 sg13g2_decap_8 FILLER_69_1133 ();
 sg13g2_decap_8 FILLER_69_1144 ();
 sg13g2_decap_8 FILLER_69_1151 ();
 sg13g2_decap_8 FILLER_69_1158 ();
 sg13g2_decap_4 FILLER_69_1165 ();
 sg13g2_decap_8 FILLER_69_1173 ();
 sg13g2_decap_8 FILLER_69_1180 ();
 sg13g2_decap_8 FILLER_69_1187 ();
 sg13g2_fill_2 FILLER_69_1194 ();
 sg13g2_decap_8 FILLER_69_1200 ();
 sg13g2_decap_8 FILLER_69_1207 ();
 sg13g2_fill_1 FILLER_69_1214 ();
 sg13g2_fill_2 FILLER_69_1246 ();
 sg13g2_fill_1 FILLER_69_1248 ();
 sg13g2_decap_8 FILLER_69_1285 ();
 sg13g2_fill_1 FILLER_69_1292 ();
 sg13g2_decap_4 FILLER_69_1319 ();
 sg13g2_decap_8 FILLER_69_1332 ();
 sg13g2_fill_2 FILLER_69_1339 ();
 sg13g2_decap_4 FILLER_69_1354 ();
 sg13g2_decap_8 FILLER_69_1366 ();
 sg13g2_fill_2 FILLER_69_1373 ();
 sg13g2_fill_1 FILLER_69_1375 ();
 sg13g2_decap_8 FILLER_69_1385 ();
 sg13g2_fill_2 FILLER_69_1392 ();
 sg13g2_fill_1 FILLER_69_1394 ();
 sg13g2_decap_4 FILLER_69_1404 ();
 sg13g2_fill_1 FILLER_69_1408 ();
 sg13g2_decap_8 FILLER_69_1413 ();
 sg13g2_fill_2 FILLER_69_1420 ();
 sg13g2_fill_1 FILLER_69_1422 ();
 sg13g2_decap_8 FILLER_69_1449 ();
 sg13g2_decap_8 FILLER_69_1456 ();
 sg13g2_decap_8 FILLER_69_1463 ();
 sg13g2_decap_8 FILLER_69_1470 ();
 sg13g2_decap_4 FILLER_69_1477 ();
 sg13g2_fill_2 FILLER_69_1481 ();
 sg13g2_decap_8 FILLER_69_1487 ();
 sg13g2_fill_2 FILLER_69_1494 ();
 sg13g2_decap_8 FILLER_69_1517 ();
 sg13g2_fill_2 FILLER_69_1524 ();
 sg13g2_fill_1 FILLER_69_1526 ();
 sg13g2_decap_8 FILLER_69_1531 ();
 sg13g2_decap_8 FILLER_69_1538 ();
 sg13g2_decap_8 FILLER_69_1545 ();
 sg13g2_fill_1 FILLER_69_1552 ();
 sg13g2_decap_4 FILLER_69_1556 ();
 sg13g2_fill_1 FILLER_69_1560 ();
 sg13g2_decap_8 FILLER_69_1570 ();
 sg13g2_decap_8 FILLER_69_1577 ();
 sg13g2_decap_4 FILLER_69_1584 ();
 sg13g2_fill_2 FILLER_69_1588 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_fill_2 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_135 ();
 sg13g2_decap_4 FILLER_70_204 ();
 sg13g2_fill_1 FILLER_70_208 ();
 sg13g2_decap_8 FILLER_70_213 ();
 sg13g2_fill_1 FILLER_70_245 ();
 sg13g2_decap_8 FILLER_70_272 ();
 sg13g2_decap_8 FILLER_70_279 ();
 sg13g2_decap_8 FILLER_70_286 ();
 sg13g2_decap_8 FILLER_70_297 ();
 sg13g2_decap_8 FILLER_70_304 ();
 sg13g2_fill_2 FILLER_70_373 ();
 sg13g2_fill_1 FILLER_70_427 ();
 sg13g2_fill_2 FILLER_70_454 ();
 sg13g2_fill_2 FILLER_70_477 ();
 sg13g2_fill_1 FILLER_70_505 ();
 sg13g2_decap_8 FILLER_70_527 ();
 sg13g2_decap_4 FILLER_70_534 ();
 sg13g2_fill_1 FILLER_70_538 ();
 sg13g2_decap_4 FILLER_70_543 ();
 sg13g2_decap_8 FILLER_70_573 ();
 sg13g2_fill_2 FILLER_70_580 ();
 sg13g2_fill_1 FILLER_70_582 ();
 sg13g2_decap_8 FILLER_70_587 ();
 sg13g2_decap_8 FILLER_70_594 ();
 sg13g2_decap_8 FILLER_70_601 ();
 sg13g2_decap_4 FILLER_70_608 ();
 sg13g2_fill_1 FILLER_70_612 ();
 sg13g2_decap_4 FILLER_70_643 ();
 sg13g2_decap_8 FILLER_70_714 ();
 sg13g2_fill_1 FILLER_70_721 ();
 sg13g2_fill_2 FILLER_70_735 ();
 sg13g2_fill_1 FILLER_70_741 ();
 sg13g2_fill_2 FILLER_70_802 ();
 sg13g2_decap_4 FILLER_70_814 ();
 sg13g2_fill_2 FILLER_70_818 ();
 sg13g2_fill_2 FILLER_70_845 ();
 sg13g2_fill_2 FILLER_70_856 ();
 sg13g2_fill_1 FILLER_70_858 ();
 sg13g2_decap_8 FILLER_70_885 ();
 sg13g2_decap_4 FILLER_70_892 ();
 sg13g2_fill_2 FILLER_70_912 ();
 sg13g2_decap_8 FILLER_70_924 ();
 sg13g2_decap_8 FILLER_70_931 ();
 sg13g2_decap_8 FILLER_70_938 ();
 sg13g2_decap_8 FILLER_70_945 ();
 sg13g2_decap_4 FILLER_70_952 ();
 sg13g2_decap_8 FILLER_70_960 ();
 sg13g2_decap_8 FILLER_70_967 ();
 sg13g2_decap_8 FILLER_70_1000 ();
 sg13g2_decap_8 FILLER_70_1007 ();
 sg13g2_decap_4 FILLER_70_1014 ();
 sg13g2_fill_2 FILLER_70_1018 ();
 sg13g2_decap_4 FILLER_70_1024 ();
 sg13g2_fill_2 FILLER_70_1031 ();
 sg13g2_fill_1 FILLER_70_1033 ();
 sg13g2_fill_2 FILLER_70_1060 ();
 sg13g2_decap_4 FILLER_70_1088 ();
 sg13g2_fill_1 FILLER_70_1092 ();
 sg13g2_decap_8 FILLER_70_1097 ();
 sg13g2_decap_8 FILLER_70_1104 ();
 sg13g2_decap_8 FILLER_70_1111 ();
 sg13g2_decap_8 FILLER_70_1118 ();
 sg13g2_decap_8 FILLER_70_1125 ();
 sg13g2_fill_1 FILLER_70_1132 ();
 sg13g2_decap_8 FILLER_70_1168 ();
 sg13g2_decap_8 FILLER_70_1175 ();
 sg13g2_decap_8 FILLER_70_1182 ();
 sg13g2_fill_2 FILLER_70_1189 ();
 sg13g2_fill_1 FILLER_70_1191 ();
 sg13g2_decap_8 FILLER_70_1196 ();
 sg13g2_decap_8 FILLER_70_1203 ();
 sg13g2_decap_8 FILLER_70_1210 ();
 sg13g2_fill_1 FILLER_70_1217 ();
 sg13g2_decap_8 FILLER_70_1256 ();
 sg13g2_decap_8 FILLER_70_1263 ();
 sg13g2_decap_8 FILLER_70_1270 ();
 sg13g2_decap_8 FILLER_70_1277 ();
 sg13g2_decap_8 FILLER_70_1284 ();
 sg13g2_decap_8 FILLER_70_1291 ();
 sg13g2_decap_8 FILLER_70_1298 ();
 sg13g2_decap_8 FILLER_70_1305 ();
 sg13g2_decap_8 FILLER_70_1312 ();
 sg13g2_decap_8 FILLER_70_1319 ();
 sg13g2_decap_4 FILLER_70_1326 ();
 sg13g2_fill_2 FILLER_70_1330 ();
 sg13g2_fill_2 FILLER_70_1360 ();
 sg13g2_fill_2 FILLER_70_1393 ();
 sg13g2_fill_1 FILLER_70_1395 ();
 sg13g2_decap_8 FILLER_70_1401 ();
 sg13g2_fill_1 FILLER_70_1408 ();
 sg13g2_decap_4 FILLER_70_1413 ();
 sg13g2_decap_8 FILLER_70_1522 ();
 sg13g2_decap_8 FILLER_70_1529 ();
 sg13g2_decap_8 FILLER_70_1536 ();
 sg13g2_decap_8 FILLER_70_1543 ();
 sg13g2_decap_4 FILLER_70_1550 ();
 sg13g2_fill_2 FILLER_70_1554 ();
 sg13g2_fill_2 FILLER_70_1561 ();
 sg13g2_fill_2 FILLER_70_1567 ();
 sg13g2_decap_8 FILLER_70_1590 ();
 sg13g2_decap_8 FILLER_70_1597 ();
 sg13g2_fill_2 FILLER_70_1604 ();
 sg13g2_fill_1 FILLER_70_1606 ();
 sg13g2_decap_8 FILLER_70_1611 ();
 sg13g2_decap_8 FILLER_70_1618 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_fill_1 FILLER_71_133 ();
 sg13g2_fill_2 FILLER_71_160 ();
 sg13g2_fill_1 FILLER_71_162 ();
 sg13g2_fill_2 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_220 ();
 sg13g2_fill_2 FILLER_71_227 ();
 sg13g2_fill_1 FILLER_71_229 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_decap_8 FILLER_71_266 ();
 sg13g2_decap_8 FILLER_71_304 ();
 sg13g2_fill_1 FILLER_71_311 ();
 sg13g2_fill_2 FILLER_71_317 ();
 sg13g2_fill_1 FILLER_71_319 ();
 sg13g2_fill_1 FILLER_71_345 ();
 sg13g2_decap_8 FILLER_71_367 ();
 sg13g2_decap_8 FILLER_71_374 ();
 sg13g2_decap_8 FILLER_71_381 ();
 sg13g2_fill_1 FILLER_71_393 ();
 sg13g2_decap_8 FILLER_71_424 ();
 sg13g2_fill_1 FILLER_71_431 ();
 sg13g2_decap_8 FILLER_71_436 ();
 sg13g2_decap_8 FILLER_71_443 ();
 sg13g2_decap_8 FILLER_71_450 ();
 sg13g2_fill_1 FILLER_71_457 ();
 sg13g2_decap_4 FILLER_71_463 ();
 sg13g2_fill_1 FILLER_71_467 ();
 sg13g2_decap_8 FILLER_71_473 ();
 sg13g2_decap_8 FILLER_71_480 ();
 sg13g2_decap_4 FILLER_71_487 ();
 sg13g2_decap_4 FILLER_71_496 ();
 sg13g2_fill_2 FILLER_71_504 ();
 sg13g2_fill_2 FILLER_71_527 ();
 sg13g2_fill_1 FILLER_71_554 ();
 sg13g2_decap_8 FILLER_71_559 ();
 sg13g2_decap_8 FILLER_71_601 ();
 sg13g2_decap_4 FILLER_71_608 ();
 sg13g2_fill_2 FILLER_71_612 ();
 sg13g2_decap_8 FILLER_71_619 ();
 sg13g2_decap_8 FILLER_71_630 ();
 sg13g2_fill_1 FILLER_71_637 ();
 sg13g2_fill_2 FILLER_71_647 ();
 sg13g2_decap_8 FILLER_71_653 ();
 sg13g2_decap_8 FILLER_71_664 ();
 sg13g2_decap_8 FILLER_71_671 ();
 sg13g2_decap_8 FILLER_71_678 ();
 sg13g2_decap_8 FILLER_71_685 ();
 sg13g2_decap_8 FILLER_71_692 ();
 sg13g2_fill_2 FILLER_71_699 ();
 sg13g2_decap_4 FILLER_71_711 ();
 sg13g2_decap_8 FILLER_71_719 ();
 sg13g2_decap_8 FILLER_71_726 ();
 sg13g2_decap_8 FILLER_71_733 ();
 sg13g2_decap_8 FILLER_71_746 ();
 sg13g2_decap_8 FILLER_71_757 ();
 sg13g2_decap_8 FILLER_71_764 ();
 sg13g2_decap_8 FILLER_71_771 ();
 sg13g2_decap_4 FILLER_71_778 ();
 sg13g2_fill_1 FILLER_71_782 ();
 sg13g2_fill_2 FILLER_71_787 ();
 sg13g2_fill_1 FILLER_71_789 ();
 sg13g2_fill_2 FILLER_71_794 ();
 sg13g2_decap_4 FILLER_71_825 ();
 sg13g2_fill_2 FILLER_71_829 ();
 sg13g2_fill_2 FILLER_71_857 ();
 sg13g2_fill_1 FILLER_71_859 ();
 sg13g2_decap_8 FILLER_71_885 ();
 sg13g2_fill_1 FILLER_71_892 ();
 sg13g2_fill_1 FILLER_71_913 ();
 sg13g2_decap_8 FILLER_71_920 ();
 sg13g2_decap_8 FILLER_71_927 ();
 sg13g2_decap_8 FILLER_71_934 ();
 sg13g2_decap_8 FILLER_71_941 ();
 sg13g2_fill_1 FILLER_71_948 ();
 sg13g2_decap_8 FILLER_71_975 ();
 sg13g2_decap_8 FILLER_71_982 ();
 sg13g2_fill_1 FILLER_71_989 ();
 sg13g2_fill_2 FILLER_71_994 ();
 sg13g2_decap_4 FILLER_71_1000 ();
 sg13g2_fill_2 FILLER_71_1009 ();
 sg13g2_fill_1 FILLER_71_1011 ();
 sg13g2_fill_2 FILLER_71_1043 ();
 sg13g2_decap_8 FILLER_71_1050 ();
 sg13g2_fill_2 FILLER_71_1057 ();
 sg13g2_fill_1 FILLER_71_1064 ();
 sg13g2_decap_8 FILLER_71_1108 ();
 sg13g2_decap_8 FILLER_71_1115 ();
 sg13g2_decap_8 FILLER_71_1122 ();
 sg13g2_decap_8 FILLER_71_1129 ();
 sg13g2_decap_4 FILLER_71_1136 ();
 sg13g2_fill_1 FILLER_71_1140 ();
 sg13g2_decap_4 FILLER_71_1147 ();
 sg13g2_fill_2 FILLER_71_1151 ();
 sg13g2_decap_4 FILLER_71_1156 ();
 sg13g2_decap_8 FILLER_71_1164 ();
 sg13g2_decap_8 FILLER_71_1171 ();
 sg13g2_fill_2 FILLER_71_1182 ();
 sg13g2_fill_1 FILLER_71_1184 ();
 sg13g2_fill_1 FILLER_71_1211 ();
 sg13g2_fill_2 FILLER_71_1238 ();
 sg13g2_fill_2 FILLER_71_1266 ();
 sg13g2_fill_2 FILLER_71_1278 ();
 sg13g2_fill_1 FILLER_71_1280 ();
 sg13g2_decap_4 FILLER_71_1302 ();
 sg13g2_fill_1 FILLER_71_1306 ();
 sg13g2_decap_4 FILLER_71_1312 ();
 sg13g2_fill_2 FILLER_71_1316 ();
 sg13g2_decap_8 FILLER_71_1323 ();
 sg13g2_decap_8 FILLER_71_1330 ();
 sg13g2_fill_1 FILLER_71_1337 ();
 sg13g2_fill_2 FILLER_71_1364 ();
 sg13g2_fill_1 FILLER_71_1366 ();
 sg13g2_decap_8 FILLER_71_1372 ();
 sg13g2_decap_8 FILLER_71_1379 ();
 sg13g2_decap_8 FILLER_71_1443 ();
 sg13g2_decap_8 FILLER_71_1450 ();
 sg13g2_decap_8 FILLER_71_1457 ();
 sg13g2_decap_4 FILLER_71_1464 ();
 sg13g2_decap_8 FILLER_71_1494 ();
 sg13g2_decap_4 FILLER_71_1501 ();
 sg13g2_decap_4 FILLER_71_1510 ();
 sg13g2_fill_1 FILLER_71_1514 ();
 sg13g2_decap_8 FILLER_71_1520 ();
 sg13g2_decap_8 FILLER_71_1527 ();
 sg13g2_decap_8 FILLER_71_1534 ();
 sg13g2_fill_2 FILLER_71_1541 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_fill_2 FILLER_72_133 ();
 sg13g2_fill_1 FILLER_72_135 ();
 sg13g2_decap_8 FILLER_72_190 ();
 sg13g2_decap_4 FILLER_72_197 ();
 sg13g2_decap_4 FILLER_72_274 ();
 sg13g2_fill_2 FILLER_72_299 ();
 sg13g2_decap_8 FILLER_72_311 ();
 sg13g2_decap_8 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_fill_2 FILLER_72_385 ();
 sg13g2_fill_1 FILLER_72_392 ();
 sg13g2_fill_2 FILLER_72_409 ();
 sg13g2_decap_4 FILLER_72_420 ();
 sg13g2_fill_1 FILLER_72_424 ();
 sg13g2_decap_4 FILLER_72_429 ();
 sg13g2_fill_2 FILLER_72_454 ();
 sg13g2_fill_1 FILLER_72_456 ();
 sg13g2_decap_8 FILLER_72_461 ();
 sg13g2_decap_8 FILLER_72_468 ();
 sg13g2_fill_1 FILLER_72_475 ();
 sg13g2_decap_8 FILLER_72_480 ();
 sg13g2_fill_1 FILLER_72_487 ();
 sg13g2_decap_8 FILLER_72_493 ();
 sg13g2_decap_8 FILLER_72_500 ();
 sg13g2_decap_8 FILLER_72_507 ();
 sg13g2_decap_8 FILLER_72_514 ();
 sg13g2_fill_1 FILLER_72_521 ();
 sg13g2_fill_2 FILLER_72_557 ();
 sg13g2_decap_8 FILLER_72_573 ();
 sg13g2_decap_8 FILLER_72_580 ();
 sg13g2_decap_8 FILLER_72_587 ();
 sg13g2_decap_8 FILLER_72_594 ();
 sg13g2_decap_8 FILLER_72_605 ();
 sg13g2_fill_2 FILLER_72_612 ();
 sg13g2_fill_1 FILLER_72_614 ();
 sg13g2_decap_8 FILLER_72_619 ();
 sg13g2_decap_8 FILLER_72_626 ();
 sg13g2_decap_8 FILLER_72_633 ();
 sg13g2_fill_1 FILLER_72_640 ();
 sg13g2_decap_8 FILLER_72_667 ();
 sg13g2_fill_2 FILLER_72_674 ();
 sg13g2_fill_1 FILLER_72_676 ();
 sg13g2_fill_1 FILLER_72_706 ();
 sg13g2_decap_8 FILLER_72_745 ();
 sg13g2_decap_8 FILLER_72_752 ();
 sg13g2_fill_2 FILLER_72_759 ();
 sg13g2_fill_1 FILLER_72_761 ();
 sg13g2_decap_8 FILLER_72_766 ();
 sg13g2_decap_8 FILLER_72_773 ();
 sg13g2_decap_8 FILLER_72_780 ();
 sg13g2_decap_8 FILLER_72_787 ();
 sg13g2_decap_8 FILLER_72_794 ();
 sg13g2_decap_8 FILLER_72_801 ();
 sg13g2_fill_2 FILLER_72_808 ();
 sg13g2_fill_1 FILLER_72_810 ();
 sg13g2_decap_8 FILLER_72_816 ();
 sg13g2_decap_8 FILLER_72_823 ();
 sg13g2_decap_8 FILLER_72_830 ();
 sg13g2_decap_8 FILLER_72_837 ();
 sg13g2_decap_8 FILLER_72_844 ();
 sg13g2_decap_8 FILLER_72_851 ();
 sg13g2_fill_1 FILLER_72_858 ();
 sg13g2_decap_8 FILLER_72_890 ();
 sg13g2_decap_8 FILLER_72_897 ();
 sg13g2_fill_1 FILLER_72_904 ();
 sg13g2_decap_4 FILLER_72_913 ();
 sg13g2_fill_2 FILLER_72_917 ();
 sg13g2_decap_8 FILLER_72_923 ();
 sg13g2_decap_4 FILLER_72_930 ();
 sg13g2_fill_2 FILLER_72_934 ();
 sg13g2_decap_4 FILLER_72_950 ();
 sg13g2_fill_1 FILLER_72_954 ();
 sg13g2_decap_4 FILLER_72_961 ();
 sg13g2_fill_1 FILLER_72_965 ();
 sg13g2_fill_2 FILLER_72_970 ();
 sg13g2_decap_8 FILLER_72_975 ();
 sg13g2_decap_8 FILLER_72_982 ();
 sg13g2_fill_2 FILLER_72_994 ();
 sg13g2_decap_4 FILLER_72_1004 ();
 sg13g2_fill_2 FILLER_72_1012 ();
 sg13g2_fill_1 FILLER_72_1014 ();
 sg13g2_decap_4 FILLER_72_1024 ();
 sg13g2_decap_8 FILLER_72_1058 ();
 sg13g2_decap_4 FILLER_72_1094 ();
 sg13g2_fill_2 FILLER_72_1118 ();
 sg13g2_fill_2 FILLER_72_1130 ();
 sg13g2_fill_1 FILLER_72_1132 ();
 sg13g2_decap_4 FILLER_72_1166 ();
 sg13g2_fill_1 FILLER_72_1175 ();
 sg13g2_decap_8 FILLER_72_1180 ();
 sg13g2_fill_2 FILLER_72_1187 ();
 sg13g2_fill_1 FILLER_72_1189 ();
 sg13g2_decap_8 FILLER_72_1219 ();
 sg13g2_decap_8 FILLER_72_1226 ();
 sg13g2_decap_8 FILLER_72_1233 ();
 sg13g2_fill_2 FILLER_72_1240 ();
 sg13g2_fill_1 FILLER_72_1242 ();
 sg13g2_decap_8 FILLER_72_1247 ();
 sg13g2_fill_1 FILLER_72_1280 ();
 sg13g2_fill_1 FILLER_72_1302 ();
 sg13g2_fill_2 FILLER_72_1334 ();
 sg13g2_fill_2 FILLER_72_1357 ();
 sg13g2_fill_1 FILLER_72_1359 ();
 sg13g2_fill_2 FILLER_72_1365 ();
 sg13g2_fill_1 FILLER_72_1367 ();
 sg13g2_decap_8 FILLER_72_1372 ();
 sg13g2_decap_4 FILLER_72_1379 ();
 sg13g2_fill_1 FILLER_72_1383 ();
 sg13g2_decap_4 FILLER_72_1409 ();
 sg13g2_fill_2 FILLER_72_1413 ();
 sg13g2_fill_2 FILLER_72_1420 ();
 sg13g2_fill_2 FILLER_72_1430 ();
 sg13g2_fill_1 FILLER_72_1432 ();
 sg13g2_fill_1 FILLER_72_1437 ();
 sg13g2_decap_8 FILLER_72_1459 ();
 sg13g2_decap_8 FILLER_72_1466 ();
 sg13g2_fill_2 FILLER_72_1473 ();
 sg13g2_decap_8 FILLER_72_1479 ();
 sg13g2_decap_8 FILLER_72_1486 ();
 sg13g2_decap_8 FILLER_72_1493 ();
 sg13g2_decap_8 FILLER_72_1500 ();
 sg13g2_decap_8 FILLER_72_1507 ();
 sg13g2_decap_4 FILLER_72_1514 ();
 sg13g2_fill_1 FILLER_72_1518 ();
 sg13g2_decap_8 FILLER_72_1540 ();
 sg13g2_fill_2 FILLER_72_1547 ();
 sg13g2_fill_1 FILLER_72_1549 ();
 sg13g2_decap_8 FILLER_72_1554 ();
 sg13g2_decap_8 FILLER_72_1561 ();
 sg13g2_decap_8 FILLER_72_1568 ();
 sg13g2_decap_8 FILLER_72_1575 ();
 sg13g2_decap_8 FILLER_72_1582 ();
 sg13g2_decap_4 FILLER_72_1589 ();
 sg13g2_fill_1 FILLER_72_1593 ();
 sg13g2_decap_8 FILLER_72_1599 ();
 sg13g2_fill_1 FILLER_72_1606 ();
 sg13g2_decap_8 FILLER_72_1611 ();
 sg13g2_decap_8 FILLER_72_1618 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_fill_2 FILLER_73_144 ();
 sg13g2_fill_1 FILLER_73_146 ();
 sg13g2_decap_4 FILLER_73_201 ();
 sg13g2_fill_2 FILLER_73_249 ();
 sg13g2_decap_8 FILLER_73_260 ();
 sg13g2_fill_1 FILLER_73_267 ();
 sg13g2_decap_8 FILLER_73_272 ();
 sg13g2_fill_2 FILLER_73_279 ();
 sg13g2_fill_1 FILLER_73_281 ();
 sg13g2_decap_8 FILLER_73_311 ();
 sg13g2_decap_4 FILLER_73_318 ();
 sg13g2_fill_1 FILLER_73_322 ();
 sg13g2_fill_2 FILLER_73_327 ();
 sg13g2_fill_2 FILLER_73_350 ();
 sg13g2_decap_8 FILLER_73_362 ();
 sg13g2_decap_4 FILLER_73_374 ();
 sg13g2_fill_1 FILLER_73_378 ();
 sg13g2_fill_2 FILLER_73_456 ();
 sg13g2_fill_2 FILLER_73_494 ();
 sg13g2_fill_2 FILLER_73_501 ();
 sg13g2_decap_8 FILLER_73_507 ();
 sg13g2_decap_8 FILLER_73_514 ();
 sg13g2_fill_2 FILLER_73_530 ();
 sg13g2_decap_8 FILLER_73_536 ();
 sg13g2_decap_8 FILLER_73_543 ();
 sg13g2_decap_8 FILLER_73_550 ();
 sg13g2_fill_1 FILLER_73_557 ();
 sg13g2_decap_4 FILLER_73_584 ();
 sg13g2_fill_2 FILLER_73_588 ();
 sg13g2_decap_8 FILLER_73_633 ();
 sg13g2_decap_8 FILLER_73_640 ();
 sg13g2_decap_8 FILLER_73_647 ();
 sg13g2_decap_8 FILLER_73_654 ();
 sg13g2_decap_8 FILLER_73_661 ();
 sg13g2_decap_8 FILLER_73_668 ();
 sg13g2_decap_8 FILLER_73_709 ();
 sg13g2_decap_4 FILLER_73_716 ();
 sg13g2_fill_1 FILLER_73_720 ();
 sg13g2_decap_8 FILLER_73_726 ();
 sg13g2_decap_8 FILLER_73_733 ();
 sg13g2_decap_8 FILLER_73_740 ();
 sg13g2_fill_2 FILLER_73_747 ();
 sg13g2_fill_1 FILLER_73_749 ();
 sg13g2_fill_1 FILLER_73_755 ();
 sg13g2_fill_1 FILLER_73_786 ();
 sg13g2_fill_1 FILLER_73_807 ();
 sg13g2_decap_4 FILLER_73_817 ();
 sg13g2_fill_1 FILLER_73_821 ();
 sg13g2_decap_4 FILLER_73_832 ();
 sg13g2_fill_2 FILLER_73_841 ();
 sg13g2_fill_1 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_848 ();
 sg13g2_decap_8 FILLER_73_855 ();
 sg13g2_fill_2 FILLER_73_862 ();
 sg13g2_decap_8 FILLER_73_877 ();
 sg13g2_decap_8 FILLER_73_899 ();
 sg13g2_decap_8 FILLER_73_906 ();
 sg13g2_fill_1 FILLER_73_918 ();
 sg13g2_decap_4 FILLER_73_933 ();
 sg13g2_decap_4 FILLER_73_941 ();
 sg13g2_fill_1 FILLER_73_959 ();
 sg13g2_fill_1 FILLER_73_965 ();
 sg13g2_fill_1 FILLER_73_977 ();
 sg13g2_decap_8 FILLER_73_982 ();
 sg13g2_fill_2 FILLER_73_989 ();
 sg13g2_fill_2 FILLER_73_1014 ();
 sg13g2_fill_1 FILLER_73_1016 ();
 sg13g2_fill_1 FILLER_73_1026 ();
 sg13g2_fill_1 FILLER_73_1032 ();
 sg13g2_fill_2 FILLER_73_1047 ();
 sg13g2_fill_2 FILLER_73_1058 ();
 sg13g2_fill_1 FILLER_73_1070 ();
 sg13g2_fill_2 FILLER_73_1075 ();
 sg13g2_fill_2 FILLER_73_1091 ();
 sg13g2_fill_1 FILLER_73_1093 ();
 sg13g2_decap_8 FILLER_73_1106 ();
 sg13g2_decap_8 FILLER_73_1113 ();
 sg13g2_fill_1 FILLER_73_1120 ();
 sg13g2_fill_2 FILLER_73_1126 ();
 sg13g2_fill_1 FILLER_73_1149 ();
 sg13g2_fill_1 FILLER_73_1175 ();
 sg13g2_fill_1 FILLER_73_1181 ();
 sg13g2_fill_2 FILLER_73_1220 ();
 sg13g2_decap_8 FILLER_73_1226 ();
 sg13g2_fill_2 FILLER_73_1247 ();
 sg13g2_fill_1 FILLER_73_1249 ();
 sg13g2_decap_4 FILLER_73_1259 ();
 sg13g2_decap_8 FILLER_73_1267 ();
 sg13g2_decap_8 FILLER_73_1279 ();
 sg13g2_decap_8 FILLER_73_1286 ();
 sg13g2_decap_8 FILLER_73_1293 ();
 sg13g2_fill_2 FILLER_73_1300 ();
 sg13g2_fill_2 FILLER_73_1333 ();
 sg13g2_fill_1 FILLER_73_1335 ();
 sg13g2_fill_2 FILLER_73_1387 ();
 sg13g2_fill_2 FILLER_73_1397 ();
 sg13g2_fill_1 FILLER_73_1399 ();
 sg13g2_fill_1 FILLER_73_1404 ();
 sg13g2_decap_8 FILLER_73_1430 ();
 sg13g2_fill_1 FILLER_73_1437 ();
 sg13g2_fill_2 FILLER_73_1464 ();
 sg13g2_fill_1 FILLER_73_1466 ();
 sg13g2_decap_4 FILLER_73_1472 ();
 sg13g2_fill_2 FILLER_73_1476 ();
 sg13g2_decap_8 FILLER_73_1482 ();
 sg13g2_fill_2 FILLER_73_1489 ();
 sg13g2_fill_1 FILLER_73_1491 ();
 sg13g2_fill_2 FILLER_73_1501 ();
 sg13g2_decap_8 FILLER_73_1507 ();
 sg13g2_decap_8 FILLER_73_1514 ();
 sg13g2_fill_2 FILLER_73_1521 ();
 sg13g2_decap_4 FILLER_73_1544 ();
 sg13g2_fill_2 FILLER_73_1548 ();
 sg13g2_decap_8 FILLER_73_1554 ();
 sg13g2_decap_8 FILLER_73_1561 ();
 sg13g2_fill_2 FILLER_73_1568 ();
 sg13g2_fill_2 FILLER_73_1591 ();
 sg13g2_fill_1 FILLER_73_1593 ();
 sg13g2_fill_1 FILLER_73_1598 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_fill_2 FILLER_74_154 ();
 sg13g2_fill_1 FILLER_74_156 ();
 sg13g2_fill_2 FILLER_74_161 ();
 sg13g2_fill_2 FILLER_74_201 ();
 sg13g2_fill_1 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_326 ();
 sg13g2_fill_2 FILLER_74_333 ();
 sg13g2_fill_1 FILLER_74_335 ();
 sg13g2_decap_8 FILLER_74_413 ();
 sg13g2_decap_8 FILLER_74_420 ();
 sg13g2_fill_2 FILLER_74_427 ();
 sg13g2_fill_2 FILLER_74_438 ();
 sg13g2_decap_4 FILLER_74_449 ();
 sg13g2_decap_4 FILLER_74_484 ();
 sg13g2_fill_2 FILLER_74_488 ();
 sg13g2_decap_4 FILLER_74_519 ();
 sg13g2_fill_1 FILLER_74_523 ();
 sg13g2_fill_2 FILLER_74_550 ();
 sg13g2_decap_8 FILLER_74_556 ();
 sg13g2_fill_2 FILLER_74_563 ();
 sg13g2_decap_8 FILLER_74_569 ();
 sg13g2_decap_8 FILLER_74_576 ();
 sg13g2_fill_2 FILLER_74_583 ();
 sg13g2_decap_8 FILLER_74_615 ();
 sg13g2_decap_8 FILLER_74_622 ();
 sg13g2_fill_1 FILLER_74_629 ();
 sg13g2_decap_8 FILLER_74_639 ();
 sg13g2_decap_8 FILLER_74_646 ();
 sg13g2_decap_8 FILLER_74_653 ();
 sg13g2_fill_2 FILLER_74_660 ();
 sg13g2_fill_1 FILLER_74_662 ();
 sg13g2_decap_8 FILLER_74_668 ();
 sg13g2_decap_4 FILLER_74_681 ();
 sg13g2_fill_1 FILLER_74_685 ();
 sg13g2_fill_1 FILLER_74_696 ();
 sg13g2_decap_8 FILLER_74_708 ();
 sg13g2_fill_1 FILLER_74_715 ();
 sg13g2_fill_1 FILLER_74_726 ();
 sg13g2_decap_8 FILLER_74_730 ();
 sg13g2_fill_1 FILLER_74_737 ();
 sg13g2_decap_8 FILLER_74_752 ();
 sg13g2_fill_2 FILLER_74_759 ();
 sg13g2_fill_2 FILLER_74_771 ();
 sg13g2_fill_1 FILLER_74_789 ();
 sg13g2_fill_2 FILLER_74_795 ();
 sg13g2_fill_1 FILLER_74_805 ();
 sg13g2_fill_1 FILLER_74_810 ();
 sg13g2_fill_1 FILLER_74_820 ();
 sg13g2_fill_2 FILLER_74_831 ();
 sg13g2_fill_2 FILLER_74_839 ();
 sg13g2_fill_1 FILLER_74_841 ();
 sg13g2_fill_2 FILLER_74_848 ();
 sg13g2_fill_1 FILLER_74_850 ();
 sg13g2_fill_2 FILLER_74_859 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_fill_2 FILLER_74_866 ();
 sg13g2_fill_1 FILLER_74_868 ();
 sg13g2_fill_2 FILLER_74_884 ();
 sg13g2_decap_4 FILLER_74_891 ();
 sg13g2_fill_2 FILLER_74_900 ();
 sg13g2_fill_1 FILLER_74_902 ();
 sg13g2_fill_2 FILLER_74_917 ();
 sg13g2_fill_1 FILLER_74_919 ();
 sg13g2_decap_8 FILLER_74_925 ();
 sg13g2_decap_8 FILLER_74_932 ();
 sg13g2_decap_8 FILLER_74_962 ();
 sg13g2_decap_4 FILLER_74_969 ();
 sg13g2_fill_2 FILLER_74_973 ();
 sg13g2_fill_1 FILLER_74_980 ();
 sg13g2_fill_2 FILLER_74_989 ();
 sg13g2_fill_2 FILLER_74_996 ();
 sg13g2_fill_2 FILLER_74_1002 ();
 sg13g2_fill_1 FILLER_74_1004 ();
 sg13g2_fill_2 FILLER_74_1010 ();
 sg13g2_decap_8 FILLER_74_1017 ();
 sg13g2_decap_8 FILLER_74_1024 ();
 sg13g2_decap_8 FILLER_74_1031 ();
 sg13g2_decap_8 FILLER_74_1038 ();
 sg13g2_fill_2 FILLER_74_1045 ();
 sg13g2_fill_1 FILLER_74_1047 ();
 sg13g2_decap_4 FILLER_74_1079 ();
 sg13g2_fill_2 FILLER_74_1088 ();
 sg13g2_fill_1 FILLER_74_1090 ();
 sg13g2_decap_8 FILLER_74_1105 ();
 sg13g2_decap_8 FILLER_74_1124 ();
 sg13g2_decap_8 FILLER_74_1131 ();
 sg13g2_decap_8 FILLER_74_1138 ();
 sg13g2_fill_2 FILLER_74_1145 ();
 sg13g2_decap_4 FILLER_74_1162 ();
 sg13g2_fill_1 FILLER_74_1166 ();
 sg13g2_decap_8 FILLER_74_1171 ();
 sg13g2_decap_8 FILLER_74_1178 ();
 sg13g2_decap_8 FILLER_74_1185 ();
 sg13g2_decap_8 FILLER_74_1192 ();
 sg13g2_decap_8 FILLER_74_1199 ();
 sg13g2_decap_4 FILLER_74_1211 ();
 sg13g2_fill_1 FILLER_74_1215 ();
 sg13g2_fill_1 FILLER_74_1242 ();
 sg13g2_decap_8 FILLER_74_1247 ();
 sg13g2_decap_4 FILLER_74_1254 ();
 sg13g2_fill_1 FILLER_74_1258 ();
 sg13g2_decap_8 FILLER_74_1287 ();
 sg13g2_decap_8 FILLER_74_1294 ();
 sg13g2_decap_8 FILLER_74_1301 ();
 sg13g2_decap_8 FILLER_74_1308 ();
 sg13g2_fill_2 FILLER_74_1315 ();
 sg13g2_fill_1 FILLER_74_1317 ();
 sg13g2_decap_8 FILLER_74_1328 ();
 sg13g2_decap_8 FILLER_74_1335 ();
 sg13g2_decap_8 FILLER_74_1342 ();
 sg13g2_decap_8 FILLER_74_1349 ();
 sg13g2_fill_2 FILLER_74_1356 ();
 sg13g2_fill_1 FILLER_74_1358 ();
 sg13g2_decap_4 FILLER_74_1362 ();
 sg13g2_fill_1 FILLER_74_1366 ();
 sg13g2_decap_8 FILLER_74_1372 ();
 sg13g2_fill_2 FILLER_74_1379 ();
 sg13g2_fill_2 FILLER_74_1412 ();
 sg13g2_decap_8 FILLER_74_1440 ();
 sg13g2_decap_8 FILLER_74_1447 ();
 sg13g2_fill_2 FILLER_74_1454 ();
 sg13g2_fill_1 FILLER_74_1456 ();
 sg13g2_decap_4 FILLER_74_1530 ();
 sg13g2_fill_1 FILLER_74_1534 ();
 sg13g2_fill_2 FILLER_74_1566 ();
 sg13g2_fill_1 FILLER_74_1568 ();
 sg13g2_decap_4 FILLER_74_1590 ();
 sg13g2_fill_2 FILLER_74_1594 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_4 FILLER_75_202 ();
 sg13g2_fill_2 FILLER_75_206 ();
 sg13g2_fill_1 FILLER_75_234 ();
 sg13g2_fill_1 FILLER_75_244 ();
 sg13g2_fill_2 FILLER_75_249 ();
 sg13g2_decap_8 FILLER_75_258 ();
 sg13g2_decap_8 FILLER_75_265 ();
 sg13g2_decap_8 FILLER_75_272 ();
 sg13g2_decap_8 FILLER_75_279 ();
 sg13g2_decap_8 FILLER_75_286 ();
 sg13g2_decap_8 FILLER_75_293 ();
 sg13g2_decap_8 FILLER_75_300 ();
 sg13g2_decap_8 FILLER_75_307 ();
 sg13g2_decap_8 FILLER_75_314 ();
 sg13g2_decap_8 FILLER_75_321 ();
 sg13g2_fill_1 FILLER_75_328 ();
 sg13g2_decap_8 FILLER_75_362 ();
 sg13g2_fill_2 FILLER_75_369 ();
 sg13g2_fill_1 FILLER_75_371 ();
 sg13g2_decap_4 FILLER_75_381 ();
 sg13g2_fill_1 FILLER_75_385 ();
 sg13g2_fill_2 FILLER_75_391 ();
 sg13g2_fill_1 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_403 ();
 sg13g2_decap_4 FILLER_75_410 ();
 sg13g2_fill_2 FILLER_75_414 ();
 sg13g2_fill_1 FILLER_75_441 ();
 sg13g2_decap_8 FILLER_75_467 ();
 sg13g2_decap_8 FILLER_75_474 ();
 sg13g2_fill_2 FILLER_75_485 ();
 sg13g2_decap_8 FILLER_75_520 ();
 sg13g2_decap_8 FILLER_75_527 ();
 sg13g2_decap_4 FILLER_75_534 ();
 sg13g2_fill_1 FILLER_75_538 ();
 sg13g2_decap_4 FILLER_75_543 ();
 sg13g2_fill_1 FILLER_75_577 ();
 sg13g2_decap_8 FILLER_75_586 ();
 sg13g2_decap_8 FILLER_75_593 ();
 sg13g2_fill_1 FILLER_75_600 ();
 sg13g2_decap_4 FILLER_75_652 ();
 sg13g2_fill_1 FILLER_75_656 ();
 sg13g2_fill_2 FILLER_75_671 ();
 sg13g2_decap_4 FILLER_75_677 ();
 sg13g2_fill_2 FILLER_75_693 ();
 sg13g2_fill_1 FILLER_75_695 ();
 sg13g2_fill_1 FILLER_75_700 ();
 sg13g2_fill_2 FILLER_75_709 ();
 sg13g2_fill_1 FILLER_75_711 ();
 sg13g2_fill_1 FILLER_75_723 ();
 sg13g2_decap_8 FILLER_75_728 ();
 sg13g2_decap_8 FILLER_75_735 ();
 sg13g2_fill_2 FILLER_75_742 ();
 sg13g2_fill_2 FILLER_75_753 ();
 sg13g2_fill_2 FILLER_75_759 ();
 sg13g2_decap_4 FILLER_75_766 ();
 sg13g2_fill_2 FILLER_75_770 ();
 sg13g2_decap_4 FILLER_75_777 ();
 sg13g2_fill_1 FILLER_75_781 ();
 sg13g2_decap_8 FILLER_75_787 ();
 sg13g2_decap_8 FILLER_75_794 ();
 sg13g2_fill_2 FILLER_75_801 ();
 sg13g2_fill_1 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_825 ();
 sg13g2_decap_4 FILLER_75_832 ();
 sg13g2_decap_8 FILLER_75_841 ();
 sg13g2_fill_1 FILLER_75_848 ();
 sg13g2_decap_8 FILLER_75_859 ();
 sg13g2_decap_8 FILLER_75_866 ();
 sg13g2_decap_8 FILLER_75_873 ();
 sg13g2_fill_1 FILLER_75_880 ();
 sg13g2_fill_1 FILLER_75_885 ();
 sg13g2_decap_8 FILLER_75_890 ();
 sg13g2_decap_4 FILLER_75_897 ();
 sg13g2_fill_2 FILLER_75_901 ();
 sg13g2_fill_2 FILLER_75_908 ();
 sg13g2_decap_8 FILLER_75_914 ();
 sg13g2_decap_8 FILLER_75_925 ();
 sg13g2_fill_1 FILLER_75_932 ();
 sg13g2_decap_8 FILLER_75_959 ();
 sg13g2_decap_8 FILLER_75_966 ();
 sg13g2_decap_8 FILLER_75_973 ();
 sg13g2_decap_8 FILLER_75_980 ();
 sg13g2_decap_8 FILLER_75_987 ();
 sg13g2_fill_1 FILLER_75_994 ();
 sg13g2_decap_4 FILLER_75_999 ();
 sg13g2_fill_2 FILLER_75_1003 ();
 sg13g2_fill_1 FILLER_75_1020 ();
 sg13g2_decap_4 FILLER_75_1025 ();
 sg13g2_fill_1 FILLER_75_1029 ();
 sg13g2_decap_4 FILLER_75_1044 ();
 sg13g2_fill_1 FILLER_75_1048 ();
 sg13g2_fill_2 FILLER_75_1083 ();
 sg13g2_fill_1 FILLER_75_1085 ();
 sg13g2_decap_4 FILLER_75_1100 ();
 sg13g2_fill_2 FILLER_75_1108 ();
 sg13g2_decap_8 FILLER_75_1136 ();
 sg13g2_decap_8 FILLER_75_1143 ();
 sg13g2_decap_8 FILLER_75_1150 ();
 sg13g2_decap_8 FILLER_75_1157 ();
 sg13g2_fill_2 FILLER_75_1164 ();
 sg13g2_fill_1 FILLER_75_1166 ();
 sg13g2_decap_8 FILLER_75_1180 ();
 sg13g2_decap_8 FILLER_75_1187 ();
 sg13g2_decap_4 FILLER_75_1194 ();
 sg13g2_fill_1 FILLER_75_1198 ();
 sg13g2_decap_8 FILLER_75_1209 ();
 sg13g2_decap_8 FILLER_75_1216 ();
 sg13g2_decap_8 FILLER_75_1223 ();
 sg13g2_fill_1 FILLER_75_1230 ();
 sg13g2_fill_2 FILLER_75_1234 ();
 sg13g2_fill_1 FILLER_75_1262 ();
 sg13g2_fill_2 FILLER_75_1272 ();
 sg13g2_decap_4 FILLER_75_1283 ();
 sg13g2_fill_1 FILLER_75_1287 ();
 sg13g2_decap_8 FILLER_75_1309 ();
 sg13g2_fill_2 FILLER_75_1316 ();
 sg13g2_fill_1 FILLER_75_1318 ();
 sg13g2_decap_8 FILLER_75_1334 ();
 sg13g2_decap_8 FILLER_75_1341 ();
 sg13g2_fill_2 FILLER_75_1348 ();
 sg13g2_fill_1 FILLER_75_1384 ();
 sg13g2_decap_8 FILLER_75_1389 ();
 sg13g2_fill_2 FILLER_75_1396 ();
 sg13g2_decap_8 FILLER_75_1402 ();
 sg13g2_decap_8 FILLER_75_1409 ();
 sg13g2_fill_2 FILLER_75_1416 ();
 sg13g2_decap_8 FILLER_75_1422 ();
 sg13g2_decap_8 FILLER_75_1429 ();
 sg13g2_fill_1 FILLER_75_1436 ();
 sg13g2_decap_8 FILLER_75_1458 ();
 sg13g2_fill_1 FILLER_75_1465 ();
 sg13g2_fill_1 FILLER_75_1470 ();
 sg13g2_decap_4 FILLER_75_1500 ();
 sg13g2_fill_2 FILLER_75_1504 ();
 sg13g2_decap_8 FILLER_75_1527 ();
 sg13g2_decap_8 FILLER_75_1534 ();
 sg13g2_fill_2 FILLER_75_1541 ();
 sg13g2_decap_4 FILLER_75_1585 ();
 sg13g2_fill_1 FILLER_75_1589 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_fill_2 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_201 ();
 sg13g2_decap_8 FILLER_76_208 ();
 sg13g2_decap_4 FILLER_76_215 ();
 sg13g2_fill_2 FILLER_76_219 ();
 sg13g2_fill_1 FILLER_76_231 ();
 sg13g2_fill_2 FILLER_76_267 ();
 sg13g2_fill_1 FILLER_76_269 ();
 sg13g2_fill_2 FILLER_76_274 ();
 sg13g2_fill_1 FILLER_76_276 ();
 sg13g2_decap_8 FILLER_76_281 ();
 sg13g2_decap_8 FILLER_76_288 ();
 sg13g2_fill_1 FILLER_76_295 ();
 sg13g2_fill_1 FILLER_76_305 ();
 sg13g2_decap_8 FILLER_76_310 ();
 sg13g2_decap_4 FILLER_76_317 ();
 sg13g2_decap_4 FILLER_76_351 ();
 sg13g2_decap_4 FILLER_76_368 ();
 sg13g2_fill_1 FILLER_76_372 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_4 FILLER_76_409 ();
 sg13g2_fill_1 FILLER_76_413 ();
 sg13g2_fill_2 FILLER_76_440 ();
 sg13g2_decap_8 FILLER_76_472 ();
 sg13g2_fill_2 FILLER_76_479 ();
 sg13g2_fill_1 FILLER_76_486 ();
 sg13g2_decap_8 FILLER_76_513 ();
 sg13g2_decap_8 FILLER_76_520 ();
 sg13g2_decap_8 FILLER_76_527 ();
 sg13g2_decap_4 FILLER_76_534 ();
 sg13g2_fill_1 FILLER_76_538 ();
 sg13g2_decap_4 FILLER_76_596 ();
 sg13g2_decap_8 FILLER_76_604 ();
 sg13g2_decap_8 FILLER_76_611 ();
 sg13g2_decap_8 FILLER_76_618 ();
 sg13g2_decap_8 FILLER_76_625 ();
 sg13g2_fill_1 FILLER_76_661 ();
 sg13g2_decap_4 FILLER_76_678 ();
 sg13g2_fill_2 FILLER_76_701 ();
 sg13g2_fill_1 FILLER_76_703 ();
 sg13g2_decap_4 FILLER_76_709 ();
 sg13g2_fill_1 FILLER_76_713 ();
 sg13g2_decap_8 FILLER_76_724 ();
 sg13g2_fill_2 FILLER_76_736 ();
 sg13g2_fill_1 FILLER_76_748 ();
 sg13g2_decap_8 FILLER_76_753 ();
 sg13g2_fill_2 FILLER_76_760 ();
 sg13g2_fill_1 FILLER_76_771 ();
 sg13g2_decap_8 FILLER_76_781 ();
 sg13g2_decap_4 FILLER_76_788 ();
 sg13g2_decap_4 FILLER_76_796 ();
 sg13g2_decap_8 FILLER_76_809 ();
 sg13g2_decap_4 FILLER_76_816 ();
 sg13g2_fill_2 FILLER_76_820 ();
 sg13g2_decap_8 FILLER_76_827 ();
 sg13g2_fill_2 FILLER_76_834 ();
 sg13g2_fill_1 FILLER_76_836 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_4 FILLER_76_849 ();
 sg13g2_decap_8 FILLER_76_862 ();
 sg13g2_fill_2 FILLER_76_869 ();
 sg13g2_decap_8 FILLER_76_875 ();
 sg13g2_decap_8 FILLER_76_882 ();
 sg13g2_decap_8 FILLER_76_889 ();
 sg13g2_decap_8 FILLER_76_896 ();
 sg13g2_fill_1 FILLER_76_903 ();
 sg13g2_decap_8 FILLER_76_959 ();
 sg13g2_decap_8 FILLER_76_966 ();
 sg13g2_decap_4 FILLER_76_973 ();
 sg13g2_decap_8 FILLER_76_986 ();
 sg13g2_decap_8 FILLER_76_993 ();
 sg13g2_decap_8 FILLER_76_1000 ();
 sg13g2_fill_2 FILLER_76_1007 ();
 sg13g2_decap_8 FILLER_76_1021 ();
 sg13g2_fill_2 FILLER_76_1028 ();
 sg13g2_fill_2 FILLER_76_1040 ();
 sg13g2_fill_1 FILLER_76_1042 ();
 sg13g2_fill_2 FILLER_76_1093 ();
 sg13g2_fill_1 FILLER_76_1095 ();
 sg13g2_fill_2 FILLER_76_1108 ();
 sg13g2_fill_1 FILLER_76_1115 ();
 sg13g2_decap_8 FILLER_76_1126 ();
 sg13g2_fill_1 FILLER_76_1133 ();
 sg13g2_decap_4 FILLER_76_1139 ();
 sg13g2_fill_1 FILLER_76_1143 ();
 sg13g2_decap_8 FILLER_76_1148 ();
 sg13g2_decap_4 FILLER_76_1155 ();
 sg13g2_fill_1 FILLER_76_1159 ();
 sg13g2_fill_1 FILLER_76_1186 ();
 sg13g2_decap_8 FILLER_76_1209 ();
 sg13g2_decap_8 FILLER_76_1216 ();
 sg13g2_decap_8 FILLER_76_1223 ();
 sg13g2_fill_1 FILLER_76_1230 ();
 sg13g2_decap_4 FILLER_76_1256 ();
 sg13g2_fill_2 FILLER_76_1286 ();
 sg13g2_fill_2 FILLER_76_1309 ();
 sg13g2_fill_1 FILLER_76_1311 ();
 sg13g2_decap_8 FILLER_76_1316 ();
 sg13g2_decap_8 FILLER_76_1323 ();
 sg13g2_decap_8 FILLER_76_1330 ();
 sg13g2_fill_1 FILLER_76_1337 ();
 sg13g2_decap_8 FILLER_76_1373 ();
 sg13g2_decap_4 FILLER_76_1380 ();
 sg13g2_fill_1 FILLER_76_1384 ();
 sg13g2_fill_1 FILLER_76_1416 ();
 sg13g2_decap_4 FILLER_76_1422 ();
 sg13g2_decap_4 FILLER_76_1430 ();
 sg13g2_decap_8 FILLER_76_1438 ();
 sg13g2_decap_8 FILLER_76_1445 ();
 sg13g2_decap_8 FILLER_76_1452 ();
 sg13g2_decap_8 FILLER_76_1459 ();
 sg13g2_fill_1 FILLER_76_1501 ();
 sg13g2_decap_8 FILLER_76_1542 ();
 sg13g2_decap_4 FILLER_76_1549 ();
 sg13g2_fill_2 FILLER_76_1579 ();
 sg13g2_fill_1 FILLER_76_1581 ();
 sg13g2_decap_8 FILLER_76_1586 ();
 sg13g2_decap_8 FILLER_76_1593 ();
 sg13g2_decap_8 FILLER_76_1600 ();
 sg13g2_decap_8 FILLER_76_1607 ();
 sg13g2_decap_8 FILLER_76_1614 ();
 sg13g2_decap_4 FILLER_76_1621 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_fill_2 FILLER_77_154 ();
 sg13g2_fill_1 FILLER_77_156 ();
 sg13g2_decap_4 FILLER_77_191 ();
 sg13g2_fill_2 FILLER_77_195 ();
 sg13g2_decap_4 FILLER_77_202 ();
 sg13g2_fill_1 FILLER_77_206 ();
 sg13g2_fill_2 FILLER_77_211 ();
 sg13g2_decap_4 FILLER_77_346 ();
 sg13g2_fill_2 FILLER_77_350 ();
 sg13g2_fill_1 FILLER_77_378 ();
 sg13g2_fill_2 FILLER_77_431 ();
 sg13g2_fill_1 FILLER_77_459 ();
 sg13g2_decap_8 FILLER_77_481 ();
 sg13g2_decap_8 FILLER_77_488 ();
 sg13g2_decap_8 FILLER_77_495 ();
 sg13g2_decap_8 FILLER_77_502 ();
 sg13g2_decap_4 FILLER_77_509 ();
 sg13g2_fill_2 FILLER_77_513 ();
 sg13g2_decap_8 FILLER_77_540 ();
 sg13g2_decap_8 FILLER_77_547 ();
 sg13g2_decap_8 FILLER_77_554 ();
 sg13g2_decap_4 FILLER_77_561 ();
 sg13g2_decap_8 FILLER_77_619 ();
 sg13g2_decap_4 FILLER_77_626 ();
 sg13g2_fill_1 FILLER_77_644 ();
 sg13g2_fill_1 FILLER_77_671 ();
 sg13g2_decap_4 FILLER_77_682 ();
 sg13g2_decap_8 FILLER_77_690 ();
 sg13g2_decap_8 FILLER_77_697 ();
 sg13g2_decap_8 FILLER_77_704 ();
 sg13g2_decap_8 FILLER_77_716 ();
 sg13g2_decap_8 FILLER_77_723 ();
 sg13g2_decap_8 FILLER_77_730 ();
 sg13g2_decap_4 FILLER_77_737 ();
 sg13g2_fill_2 FILLER_77_741 ();
 sg13g2_decap_8 FILLER_77_769 ();
 sg13g2_decap_8 FILLER_77_776 ();
 sg13g2_fill_2 FILLER_77_783 ();
 sg13g2_fill_1 FILLER_77_785 ();
 sg13g2_decap_8 FILLER_77_812 ();
 sg13g2_fill_2 FILLER_77_845 ();
 sg13g2_fill_1 FILLER_77_847 ();
 sg13g2_fill_1 FILLER_77_856 ();
 sg13g2_fill_1 FILLER_77_888 ();
 sg13g2_fill_2 FILLER_77_899 ();
 sg13g2_decap_8 FILLER_77_907 ();
 sg13g2_decap_8 FILLER_77_914 ();
 sg13g2_decap_8 FILLER_77_921 ();
 sg13g2_fill_1 FILLER_77_928 ();
 sg13g2_fill_2 FILLER_77_967 ();
 sg13g2_fill_2 FILLER_77_973 ();
 sg13g2_fill_1 FILLER_77_975 ();
 sg13g2_decap_8 FILLER_77_981 ();
 sg13g2_fill_2 FILLER_77_988 ();
 sg13g2_decap_4 FILLER_77_1009 ();
 sg13g2_decap_4 FILLER_77_1017 ();
 sg13g2_fill_1 FILLER_77_1033 ();
 sg13g2_fill_2 FILLER_77_1038 ();
 sg13g2_fill_1 FILLER_77_1040 ();
 sg13g2_decap_4 FILLER_77_1046 ();
 sg13g2_fill_2 FILLER_77_1050 ();
 sg13g2_fill_2 FILLER_77_1060 ();
 sg13g2_fill_1 FILLER_77_1062 ();
 sg13g2_decap_8 FILLER_77_1157 ();
 sg13g2_decap_4 FILLER_77_1164 ();
 sg13g2_fill_2 FILLER_77_1168 ();
 sg13g2_decap_8 FILLER_77_1180 ();
 sg13g2_fill_2 FILLER_77_1187 ();
 sg13g2_fill_2 FILLER_77_1209 ();
 sg13g2_fill_1 FILLER_77_1211 ();
 sg13g2_fill_2 FILLER_77_1220 ();
 sg13g2_fill_1 FILLER_77_1222 ();
 sg13g2_decap_8 FILLER_77_1229 ();
 sg13g2_decap_8 FILLER_77_1236 ();
 sg13g2_fill_1 FILLER_77_1243 ();
 sg13g2_decap_8 FILLER_77_1250 ();
 sg13g2_decap_8 FILLER_77_1257 ();
 sg13g2_fill_2 FILLER_77_1264 ();
 sg13g2_decap_8 FILLER_77_1270 ();
 sg13g2_fill_2 FILLER_77_1282 ();
 sg13g2_fill_1 FILLER_77_1284 ();
 sg13g2_decap_4 FILLER_77_1289 ();
 sg13g2_fill_2 FILLER_77_1293 ();
 sg13g2_decap_8 FILLER_77_1330 ();
 sg13g2_decap_8 FILLER_77_1342 ();
 sg13g2_decap_8 FILLER_77_1349 ();
 sg13g2_decap_8 FILLER_77_1356 ();
 sg13g2_decap_4 FILLER_77_1363 ();
 sg13g2_decap_4 FILLER_77_1372 ();
 sg13g2_fill_2 FILLER_77_1376 ();
 sg13g2_decap_8 FILLER_77_1388 ();
 sg13g2_decap_4 FILLER_77_1395 ();
 sg13g2_decap_8 FILLER_77_1404 ();
 sg13g2_decap_8 FILLER_77_1411 ();
 sg13g2_fill_2 FILLER_77_1444 ();
 sg13g2_fill_1 FILLER_77_1446 ();
 sg13g2_decap_8 FILLER_77_1468 ();
 sg13g2_decap_8 FILLER_77_1475 ();
 sg13g2_decap_8 FILLER_77_1482 ();
 sg13g2_fill_1 FILLER_77_1489 ();
 sg13g2_decap_8 FILLER_77_1500 ();
 sg13g2_decap_8 FILLER_77_1507 ();
 sg13g2_decap_4 FILLER_77_1514 ();
 sg13g2_decap_8 FILLER_77_1522 ();
 sg13g2_decap_8 FILLER_77_1529 ();
 sg13g2_decap_4 FILLER_77_1536 ();
 sg13g2_decap_8 FILLER_77_1544 ();
 sg13g2_decap_8 FILLER_77_1551 ();
 sg13g2_decap_8 FILLER_77_1558 ();
 sg13g2_decap_8 FILLER_77_1565 ();
 sg13g2_fill_2 FILLER_77_1572 ();
 sg13g2_decap_8 FILLER_77_1600 ();
 sg13g2_fill_1 FILLER_77_1607 ();
 sg13g2_decap_8 FILLER_77_1612 ();
 sg13g2_decap_4 FILLER_77_1619 ();
 sg13g2_fill_2 FILLER_77_1623 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_4 FILLER_78_175 ();
 sg13g2_fill_1 FILLER_78_179 ();
 sg13g2_fill_2 FILLER_78_188 ();
 sg13g2_decap_4 FILLER_78_216 ();
 sg13g2_fill_1 FILLER_78_220 ();
 sg13g2_decap_8 FILLER_78_247 ();
 sg13g2_decap_8 FILLER_78_254 ();
 sg13g2_decap_4 FILLER_78_261 ();
 sg13g2_fill_2 FILLER_78_265 ();
 sg13g2_decap_8 FILLER_78_272 ();
 sg13g2_decap_4 FILLER_78_279 ();
 sg13g2_decap_8 FILLER_78_298 ();
 sg13g2_decap_8 FILLER_78_305 ();
 sg13g2_decap_8 FILLER_78_312 ();
 sg13g2_decap_8 FILLER_78_319 ();
 sg13g2_decap_8 FILLER_78_326 ();
 sg13g2_decap_8 FILLER_78_333 ();
 sg13g2_decap_8 FILLER_78_340 ();
 sg13g2_decap_8 FILLER_78_347 ();
 sg13g2_decap_4 FILLER_78_354 ();
 sg13g2_fill_2 FILLER_78_363 ();
 sg13g2_fill_2 FILLER_78_432 ();
 sg13g2_fill_1 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_467 ();
 sg13g2_decap_4 FILLER_78_474 ();
 sg13g2_fill_2 FILLER_78_478 ();
 sg13g2_fill_1 FILLER_78_484 ();
 sg13g2_fill_2 FILLER_78_511 ();
 sg13g2_fill_1 FILLER_78_534 ();
 sg13g2_fill_2 FILLER_78_540 ();
 sg13g2_decap_8 FILLER_78_546 ();
 sg13g2_decap_8 FILLER_78_553 ();
 sg13g2_fill_2 FILLER_78_560 ();
 sg13g2_fill_1 FILLER_78_562 ();
 sg13g2_decap_8 FILLER_78_598 ();
 sg13g2_decap_8 FILLER_78_605 ();
 sg13g2_decap_8 FILLER_78_612 ();
 sg13g2_decap_8 FILLER_78_619 ();
 sg13g2_decap_4 FILLER_78_631 ();
 sg13g2_fill_1 FILLER_78_639 ();
 sg13g2_decap_4 FILLER_78_651 ();
 sg13g2_fill_1 FILLER_78_655 ();
 sg13g2_fill_1 FILLER_78_662 ();
 sg13g2_decap_8 FILLER_78_669 ();
 sg13g2_fill_1 FILLER_78_680 ();
 sg13g2_fill_2 FILLER_78_686 ();
 sg13g2_fill_1 FILLER_78_694 ();
 sg13g2_fill_1 FILLER_78_700 ();
 sg13g2_fill_1 FILLER_78_707 ();
 sg13g2_fill_1 FILLER_78_713 ();
 sg13g2_decap_8 FILLER_78_719 ();
 sg13g2_fill_1 FILLER_78_726 ();
 sg13g2_decap_8 FILLER_78_746 ();
 sg13g2_decap_8 FILLER_78_753 ();
 sg13g2_decap_8 FILLER_78_760 ();
 sg13g2_decap_8 FILLER_78_767 ();
 sg13g2_decap_8 FILLER_78_774 ();
 sg13g2_decap_8 FILLER_78_781 ();
 sg13g2_fill_2 FILLER_78_788 ();
 sg13g2_decap_8 FILLER_78_799 ();
 sg13g2_decap_8 FILLER_78_806 ();
 sg13g2_decap_8 FILLER_78_813 ();
 sg13g2_decap_4 FILLER_78_820 ();
 sg13g2_fill_2 FILLER_78_824 ();
 sg13g2_decap_8 FILLER_78_830 ();
 sg13g2_decap_4 FILLER_78_837 ();
 sg13g2_fill_2 FILLER_78_841 ();
 sg13g2_decap_8 FILLER_78_848 ();
 sg13g2_fill_1 FILLER_78_855 ();
 sg13g2_decap_4 FILLER_78_860 ();
 sg13g2_fill_1 FILLER_78_868 ();
 sg13g2_fill_2 FILLER_78_875 ();
 sg13g2_decap_4 FILLER_78_882 ();
 sg13g2_fill_2 FILLER_78_886 ();
 sg13g2_fill_1 FILLER_78_929 ();
 sg13g2_fill_1 FILLER_78_945 ();
 sg13g2_decap_4 FILLER_78_951 ();
 sg13g2_fill_2 FILLER_78_955 ();
 sg13g2_fill_1 FILLER_78_961 ();
 sg13g2_fill_1 FILLER_78_982 ();
 sg13g2_decap_4 FILLER_78_991 ();
 sg13g2_fill_1 FILLER_78_995 ();
 sg13g2_fill_2 FILLER_78_1013 ();
 sg13g2_fill_1 FILLER_78_1015 ();
 sg13g2_fill_2 FILLER_78_1026 ();
 sg13g2_fill_2 FILLER_78_1032 ();
 sg13g2_decap_8 FILLER_78_1039 ();
 sg13g2_decap_8 FILLER_78_1046 ();
 sg13g2_fill_1 FILLER_78_1053 ();
 sg13g2_fill_2 FILLER_78_1058 ();
 sg13g2_fill_1 FILLER_78_1081 ();
 sg13g2_decap_8 FILLER_78_1139 ();
 sg13g2_decap_4 FILLER_78_1146 ();
 sg13g2_fill_1 FILLER_78_1150 ();
 sg13g2_fill_2 FILLER_78_1163 ();
 sg13g2_fill_1 FILLER_78_1165 ();
 sg13g2_decap_8 FILLER_78_1176 ();
 sg13g2_decap_4 FILLER_78_1183 ();
 sg13g2_fill_1 FILLER_78_1203 ();
 sg13g2_decap_8 FILLER_78_1217 ();
 sg13g2_decap_4 FILLER_78_1224 ();
 sg13g2_fill_2 FILLER_78_1228 ();
 sg13g2_fill_2 FILLER_78_1242 ();
 sg13g2_decap_8 FILLER_78_1256 ();
 sg13g2_decap_8 FILLER_78_1263 ();
 sg13g2_decap_8 FILLER_78_1296 ();
 sg13g2_decap_4 FILLER_78_1303 ();
 sg13g2_fill_2 FILLER_78_1307 ();
 sg13g2_decap_8 FILLER_78_1313 ();
 sg13g2_fill_1 FILLER_78_1320 ();
 sg13g2_decap_8 FILLER_78_1325 ();
 sg13g2_fill_2 FILLER_78_1332 ();
 sg13g2_fill_1 FILLER_78_1334 ();
 sg13g2_decap_8 FILLER_78_1339 ();
 sg13g2_decap_8 FILLER_78_1346 ();
 sg13g2_decap_4 FILLER_78_1353 ();
 sg13g2_fill_1 FILLER_78_1357 ();
 sg13g2_decap_8 FILLER_78_1367 ();
 sg13g2_fill_2 FILLER_78_1374 ();
 sg13g2_fill_2 FILLER_78_1381 ();
 sg13g2_decap_8 FILLER_78_1416 ();
 sg13g2_decap_8 FILLER_78_1428 ();
 sg13g2_decap_8 FILLER_78_1435 ();
 sg13g2_decap_8 FILLER_78_1442 ();
 sg13g2_decap_8 FILLER_78_1449 ();
 sg13g2_decap_8 FILLER_78_1466 ();
 sg13g2_decap_8 FILLER_78_1473 ();
 sg13g2_decap_4 FILLER_78_1480 ();
 sg13g2_fill_1 FILLER_78_1484 ();
 sg13g2_fill_2 FILLER_78_1490 ();
 sg13g2_fill_1 FILLER_78_1492 ();
 sg13g2_decap_8 FILLER_78_1501 ();
 sg13g2_decap_8 FILLER_78_1508 ();
 sg13g2_decap_4 FILLER_78_1528 ();
 sg13g2_fill_1 FILLER_78_1532 ();
 sg13g2_decap_4 FILLER_78_1569 ();
 sg13g2_decap_8 FILLER_78_1582 ();
 sg13g2_fill_1 FILLER_78_1589 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_4 FILLER_79_147 ();
 sg13g2_fill_1 FILLER_79_151 ();
 sg13g2_decap_8 FILLER_79_156 ();
 sg13g2_fill_2 FILLER_79_163 ();
 sg13g2_decap_4 FILLER_79_170 ();
 sg13g2_fill_2 FILLER_79_225 ();
 sg13g2_fill_1 FILLER_79_227 ();
 sg13g2_fill_1 FILLER_79_232 ();
 sg13g2_decap_4 FILLER_79_273 ();
 sg13g2_fill_2 FILLER_79_277 ();
 sg13g2_decap_8 FILLER_79_325 ();
 sg13g2_decap_8 FILLER_79_332 ();
 sg13g2_decap_4 FILLER_79_354 ();
 sg13g2_fill_1 FILLER_79_358 ();
 sg13g2_fill_1 FILLER_79_364 ();
 sg13g2_fill_2 FILLER_79_369 ();
 sg13g2_fill_1 FILLER_79_426 ();
 sg13g2_decap_4 FILLER_79_488 ();
 sg13g2_decap_8 FILLER_79_496 ();
 sg13g2_decap_8 FILLER_79_503 ();
 sg13g2_fill_1 FILLER_79_510 ();
 sg13g2_decap_8 FILLER_79_515 ();
 sg13g2_fill_1 FILLER_79_522 ();
 sg13g2_decap_4 FILLER_79_527 ();
 sg13g2_fill_2 FILLER_79_531 ();
 sg13g2_decap_4 FILLER_79_564 ();
 sg13g2_decap_8 FILLER_79_576 ();
 sg13g2_decap_4 FILLER_79_583 ();
 sg13g2_fill_1 FILLER_79_587 ();
 sg13g2_decap_8 FILLER_79_619 ();
 sg13g2_fill_2 FILLER_79_626 ();
 sg13g2_fill_1 FILLER_79_628 ();
 sg13g2_decap_8 FILLER_79_646 ();
 sg13g2_fill_1 FILLER_79_653 ();
 sg13g2_fill_1 FILLER_79_660 ();
 sg13g2_fill_2 FILLER_79_667 ();
 sg13g2_fill_1 FILLER_79_669 ();
 sg13g2_fill_2 FILLER_79_676 ();
 sg13g2_fill_1 FILLER_79_678 ();
 sg13g2_decap_4 FILLER_79_692 ();
 sg13g2_fill_2 FILLER_79_696 ();
 sg13g2_fill_2 FILLER_79_724 ();
 sg13g2_decap_8 FILLER_79_744 ();
 sg13g2_decap_8 FILLER_79_751 ();
 sg13g2_decap_4 FILLER_79_758 ();
 sg13g2_fill_1 FILLER_79_762 ();
 sg13g2_fill_2 FILLER_79_774 ();
 sg13g2_fill_1 FILLER_79_788 ();
 sg13g2_fill_2 FILLER_79_815 ();
 sg13g2_fill_2 FILLER_79_821 ();
 sg13g2_decap_4 FILLER_79_831 ();
 sg13g2_fill_1 FILLER_79_835 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_4 FILLER_79_848 ();
 sg13g2_fill_2 FILLER_79_852 ();
 sg13g2_decap_8 FILLER_79_865 ();
 sg13g2_decap_8 FILLER_79_872 ();
 sg13g2_decap_8 FILLER_79_879 ();
 sg13g2_decap_8 FILLER_79_886 ();
 sg13g2_decap_8 FILLER_79_893 ();
 sg13g2_fill_2 FILLER_79_905 ();
 sg13g2_fill_1 FILLER_79_907 ();
 sg13g2_fill_2 FILLER_79_912 ();
 sg13g2_fill_2 FILLER_79_919 ();
 sg13g2_fill_1 FILLER_79_921 ();
 sg13g2_fill_1 FILLER_79_926 ();
 sg13g2_fill_2 FILLER_79_935 ();
 sg13g2_fill_1 FILLER_79_937 ();
 sg13g2_decap_8 FILLER_79_943 ();
 sg13g2_decap_8 FILLER_79_950 ();
 sg13g2_decap_8 FILLER_79_957 ();
 sg13g2_decap_8 FILLER_79_964 ();
 sg13g2_decap_8 FILLER_79_971 ();
 sg13g2_decap_8 FILLER_79_978 ();
 sg13g2_decap_8 FILLER_79_985 ();
 sg13g2_fill_2 FILLER_79_992 ();
 sg13g2_fill_2 FILLER_79_1020 ();
 sg13g2_fill_1 FILLER_79_1022 ();
 sg13g2_decap_8 FILLER_79_1028 ();
 sg13g2_decap_8 FILLER_79_1035 ();
 sg13g2_decap_4 FILLER_79_1042 ();
 sg13g2_fill_1 FILLER_79_1046 ();
 sg13g2_decap_4 FILLER_79_1055 ();
 sg13g2_fill_1 FILLER_79_1059 ();
 sg13g2_fill_1 FILLER_79_1070 ();
 sg13g2_fill_2 FILLER_79_1079 ();
 sg13g2_fill_1 FILLER_79_1081 ();
 sg13g2_fill_1 FILLER_79_1100 ();
 sg13g2_decap_8 FILLER_79_1145 ();
 sg13g2_fill_1 FILLER_79_1152 ();
 sg13g2_decap_8 FILLER_79_1164 ();
 sg13g2_decap_8 FILLER_79_1171 ();
 sg13g2_decap_8 FILLER_79_1178 ();
 sg13g2_decap_4 FILLER_79_1185 ();
 sg13g2_decap_8 FILLER_79_1203 ();
 sg13g2_fill_2 FILLER_79_1210 ();
 sg13g2_decap_8 FILLER_79_1220 ();
 sg13g2_fill_2 FILLER_79_1227 ();
 sg13g2_fill_1 FILLER_79_1229 ();
 sg13g2_decap_8 FILLER_79_1235 ();
 sg13g2_decap_8 FILLER_79_1242 ();
 sg13g2_decap_8 FILLER_79_1249 ();
 sg13g2_fill_2 FILLER_79_1256 ();
 sg13g2_fill_2 FILLER_79_1263 ();
 sg13g2_fill_1 FILLER_79_1265 ();
 sg13g2_decap_4 FILLER_79_1299 ();
 sg13g2_fill_1 FILLER_79_1334 ();
 sg13g2_decap_4 FILLER_79_1344 ();
 sg13g2_fill_1 FILLER_79_1348 ();
 sg13g2_decap_8 FILLER_79_1431 ();
 sg13g2_fill_1 FILLER_79_1438 ();
 sg13g2_decap_8 FILLER_79_1448 ();
 sg13g2_decap_8 FILLER_79_1472 ();
 sg13g2_decap_8 FILLER_79_1479 ();
 sg13g2_fill_1 FILLER_79_1486 ();
 sg13g2_fill_2 FILLER_79_1513 ();
 sg13g2_decap_4 FILLER_79_1541 ();
 sg13g2_fill_1 FILLER_79_1545 ();
 sg13g2_decap_8 FILLER_79_1555 ();
 sg13g2_decap_4 FILLER_79_1562 ();
 sg13g2_fill_2 FILLER_79_1591 ();
 sg13g2_fill_1 FILLER_79_1593 ();
 sg13g2_fill_1 FILLER_79_1599 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_77 ();
 sg13g2_decap_8 FILLER_80_84 ();
 sg13g2_decap_8 FILLER_80_91 ();
 sg13g2_decap_8 FILLER_80_98 ();
 sg13g2_decap_8 FILLER_80_105 ();
 sg13g2_decap_8 FILLER_80_112 ();
 sg13g2_decap_8 FILLER_80_119 ();
 sg13g2_decap_8 FILLER_80_126 ();
 sg13g2_decap_8 FILLER_80_133 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_decap_8 FILLER_80_221 ();
 sg13g2_decap_4 FILLER_80_228 ();
 sg13g2_fill_2 FILLER_80_232 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_254 ();
 sg13g2_decap_8 FILLER_80_261 ();
 sg13g2_fill_2 FILLER_80_268 ();
 sg13g2_fill_1 FILLER_80_270 ();
 sg13g2_decap_4 FILLER_80_322 ();
 sg13g2_fill_2 FILLER_80_326 ();
 sg13g2_decap_8 FILLER_80_349 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_decap_8 FILLER_80_415 ();
 sg13g2_decap_8 FILLER_80_422 ();
 sg13g2_fill_2 FILLER_80_429 ();
 sg13g2_fill_2 FILLER_80_457 ();
 sg13g2_decap_8 FILLER_80_480 ();
 sg13g2_decap_8 FILLER_80_491 ();
 sg13g2_fill_1 FILLER_80_498 ();
 sg13g2_decap_8 FILLER_80_503 ();
 sg13g2_decap_8 FILLER_80_541 ();
 sg13g2_decap_8 FILLER_80_548 ();
 sg13g2_decap_8 FILLER_80_555 ();
 sg13g2_decap_8 FILLER_80_562 ();
 sg13g2_decap_8 FILLER_80_569 ();
 sg13g2_decap_8 FILLER_80_576 ();
 sg13g2_decap_8 FILLER_80_583 ();
 sg13g2_decap_8 FILLER_80_590 ();
 sg13g2_decap_8 FILLER_80_597 ();
 sg13g2_decap_8 FILLER_80_604 ();
 sg13g2_decap_4 FILLER_80_611 ();
 sg13g2_decap_4 FILLER_80_631 ();
 sg13g2_fill_2 FILLER_80_635 ();
 sg13g2_fill_2 FILLER_80_642 ();
 sg13g2_fill_1 FILLER_80_644 ();
 sg13g2_decap_8 FILLER_80_661 ();
 sg13g2_decap_8 FILLER_80_668 ();
 sg13g2_fill_2 FILLER_80_675 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_4 FILLER_80_704 ();
 sg13g2_fill_2 FILLER_80_708 ();
 sg13g2_fill_1 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_724 ();
 sg13g2_fill_2 FILLER_80_731 ();
 sg13g2_fill_1 FILLER_80_733 ();
 sg13g2_fill_2 FILLER_80_738 ();
 sg13g2_decap_4 FILLER_80_750 ();
 sg13g2_fill_1 FILLER_80_754 ();
 sg13g2_decap_4 FILLER_80_767 ();
 sg13g2_fill_1 FILLER_80_771 ();
 sg13g2_fill_1 FILLER_80_790 ();
 sg13g2_decap_4 FILLER_80_814 ();
 sg13g2_fill_1 FILLER_80_818 ();
 sg13g2_decap_4 FILLER_80_838 ();
 sg13g2_decap_4 FILLER_80_847 ();
 sg13g2_fill_2 FILLER_80_851 ();
 sg13g2_decap_4 FILLER_80_863 ();
 sg13g2_fill_1 FILLER_80_867 ();
 sg13g2_decap_8 FILLER_80_873 ();
 sg13g2_fill_2 FILLER_80_880 ();
 sg13g2_decap_8 FILLER_80_902 ();
 sg13g2_decap_8 FILLER_80_909 ();
 sg13g2_fill_2 FILLER_80_916 ();
 sg13g2_fill_1 FILLER_80_918 ();
 sg13g2_decap_8 FILLER_80_924 ();
 sg13g2_fill_2 FILLER_80_931 ();
 sg13g2_decap_8 FILLER_80_942 ();
 sg13g2_decap_8 FILLER_80_949 ();
 sg13g2_decap_8 FILLER_80_956 ();
 sg13g2_decap_8 FILLER_80_963 ();
 sg13g2_decap_4 FILLER_80_970 ();
 sg13g2_decap_8 FILLER_80_986 ();
 sg13g2_decap_8 FILLER_80_993 ();
 sg13g2_fill_1 FILLER_80_1000 ();
 sg13g2_decap_8 FILLER_80_1005 ();
 sg13g2_fill_2 FILLER_80_1012 ();
 sg13g2_decap_8 FILLER_80_1026 ();
 sg13g2_decap_8 FILLER_80_1041 ();
 sg13g2_decap_8 FILLER_80_1048 ();
 sg13g2_decap_4 FILLER_80_1055 ();
 sg13g2_fill_2 FILLER_80_1059 ();
 sg13g2_decap_8 FILLER_80_1066 ();
 sg13g2_fill_2 FILLER_80_1114 ();
 sg13g2_decap_8 FILLER_80_1138 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_fill_2 FILLER_80_1158 ();
 sg13g2_decap_4 FILLER_80_1165 ();
 sg13g2_fill_1 FILLER_80_1169 ();
 sg13g2_decap_8 FILLER_80_1175 ();
 sg13g2_fill_2 FILLER_80_1182 ();
 sg13g2_fill_1 FILLER_80_1184 ();
 sg13g2_decap_4 FILLER_80_1189 ();
 sg13g2_fill_2 FILLER_80_1193 ();
 sg13g2_fill_2 FILLER_80_1229 ();
 sg13g2_decap_4 FILLER_80_1354 ();
 sg13g2_fill_2 FILLER_80_1358 ();
 sg13g2_decap_8 FILLER_80_1364 ();
 sg13g2_decap_8 FILLER_80_1371 ();
 sg13g2_fill_1 FILLER_80_1378 ();
 sg13g2_decap_8 FILLER_80_1383 ();
 sg13g2_fill_2 FILLER_80_1403 ();
 sg13g2_decap_4 FILLER_80_1486 ();
 sg13g2_decap_8 FILLER_80_1494 ();
 sg13g2_decap_4 FILLER_80_1501 ();
 sg13g2_fill_2 FILLER_80_1505 ();
 sg13g2_decap_8 FILLER_81_0 ();
 sg13g2_decap_8 FILLER_81_7 ();
 sg13g2_decap_8 FILLER_81_14 ();
 sg13g2_decap_8 FILLER_81_21 ();
 sg13g2_decap_8 FILLER_81_28 ();
 sg13g2_decap_8 FILLER_81_35 ();
 sg13g2_decap_8 FILLER_81_42 ();
 sg13g2_decap_8 FILLER_81_49 ();
 sg13g2_decap_8 FILLER_81_56 ();
 sg13g2_decap_8 FILLER_81_63 ();
 sg13g2_decap_8 FILLER_81_70 ();
 sg13g2_decap_8 FILLER_81_77 ();
 sg13g2_decap_8 FILLER_81_84 ();
 sg13g2_decap_8 FILLER_81_91 ();
 sg13g2_decap_8 FILLER_81_98 ();
 sg13g2_decap_8 FILLER_81_105 ();
 sg13g2_decap_8 FILLER_81_112 ();
 sg13g2_decap_8 FILLER_81_119 ();
 sg13g2_decap_8 FILLER_81_126 ();
 sg13g2_decap_8 FILLER_81_133 ();
 sg13g2_decap_8 FILLER_81_140 ();
 sg13g2_decap_8 FILLER_81_147 ();
 sg13g2_decap_8 FILLER_81_154 ();
 sg13g2_fill_2 FILLER_81_161 ();
 sg13g2_fill_1 FILLER_81_163 ();
 sg13g2_decap_4 FILLER_81_173 ();
 sg13g2_fill_1 FILLER_81_177 ();
 sg13g2_decap_8 FILLER_81_182 ();
 sg13g2_decap_8 FILLER_81_189 ();
 sg13g2_decap_8 FILLER_81_196 ();
 sg13g2_decap_4 FILLER_81_203 ();
 sg13g2_decap_8 FILLER_81_211 ();
 sg13g2_decap_4 FILLER_81_218 ();
 sg13g2_fill_1 FILLER_81_222 ();
 sg13g2_decap_8 FILLER_81_249 ();
 sg13g2_decap_8 FILLER_81_256 ();
 sg13g2_decap_8 FILLER_81_263 ();
 sg13g2_decap_8 FILLER_81_270 ();
 sg13g2_decap_8 FILLER_81_281 ();
 sg13g2_decap_8 FILLER_81_288 ();
 sg13g2_decap_8 FILLER_81_295 ();
 sg13g2_decap_8 FILLER_81_302 ();
 sg13g2_decap_8 FILLER_81_309 ();
 sg13g2_decap_4 FILLER_81_316 ();
 sg13g2_fill_2 FILLER_81_356 ();
 sg13g2_fill_1 FILLER_81_358 ();
 sg13g2_fill_2 FILLER_81_384 ();
 sg13g2_fill_1 FILLER_81_386 ();
 sg13g2_decap_8 FILLER_81_418 ();
 sg13g2_decap_8 FILLER_81_425 ();
 sg13g2_decap_4 FILLER_81_432 ();
 sg13g2_fill_2 FILLER_81_436 ();
 sg13g2_decap_8 FILLER_81_442 ();
 sg13g2_decap_4 FILLER_81_449 ();
 sg13g2_fill_1 FILLER_81_453 ();
 sg13g2_decap_8 FILLER_81_463 ();
 sg13g2_decap_8 FILLER_81_470 ();
 sg13g2_decap_4 FILLER_81_477 ();
 sg13g2_fill_1 FILLER_81_481 ();
 sg13g2_fill_2 FILLER_81_485 ();
 sg13g2_decap_4 FILLER_81_518 ();
 sg13g2_fill_2 FILLER_81_522 ();
 sg13g2_decap_8 FILLER_81_554 ();
 sg13g2_decap_8 FILLER_81_570 ();
 sg13g2_decap_4 FILLER_81_577 ();
 sg13g2_fill_2 FILLER_81_586 ();
 sg13g2_fill_1 FILLER_81_588 ();
 sg13g2_decap_8 FILLER_81_593 ();
 sg13g2_decap_4 FILLER_81_600 ();
 sg13g2_fill_2 FILLER_81_641 ();
 sg13g2_fill_1 FILLER_81_643 ();
 sg13g2_fill_2 FILLER_81_648 ();
 sg13g2_fill_1 FILLER_81_650 ();
 sg13g2_fill_2 FILLER_81_655 ();
 sg13g2_decap_8 FILLER_81_665 ();
 sg13g2_decap_8 FILLER_81_672 ();
 sg13g2_fill_2 FILLER_81_679 ();
 sg13g2_fill_1 FILLER_81_681 ();
 sg13g2_fill_2 FILLER_81_686 ();
 sg13g2_fill_1 FILLER_81_688 ();
 sg13g2_decap_8 FILLER_81_697 ();
 sg13g2_fill_2 FILLER_81_704 ();
 sg13g2_fill_1 FILLER_81_706 ();
 sg13g2_decap_8 FILLER_81_726 ();
 sg13g2_decap_8 FILLER_81_733 ();
 sg13g2_decap_4 FILLER_81_740 ();
 sg13g2_decap_8 FILLER_81_784 ();
 sg13g2_fill_2 FILLER_81_791 ();
 sg13g2_decap_4 FILLER_81_797 ();
 sg13g2_fill_1 FILLER_81_801 ();
 sg13g2_decap_8 FILLER_81_811 ();
 sg13g2_decap_8 FILLER_81_818 ();
 sg13g2_decap_8 FILLER_81_825 ();
 sg13g2_decap_8 FILLER_81_832 ();
 sg13g2_decap_8 FILLER_81_839 ();
 sg13g2_decap_4 FILLER_81_846 ();
 sg13g2_fill_2 FILLER_81_850 ();
 sg13g2_decap_8 FILLER_81_877 ();
 sg13g2_decap_8 FILLER_81_917 ();
 sg13g2_decap_8 FILLER_81_924 ();
 sg13g2_fill_2 FILLER_81_931 ();
 sg13g2_decap_8 FILLER_81_941 ();
 sg13g2_fill_2 FILLER_81_948 ();
 sg13g2_decap_4 FILLER_81_958 ();
 sg13g2_fill_2 FILLER_81_962 ();
 sg13g2_decap_4 FILLER_81_968 ();
 sg13g2_fill_1 FILLER_81_972 ();
 sg13g2_decap_8 FILLER_81_985 ();
 sg13g2_decap_8 FILLER_81_992 ();
 sg13g2_decap_4 FILLER_81_999 ();
 sg13g2_fill_1 FILLER_81_1003 ();
 sg13g2_decap_4 FILLER_81_1009 ();
 sg13g2_fill_2 FILLER_81_1013 ();
 sg13g2_fill_2 FILLER_81_1039 ();
 sg13g2_fill_1 FILLER_81_1050 ();
 sg13g2_fill_1 FILLER_81_1134 ();
 sg13g2_fill_1 FILLER_81_1140 ();
 sg13g2_fill_1 FILLER_81_1145 ();
 sg13g2_fill_2 FILLER_81_1151 ();
 sg13g2_decap_8 FILLER_81_1165 ();
 sg13g2_fill_1 FILLER_81_1172 ();
 sg13g2_decap_8 FILLER_81_1209 ();
 sg13g2_decap_8 FILLER_81_1248 ();
 sg13g2_decap_8 FILLER_81_1255 ();
 sg13g2_fill_2 FILLER_81_1265 ();
 sg13g2_fill_2 FILLER_81_1276 ();
 sg13g2_fill_1 FILLER_81_1278 ();
 sg13g2_decap_4 FILLER_81_1310 ();
 sg13g2_fill_2 FILLER_81_1318 ();
 sg13g2_fill_1 FILLER_81_1320 ();
 sg13g2_fill_2 FILLER_81_1384 ();
 sg13g2_fill_1 FILLER_81_1442 ();
 sg13g2_decap_8 FILLER_81_1509 ();
 sg13g2_decap_8 FILLER_81_1516 ();
 sg13g2_decap_8 FILLER_81_1523 ();
 sg13g2_decap_8 FILLER_81_1530 ();
 sg13g2_decap_8 FILLER_81_1537 ();
 sg13g2_fill_1 FILLER_81_1544 ();
 sg13g2_decap_8 FILLER_81_1571 ();
 sg13g2_decap_8 FILLER_81_1578 ();
 sg13g2_decap_8 FILLER_81_1585 ();
 sg13g2_decap_8 FILLER_81_1592 ();
 sg13g2_decap_8 FILLER_81_1599 ();
 sg13g2_fill_2 FILLER_81_1606 ();
 sg13g2_decap_8 FILLER_81_1612 ();
 sg13g2_decap_4 FILLER_81_1619 ();
 sg13g2_fill_2 FILLER_81_1623 ();
 sg13g2_decap_8 FILLER_82_0 ();
 sg13g2_decap_8 FILLER_82_7 ();
 sg13g2_decap_8 FILLER_82_14 ();
 sg13g2_decap_8 FILLER_82_21 ();
 sg13g2_decap_8 FILLER_82_28 ();
 sg13g2_decap_8 FILLER_82_35 ();
 sg13g2_decap_8 FILLER_82_42 ();
 sg13g2_decap_8 FILLER_82_49 ();
 sg13g2_decap_8 FILLER_82_56 ();
 sg13g2_decap_8 FILLER_82_63 ();
 sg13g2_decap_8 FILLER_82_70 ();
 sg13g2_decap_8 FILLER_82_77 ();
 sg13g2_decap_8 FILLER_82_84 ();
 sg13g2_decap_8 FILLER_82_91 ();
 sg13g2_decap_8 FILLER_82_98 ();
 sg13g2_decap_8 FILLER_82_105 ();
 sg13g2_decap_8 FILLER_82_112 ();
 sg13g2_decap_8 FILLER_82_119 ();
 sg13g2_decap_8 FILLER_82_126 ();
 sg13g2_decap_8 FILLER_82_133 ();
 sg13g2_fill_2 FILLER_82_140 ();
 sg13g2_fill_2 FILLER_82_178 ();
 sg13g2_fill_1 FILLER_82_184 ();
 sg13g2_decap_4 FILLER_82_194 ();
 sg13g2_fill_2 FILLER_82_198 ();
 sg13g2_decap_4 FILLER_82_221 ();
 sg13g2_fill_2 FILLER_82_225 ();
 sg13g2_decap_4 FILLER_82_234 ();
 sg13g2_fill_2 FILLER_82_247 ();
 sg13g2_decap_4 FILLER_82_270 ();
 sg13g2_fill_1 FILLER_82_274 ();
 sg13g2_decap_8 FILLER_82_296 ();
 sg13g2_fill_2 FILLER_82_303 ();
 sg13g2_decap_8 FILLER_82_315 ();
 sg13g2_decap_8 FILLER_82_322 ();
 sg13g2_decap_8 FILLER_82_329 ();
 sg13g2_fill_1 FILLER_82_336 ();
 sg13g2_decap_4 FILLER_82_342 ();
 sg13g2_fill_2 FILLER_82_346 ();
 sg13g2_fill_2 FILLER_82_388 ();
 sg13g2_fill_1 FILLER_82_390 ();
 sg13g2_fill_2 FILLER_82_420 ();
 sg13g2_fill_1 FILLER_82_422 ();
 sg13g2_decap_8 FILLER_82_444 ();
 sg13g2_decap_8 FILLER_82_451 ();
 sg13g2_decap_8 FILLER_82_526 ();
 sg13g2_decap_4 FILLER_82_533 ();
 sg13g2_fill_2 FILLER_82_537 ();
 sg13g2_fill_1 FILLER_82_543 ();
 sg13g2_fill_2 FILLER_82_553 ();
 sg13g2_fill_1 FILLER_82_555 ();
 sg13g2_fill_1 FILLER_82_647 ();
 sg13g2_decap_4 FILLER_82_653 ();
 sg13g2_decap_8 FILLER_82_665 ();
 sg13g2_fill_2 FILLER_82_672 ();
 sg13g2_decap_4 FILLER_82_700 ();
 sg13g2_fill_1 FILLER_82_732 ();
 sg13g2_fill_1 FILLER_82_741 ();
 sg13g2_decap_8 FILLER_82_746 ();
 sg13g2_fill_1 FILLER_82_753 ();
 sg13g2_decap_8 FILLER_82_758 ();
 sg13g2_decap_8 FILLER_82_765 ();
 sg13g2_decap_8 FILLER_82_772 ();
 sg13g2_decap_8 FILLER_82_779 ();
 sg13g2_decap_8 FILLER_82_786 ();
 sg13g2_decap_8 FILLER_82_793 ();
 sg13g2_decap_4 FILLER_82_800 ();
 sg13g2_fill_2 FILLER_82_804 ();
 sg13g2_decap_8 FILLER_82_811 ();
 sg13g2_fill_2 FILLER_82_818 ();
 sg13g2_fill_2 FILLER_82_836 ();
 sg13g2_fill_1 FILLER_82_838 ();
 sg13g2_fill_2 FILLER_82_844 ();
 sg13g2_fill_1 FILLER_82_846 ();
 sg13g2_fill_2 FILLER_82_855 ();
 sg13g2_fill_1 FILLER_82_861 ();
 sg13g2_decap_8 FILLER_82_867 ();
 sg13g2_decap_8 FILLER_82_874 ();
 sg13g2_decap_8 FILLER_82_881 ();
 sg13g2_decap_8 FILLER_82_888 ();
 sg13g2_fill_2 FILLER_82_895 ();
 sg13g2_fill_1 FILLER_82_897 ();
 sg13g2_decap_8 FILLER_82_902 ();
 sg13g2_fill_1 FILLER_82_909 ();
 sg13g2_decap_8 FILLER_82_918 ();
 sg13g2_decap_4 FILLER_82_925 ();
 sg13g2_fill_1 FILLER_82_929 ();
 sg13g2_fill_2 FILLER_82_933 ();
 sg13g2_fill_1 FILLER_82_935 ();
 sg13g2_fill_2 FILLER_82_943 ();
 sg13g2_fill_2 FILLER_82_950 ();
 sg13g2_fill_1 FILLER_82_970 ();
 sg13g2_decap_8 FILLER_82_976 ();
 sg13g2_decap_8 FILLER_82_983 ();
 sg13g2_decap_8 FILLER_82_990 ();
 sg13g2_decap_8 FILLER_82_997 ();
 sg13g2_decap_4 FILLER_82_1004 ();
 sg13g2_fill_1 FILLER_82_1008 ();
 sg13g2_decap_8 FILLER_82_1017 ();
 sg13g2_decap_8 FILLER_82_1034 ();
 sg13g2_decap_8 FILLER_82_1041 ();
 sg13g2_fill_2 FILLER_82_1048 ();
 sg13g2_fill_1 FILLER_82_1072 ();
 sg13g2_fill_1 FILLER_82_1110 ();
 sg13g2_fill_2 FILLER_82_1122 ();
 sg13g2_decap_8 FILLER_82_1133 ();
 sg13g2_decap_8 FILLER_82_1140 ();
 sg13g2_fill_2 FILLER_82_1166 ();
 sg13g2_fill_1 FILLER_82_1168 ();
 sg13g2_fill_1 FILLER_82_1181 ();
 sg13g2_fill_2 FILLER_82_1186 ();
 sg13g2_fill_2 FILLER_82_1196 ();
 sg13g2_decap_4 FILLER_82_1205 ();
 sg13g2_decap_8 FILLER_82_1214 ();
 sg13g2_decap_4 FILLER_82_1221 ();
 sg13g2_decap_8 FILLER_82_1251 ();
 sg13g2_decap_8 FILLER_82_1258 ();
 sg13g2_fill_1 FILLER_82_1265 ();
 sg13g2_fill_1 FILLER_82_1300 ();
 sg13g2_fill_1 FILLER_82_1336 ();
 sg13g2_decap_4 FILLER_82_1423 ();
 sg13g2_decap_8 FILLER_82_1507 ();
 sg13g2_decap_8 FILLER_82_1514 ();
 sg13g2_fill_1 FILLER_82_1521 ();
 sg13g2_decap_8 FILLER_82_1543 ();
 sg13g2_fill_2 FILLER_82_1550 ();
 sg13g2_decap_8 FILLER_82_1556 ();
 sg13g2_decap_8 FILLER_82_1563 ();
 sg13g2_decap_8 FILLER_82_1591 ();
 sg13g2_decap_4 FILLER_82_1598 ();
 sg13g2_fill_1 FILLER_82_1602 ();
 sg13g2_decap_8 FILLER_82_1611 ();
 sg13g2_decap_8 FILLER_82_1618 ();
 sg13g2_decap_8 FILLER_83_0 ();
 sg13g2_decap_8 FILLER_83_7 ();
 sg13g2_decap_8 FILLER_83_14 ();
 sg13g2_decap_8 FILLER_83_21 ();
 sg13g2_decap_8 FILLER_83_28 ();
 sg13g2_decap_8 FILLER_83_35 ();
 sg13g2_decap_8 FILLER_83_42 ();
 sg13g2_decap_8 FILLER_83_49 ();
 sg13g2_decap_8 FILLER_83_56 ();
 sg13g2_decap_8 FILLER_83_63 ();
 sg13g2_decap_8 FILLER_83_70 ();
 sg13g2_decap_8 FILLER_83_77 ();
 sg13g2_decap_8 FILLER_83_84 ();
 sg13g2_decap_8 FILLER_83_91 ();
 sg13g2_decap_8 FILLER_83_98 ();
 sg13g2_decap_8 FILLER_83_105 ();
 sg13g2_decap_8 FILLER_83_112 ();
 sg13g2_decap_8 FILLER_83_119 ();
 sg13g2_decap_8 FILLER_83_126 ();
 sg13g2_decap_8 FILLER_83_133 ();
 sg13g2_decap_4 FILLER_83_140 ();
 sg13g2_fill_1 FILLER_83_144 ();
 sg13g2_fill_1 FILLER_83_171 ();
 sg13g2_fill_2 FILLER_83_198 ();
 sg13g2_fill_2 FILLER_83_221 ();
 sg13g2_fill_2 FILLER_83_252 ();
 sg13g2_fill_1 FILLER_83_254 ();
 sg13g2_decap_8 FILLER_83_276 ();
 sg13g2_decap_8 FILLER_83_283 ();
 sg13g2_decap_4 FILLER_83_311 ();
 sg13g2_fill_2 FILLER_83_315 ();
 sg13g2_fill_2 FILLER_83_343 ();
 sg13g2_fill_1 FILLER_83_345 ();
 sg13g2_decap_8 FILLER_83_350 ();
 sg13g2_fill_2 FILLER_83_357 ();
 sg13g2_fill_1 FILLER_83_359 ();
 sg13g2_fill_1 FILLER_83_394 ();
 sg13g2_fill_1 FILLER_83_399 ();
 sg13g2_decap_4 FILLER_83_421 ();
 sg13g2_decap_8 FILLER_83_474 ();
 sg13g2_decap_8 FILLER_83_481 ();
 sg13g2_decap_8 FILLER_83_488 ();
 sg13g2_decap_8 FILLER_83_495 ();
 sg13g2_fill_2 FILLER_83_502 ();
 sg13g2_fill_2 FILLER_83_530 ();
 sg13g2_fill_1 FILLER_83_532 ();
 sg13g2_fill_2 FILLER_83_559 ();
 sg13g2_fill_1 FILLER_83_561 ();
 sg13g2_decap_4 FILLER_83_566 ();
 sg13g2_decap_8 FILLER_83_575 ();
 sg13g2_fill_2 FILLER_83_586 ();
 sg13g2_fill_2 FILLER_83_617 ();
 sg13g2_fill_2 FILLER_83_630 ();
 sg13g2_decap_4 FILLER_83_646 ();
 sg13g2_fill_1 FILLER_83_650 ();
 sg13g2_decap_8 FILLER_83_671 ();
 sg13g2_decap_8 FILLER_83_678 ();
 sg13g2_decap_8 FILLER_83_685 ();
 sg13g2_decap_8 FILLER_83_692 ();
 sg13g2_fill_2 FILLER_83_699 ();
 sg13g2_fill_1 FILLER_83_701 ();
 sg13g2_fill_2 FILLER_83_707 ();
 sg13g2_decap_8 FILLER_83_716 ();
 sg13g2_decap_8 FILLER_83_723 ();
 sg13g2_decap_8 FILLER_83_730 ();
 sg13g2_decap_8 FILLER_83_737 ();
 sg13g2_decap_8 FILLER_83_744 ();
 sg13g2_decap_8 FILLER_83_751 ();
 sg13g2_decap_8 FILLER_83_758 ();
 sg13g2_decap_8 FILLER_83_765 ();
 sg13g2_decap_4 FILLER_83_772 ();
 sg13g2_fill_2 FILLER_83_776 ();
 sg13g2_fill_2 FILLER_83_786 ();
 sg13g2_fill_2 FILLER_83_813 ();
 sg13g2_fill_1 FILLER_83_815 ();
 sg13g2_fill_1 FILLER_83_821 ();
 sg13g2_decap_4 FILLER_83_826 ();
 sg13g2_fill_1 FILLER_83_830 ();
 sg13g2_fill_2 FILLER_83_853 ();
 sg13g2_fill_1 FILLER_83_860 ();
 sg13g2_decap_8 FILLER_83_866 ();
 sg13g2_fill_2 FILLER_83_873 ();
 sg13g2_fill_2 FILLER_83_880 ();
 sg13g2_fill_1 FILLER_83_882 ();
 sg13g2_decap_8 FILLER_83_896 ();
 sg13g2_decap_8 FILLER_83_903 ();
 sg13g2_fill_2 FILLER_83_910 ();
 sg13g2_decap_4 FILLER_83_916 ();
 sg13g2_fill_1 FILLER_83_930 ();
 sg13g2_fill_2 FILLER_83_936 ();
 sg13g2_fill_1 FILLER_83_946 ();
 sg13g2_fill_2 FILLER_83_952 ();
 sg13g2_fill_2 FILLER_83_959 ();
 sg13g2_decap_8 FILLER_83_982 ();
 sg13g2_decap_8 FILLER_83_989 ();
 sg13g2_fill_2 FILLER_83_996 ();
 sg13g2_fill_1 FILLER_83_998 ();
 sg13g2_decap_4 FILLER_83_1005 ();
 sg13g2_fill_1 FILLER_83_1009 ();
 sg13g2_decap_8 FILLER_83_1025 ();
 sg13g2_decap_8 FILLER_83_1032 ();
 sg13g2_fill_2 FILLER_83_1039 ();
 sg13g2_fill_1 FILLER_83_1041 ();
 sg13g2_fill_1 FILLER_83_1055 ();
 sg13g2_fill_1 FILLER_83_1061 ();
 sg13g2_decap_8 FILLER_83_1066 ();
 sg13g2_decap_8 FILLER_83_1073 ();
 sg13g2_decap_4 FILLER_83_1080 ();
 sg13g2_fill_2 FILLER_83_1084 ();
 sg13g2_decap_4 FILLER_83_1091 ();
 sg13g2_fill_1 FILLER_83_1112 ();
 sg13g2_fill_2 FILLER_83_1131 ();
 sg13g2_decap_4 FILLER_83_1144 ();
 sg13g2_fill_2 FILLER_83_1148 ();
 sg13g2_decap_8 FILLER_83_1155 ();
 sg13g2_decap_8 FILLER_83_1162 ();
 sg13g2_decap_8 FILLER_83_1169 ();
 sg13g2_decap_4 FILLER_83_1176 ();
 sg13g2_fill_1 FILLER_83_1180 ();
 sg13g2_decap_8 FILLER_83_1191 ();
 sg13g2_fill_1 FILLER_83_1198 ();
 sg13g2_fill_2 FILLER_83_1209 ();
 sg13g2_decap_8 FILLER_83_1241 ();
 sg13g2_decap_8 FILLER_83_1248 ();
 sg13g2_decap_8 FILLER_83_1255 ();
 sg13g2_fill_2 FILLER_83_1262 ();
 sg13g2_fill_1 FILLER_83_1264 ();
 sg13g2_decap_4 FILLER_83_1345 ();
 sg13g2_fill_1 FILLER_83_1349 ();
 sg13g2_decap_8 FILLER_83_1383 ();
 sg13g2_decap_8 FILLER_83_1390 ();
 sg13g2_fill_2 FILLER_83_1397 ();
 sg13g2_fill_1 FILLER_83_1399 ();
 sg13g2_decap_8 FILLER_83_1404 ();
 sg13g2_decap_8 FILLER_83_1411 ();
 sg13g2_fill_1 FILLER_83_1418 ();
 sg13g2_fill_2 FILLER_83_1440 ();
 sg13g2_fill_1 FILLER_83_1442 ();
 sg13g2_decap_8 FILLER_83_1477 ();
 sg13g2_fill_1 FILLER_83_1484 ();
 sg13g2_decap_8 FILLER_83_1536 ();
 sg13g2_fill_2 FILLER_83_1543 ();
 sg13g2_fill_1 FILLER_83_1545 ();
 sg13g2_decap_4 FILLER_83_1563 ();
 sg13g2_fill_2 FILLER_83_1567 ();
 sg13g2_decap_8 FILLER_84_0 ();
 sg13g2_decap_8 FILLER_84_7 ();
 sg13g2_decap_8 FILLER_84_14 ();
 sg13g2_decap_8 FILLER_84_21 ();
 sg13g2_decap_8 FILLER_84_28 ();
 sg13g2_decap_8 FILLER_84_35 ();
 sg13g2_decap_8 FILLER_84_42 ();
 sg13g2_decap_8 FILLER_84_49 ();
 sg13g2_decap_8 FILLER_84_56 ();
 sg13g2_decap_8 FILLER_84_63 ();
 sg13g2_decap_8 FILLER_84_70 ();
 sg13g2_decap_8 FILLER_84_77 ();
 sg13g2_decap_8 FILLER_84_84 ();
 sg13g2_decap_8 FILLER_84_91 ();
 sg13g2_decap_8 FILLER_84_98 ();
 sg13g2_decap_8 FILLER_84_105 ();
 sg13g2_decap_8 FILLER_84_112 ();
 sg13g2_decap_8 FILLER_84_119 ();
 sg13g2_decap_8 FILLER_84_126 ();
 sg13g2_decap_8 FILLER_84_133 ();
 sg13g2_decap_8 FILLER_84_140 ();
 sg13g2_decap_8 FILLER_84_147 ();
 sg13g2_decap_4 FILLER_84_154 ();
 sg13g2_fill_1 FILLER_84_158 ();
 sg13g2_decap_8 FILLER_84_253 ();
 sg13g2_decap_8 FILLER_84_260 ();
 sg13g2_decap_8 FILLER_84_267 ();
 sg13g2_fill_2 FILLER_84_274 ();
 sg13g2_decap_8 FILLER_84_297 ();
 sg13g2_decap_8 FILLER_84_304 ();
 sg13g2_decap_4 FILLER_84_311 ();
 sg13g2_fill_2 FILLER_84_315 ();
 sg13g2_fill_2 FILLER_84_364 ();
 sg13g2_fill_1 FILLER_84_366 ();
 sg13g2_decap_8 FILLER_84_417 ();
 sg13g2_decap_8 FILLER_84_424 ();
 sg13g2_decap_8 FILLER_84_431 ();
 sg13g2_decap_8 FILLER_84_438 ();
 sg13g2_decap_8 FILLER_84_445 ();
 sg13g2_decap_4 FILLER_84_452 ();
 sg13g2_fill_2 FILLER_84_456 ();
 sg13g2_fill_2 FILLER_84_488 ();
 sg13g2_fill_1 FILLER_84_490 ();
 sg13g2_decap_8 FILLER_84_495 ();
 sg13g2_decap_8 FILLER_84_502 ();
 sg13g2_decap_8 FILLER_84_509 ();
 sg13g2_fill_2 FILLER_84_516 ();
 sg13g2_fill_1 FILLER_84_518 ();
 sg13g2_fill_1 FILLER_84_548 ();
 sg13g2_fill_2 FILLER_84_553 ();
 sg13g2_fill_2 FILLER_84_559 ();
 sg13g2_decap_8 FILLER_84_571 ();
 sg13g2_decap_8 FILLER_84_578 ();
 sg13g2_decap_8 FILLER_84_585 ();
 sg13g2_fill_1 FILLER_84_623 ();
 sg13g2_decap_8 FILLER_84_642 ();
 sg13g2_decap_8 FILLER_84_649 ();
 sg13g2_decap_8 FILLER_84_656 ();
 sg13g2_decap_8 FILLER_84_663 ();
 sg13g2_decap_8 FILLER_84_670 ();
 sg13g2_fill_2 FILLER_84_677 ();
 sg13g2_decap_8 FILLER_84_695 ();
 sg13g2_decap_4 FILLER_84_702 ();
 sg13g2_decap_4 FILLER_84_714 ();
 sg13g2_fill_2 FILLER_84_718 ();
 sg13g2_decap_4 FILLER_84_730 ();
 sg13g2_decap_4 FILLER_84_742 ();
 sg13g2_fill_1 FILLER_84_746 ();
 sg13g2_fill_2 FILLER_84_756 ();
 sg13g2_decap_4 FILLER_84_773 ();
 sg13g2_fill_2 FILLER_84_777 ();
 sg13g2_fill_1 FILLER_84_783 ();
 sg13g2_decap_8 FILLER_84_794 ();
 sg13g2_decap_8 FILLER_84_801 ();
 sg13g2_decap_8 FILLER_84_808 ();
 sg13g2_decap_8 FILLER_84_815 ();
 sg13g2_decap_8 FILLER_84_822 ();
 sg13g2_decap_8 FILLER_84_837 ();
 sg13g2_decap_8 FILLER_84_844 ();
 sg13g2_fill_2 FILLER_84_851 ();
 sg13g2_fill_1 FILLER_84_853 ();
 sg13g2_decap_4 FILLER_84_862 ();
 sg13g2_fill_1 FILLER_84_866 ();
 sg13g2_decap_4 FILLER_84_883 ();
 sg13g2_fill_2 FILLER_84_892 ();
 sg13g2_decap_8 FILLER_84_899 ();
 sg13g2_fill_1 FILLER_84_906 ();
 sg13g2_fill_1 FILLER_84_911 ();
 sg13g2_decap_8 FILLER_84_930 ();
 sg13g2_decap_8 FILLER_84_937 ();
 sg13g2_fill_2 FILLER_84_944 ();
 sg13g2_fill_1 FILLER_84_946 ();
 sg13g2_fill_1 FILLER_84_953 ();
 sg13g2_fill_1 FILLER_84_958 ();
 sg13g2_fill_1 FILLER_84_969 ();
 sg13g2_fill_2 FILLER_84_978 ();
 sg13g2_fill_1 FILLER_84_1002 ();
 sg13g2_fill_1 FILLER_84_1008 ();
 sg13g2_fill_1 FILLER_84_1018 ();
 sg13g2_fill_1 FILLER_84_1029 ();
 sg13g2_fill_1 FILLER_84_1042 ();
 sg13g2_fill_1 FILLER_84_1049 ();
 sg13g2_fill_1 FILLER_84_1060 ();
 sg13g2_fill_2 FILLER_84_1074 ();
 sg13g2_fill_1 FILLER_84_1076 ();
 sg13g2_decap_4 FILLER_84_1098 ();
 sg13g2_decap_8 FILLER_84_1107 ();
 sg13g2_fill_2 FILLER_84_1114 ();
 sg13g2_fill_2 FILLER_84_1121 ();
 sg13g2_decap_4 FILLER_84_1126 ();
 sg13g2_fill_2 FILLER_84_1130 ();
 sg13g2_fill_2 FILLER_84_1148 ();
 sg13g2_fill_1 FILLER_84_1168 ();
 sg13g2_decap_8 FILLER_84_1177 ();
 sg13g2_decap_8 FILLER_84_1199 ();
 sg13g2_decap_8 FILLER_84_1206 ();
 sg13g2_decap_4 FILLER_84_1213 ();
 sg13g2_fill_2 FILLER_84_1227 ();
 sg13g2_fill_1 FILLER_84_1229 ();
 sg13g2_fill_1 FILLER_84_1256 ();
 sg13g2_decap_8 FILLER_84_1313 ();
 sg13g2_decap_4 FILLER_84_1341 ();
 sg13g2_fill_2 FILLER_84_1345 ();
 sg13g2_fill_2 FILLER_84_1352 ();
 sg13g2_decap_8 FILLER_84_1368 ();
 sg13g2_decap_8 FILLER_84_1375 ();
 sg13g2_decap_8 FILLER_84_1382 ();
 sg13g2_decap_4 FILLER_84_1389 ();
 sg13g2_fill_2 FILLER_84_1393 ();
 sg13g2_fill_2 FILLER_84_1404 ();
 sg13g2_decap_8 FILLER_84_1410 ();
 sg13g2_decap_4 FILLER_84_1417 ();
 sg13g2_fill_1 FILLER_84_1421 ();
 sg13g2_decap_4 FILLER_84_1493 ();
 sg13g2_fill_1 FILLER_84_1497 ();
 sg13g2_decap_4 FILLER_84_1536 ();
 sg13g2_decap_8 FILLER_84_1569 ();
 sg13g2_decap_8 FILLER_84_1576 ();
 sg13g2_decap_8 FILLER_84_1583 ();
 sg13g2_fill_1 FILLER_84_1590 ();
 sg13g2_decap_8 FILLER_85_0 ();
 sg13g2_decap_8 FILLER_85_7 ();
 sg13g2_decap_8 FILLER_85_14 ();
 sg13g2_decap_8 FILLER_85_21 ();
 sg13g2_decap_8 FILLER_85_28 ();
 sg13g2_decap_8 FILLER_85_35 ();
 sg13g2_decap_8 FILLER_85_42 ();
 sg13g2_decap_8 FILLER_85_49 ();
 sg13g2_decap_8 FILLER_85_56 ();
 sg13g2_decap_8 FILLER_85_63 ();
 sg13g2_decap_8 FILLER_85_70 ();
 sg13g2_decap_8 FILLER_85_77 ();
 sg13g2_decap_8 FILLER_85_84 ();
 sg13g2_decap_8 FILLER_85_91 ();
 sg13g2_decap_8 FILLER_85_98 ();
 sg13g2_decap_8 FILLER_85_105 ();
 sg13g2_decap_8 FILLER_85_112 ();
 sg13g2_decap_8 FILLER_85_119 ();
 sg13g2_decap_8 FILLER_85_126 ();
 sg13g2_decap_8 FILLER_85_133 ();
 sg13g2_decap_8 FILLER_85_140 ();
 sg13g2_decap_8 FILLER_85_147 ();
 sg13g2_fill_2 FILLER_85_154 ();
 sg13g2_fill_2 FILLER_85_220 ();
 sg13g2_decap_4 FILLER_85_260 ();
 sg13g2_fill_1 FILLER_85_264 ();
 sg13g2_fill_2 FILLER_85_269 ();
 sg13g2_fill_1 FILLER_85_271 ();
 sg13g2_fill_2 FILLER_85_293 ();
 sg13g2_decap_8 FILLER_85_299 ();
 sg13g2_decap_8 FILLER_85_306 ();
 sg13g2_fill_1 FILLER_85_313 ();
 sg13g2_decap_8 FILLER_85_319 ();
 sg13g2_decap_8 FILLER_85_326 ();
 sg13g2_decap_4 FILLER_85_333 ();
 sg13g2_fill_2 FILLER_85_337 ();
 sg13g2_decap_8 FILLER_85_343 ();
 sg13g2_fill_2 FILLER_85_350 ();
 sg13g2_fill_1 FILLER_85_352 ();
 sg13g2_decap_8 FILLER_85_419 ();
 sg13g2_decap_8 FILLER_85_430 ();
 sg13g2_fill_1 FILLER_85_437 ();
 sg13g2_decap_8 FILLER_85_447 ();
 sg13g2_fill_2 FILLER_85_454 ();
 sg13g2_decap_4 FILLER_85_509 ();
 sg13g2_fill_2 FILLER_85_513 ();
 sg13g2_decap_4 FILLER_85_546 ();
 sg13g2_fill_1 FILLER_85_550 ();
 sg13g2_decap_8 FILLER_85_556 ();
 sg13g2_decap_8 FILLER_85_563 ();
 sg13g2_decap_4 FILLER_85_574 ();
 sg13g2_fill_2 FILLER_85_578 ();
 sg13g2_decap_8 FILLER_85_584 ();
 sg13g2_decap_8 FILLER_85_591 ();
 sg13g2_decap_8 FILLER_85_598 ();
 sg13g2_decap_4 FILLER_85_605 ();
 sg13g2_fill_1 FILLER_85_609 ();
 sg13g2_decap_8 FILLER_85_619 ();
 sg13g2_decap_8 FILLER_85_626 ();
 sg13g2_decap_8 FILLER_85_633 ();
 sg13g2_decap_4 FILLER_85_640 ();
 sg13g2_decap_8 FILLER_85_648 ();
 sg13g2_decap_4 FILLER_85_655 ();
 sg13g2_decap_4 FILLER_85_673 ();
 sg13g2_fill_1 FILLER_85_677 ();
 sg13g2_decap_8 FILLER_85_682 ();
 sg13g2_decap_4 FILLER_85_689 ();
 sg13g2_fill_1 FILLER_85_693 ();
 sg13g2_decap_4 FILLER_85_730 ();
 sg13g2_fill_1 FILLER_85_734 ();
 sg13g2_decap_4 FILLER_85_740 ();
 sg13g2_fill_1 FILLER_85_762 ();
 sg13g2_fill_2 FILLER_85_767 ();
 sg13g2_fill_2 FILLER_85_777 ();
 sg13g2_fill_1 FILLER_85_779 ();
 sg13g2_decap_8 FILLER_85_793 ();
 sg13g2_fill_2 FILLER_85_819 ();
 sg13g2_decap_8 FILLER_85_834 ();
 sg13g2_fill_1 FILLER_85_841 ();
 sg13g2_decap_4 FILLER_85_848 ();
 sg13g2_fill_1 FILLER_85_852 ();
 sg13g2_fill_1 FILLER_85_863 ();
 sg13g2_fill_1 FILLER_85_875 ();
 sg13g2_fill_2 FILLER_85_890 ();
 sg13g2_fill_2 FILLER_85_898 ();
 sg13g2_decap_8 FILLER_85_936 ();
 sg13g2_decap_4 FILLER_85_943 ();
 sg13g2_decap_8 FILLER_85_952 ();
 sg13g2_decap_8 FILLER_85_959 ();
 sg13g2_fill_1 FILLER_85_966 ();
 sg13g2_decap_8 FILLER_85_973 ();
 sg13g2_decap_8 FILLER_85_980 ();
 sg13g2_fill_2 FILLER_85_987 ();
 sg13g2_fill_1 FILLER_85_989 ();
 sg13g2_decap_8 FILLER_85_995 ();
 sg13g2_decap_4 FILLER_85_1007 ();
 sg13g2_fill_1 FILLER_85_1011 ();
 sg13g2_decap_4 FILLER_85_1020 ();
 sg13g2_fill_1 FILLER_85_1060 ();
 sg13g2_fill_1 FILLER_85_1082 ();
 sg13g2_decap_8 FILLER_85_1087 ();
 sg13g2_decap_8 FILLER_85_1094 ();
 sg13g2_decap_8 FILLER_85_1101 ();
 sg13g2_decap_4 FILLER_85_1108 ();
 sg13g2_fill_2 FILLER_85_1161 ();
 sg13g2_decap_8 FILLER_85_1172 ();
 sg13g2_decap_8 FILLER_85_1179 ();
 sg13g2_decap_4 FILLER_85_1186 ();
 sg13g2_fill_1 FILLER_85_1190 ();
 sg13g2_decap_8 FILLER_85_1207 ();
 sg13g2_decap_8 FILLER_85_1214 ();
 sg13g2_decap_8 FILLER_85_1221 ();
 sg13g2_decap_8 FILLER_85_1228 ();
 sg13g2_decap_8 FILLER_85_1235 ();
 sg13g2_decap_8 FILLER_85_1242 ();
 sg13g2_decap_8 FILLER_85_1249 ();
 sg13g2_decap_4 FILLER_85_1256 ();
 sg13g2_decap_4 FILLER_85_1264 ();
 sg13g2_decap_4 FILLER_85_1345 ();
 sg13g2_fill_2 FILLER_85_1396 ();
 sg13g2_fill_1 FILLER_85_1398 ();
 sg13g2_decap_8 FILLER_85_1425 ();
 sg13g2_decap_8 FILLER_85_1432 ();
 sg13g2_decap_8 FILLER_85_1439 ();
 sg13g2_decap_4 FILLER_85_1446 ();
 sg13g2_fill_2 FILLER_85_1450 ();
 sg13g2_decap_8 FILLER_85_1478 ();
 sg13g2_decap_8 FILLER_85_1485 ();
 sg13g2_decap_4 FILLER_85_1492 ();
 sg13g2_fill_1 FILLER_85_1496 ();
 sg13g2_decap_4 FILLER_85_1594 ();
 sg13g2_fill_1 FILLER_85_1598 ();
 sg13g2_decap_8 FILLER_86_0 ();
 sg13g2_decap_8 FILLER_86_7 ();
 sg13g2_decap_8 FILLER_86_14 ();
 sg13g2_decap_8 FILLER_86_21 ();
 sg13g2_decap_8 FILLER_86_28 ();
 sg13g2_decap_8 FILLER_86_35 ();
 sg13g2_decap_8 FILLER_86_42 ();
 sg13g2_decap_8 FILLER_86_49 ();
 sg13g2_decap_8 FILLER_86_56 ();
 sg13g2_decap_8 FILLER_86_63 ();
 sg13g2_decap_8 FILLER_86_70 ();
 sg13g2_decap_8 FILLER_86_77 ();
 sg13g2_decap_8 FILLER_86_84 ();
 sg13g2_decap_8 FILLER_86_91 ();
 sg13g2_decap_8 FILLER_86_98 ();
 sg13g2_fill_2 FILLER_86_105 ();
 sg13g2_fill_1 FILLER_86_107 ();
 sg13g2_fill_2 FILLER_86_112 ();
 sg13g2_fill_1 FILLER_86_114 ();
 sg13g2_decap_8 FILLER_86_119 ();
 sg13g2_decap_8 FILLER_86_126 ();
 sg13g2_decap_8 FILLER_86_133 ();
 sg13g2_fill_2 FILLER_86_140 ();
 sg13g2_fill_1 FILLER_86_142 ();
 sg13g2_decap_8 FILLER_86_147 ();
 sg13g2_fill_2 FILLER_86_154 ();
 sg13g2_fill_1 FILLER_86_156 ();
 sg13g2_decap_4 FILLER_86_284 ();
 sg13g2_fill_1 FILLER_86_288 ();
 sg13g2_decap_8 FILLER_86_328 ();
 sg13g2_fill_1 FILLER_86_344 ();
 sg13g2_decap_8 FILLER_86_349 ();
 sg13g2_decap_8 FILLER_86_356 ();
 sg13g2_decap_8 FILLER_86_363 ();
 sg13g2_decap_8 FILLER_86_370 ();
 sg13g2_fill_2 FILLER_86_377 ();
 sg13g2_fill_1 FILLER_86_379 ();
 sg13g2_decap_8 FILLER_86_385 ();
 sg13g2_decap_8 FILLER_86_395 ();
 sg13g2_fill_2 FILLER_86_402 ();
 sg13g2_fill_1 FILLER_86_404 ();
 sg13g2_fill_1 FILLER_86_478 ();
 sg13g2_decap_8 FILLER_86_510 ();
 sg13g2_decap_8 FILLER_86_517 ();
 sg13g2_decap_8 FILLER_86_524 ();
 sg13g2_decap_8 FILLER_86_531 ();
 sg13g2_decap_8 FILLER_86_538 ();
 sg13g2_decap_8 FILLER_86_555 ();
 sg13g2_fill_1 FILLER_86_594 ();
 sg13g2_decap_8 FILLER_86_600 ();
 sg13g2_decap_8 FILLER_86_607 ();
 sg13g2_fill_1 FILLER_86_614 ();
 sg13g2_fill_1 FILLER_86_633 ();
 sg13g2_fill_1 FILLER_86_651 ();
 sg13g2_fill_2 FILLER_86_675 ();
 sg13g2_decap_8 FILLER_86_695 ();
 sg13g2_decap_8 FILLER_86_702 ();
 sg13g2_decap_8 FILLER_86_709 ();
 sg13g2_decap_8 FILLER_86_716 ();
 sg13g2_decap_8 FILLER_86_727 ();
 sg13g2_decap_8 FILLER_86_734 ();
 sg13g2_fill_2 FILLER_86_741 ();
 sg13g2_decap_4 FILLER_86_751 ();
 sg13g2_fill_2 FILLER_86_755 ();
 sg13g2_decap_4 FILLER_86_763 ();
 sg13g2_decap_4 FILLER_86_775 ();
 sg13g2_fill_2 FILLER_86_779 ();
 sg13g2_decap_8 FILLER_86_786 ();
 sg13g2_decap_4 FILLER_86_793 ();
 sg13g2_fill_1 FILLER_86_802 ();
 sg13g2_fill_1 FILLER_86_808 ();
 sg13g2_fill_1 FILLER_86_828 ();
 sg13g2_decap_8 FILLER_86_835 ();
 sg13g2_decap_8 FILLER_86_842 ();
 sg13g2_fill_1 FILLER_86_849 ();
 sg13g2_decap_8 FILLER_86_858 ();
 sg13g2_decap_8 FILLER_86_865 ();
 sg13g2_decap_8 FILLER_86_872 ();
 sg13g2_fill_2 FILLER_86_879 ();
 sg13g2_fill_1 FILLER_86_881 ();
 sg13g2_fill_1 FILLER_86_928 ();
 sg13g2_decap_8 FILLER_86_942 ();
 sg13g2_decap_8 FILLER_86_953 ();
 sg13g2_decap_8 FILLER_86_960 ();
 sg13g2_fill_1 FILLER_86_967 ();
 sg13g2_decap_8 FILLER_86_973 ();
 sg13g2_decap_8 FILLER_86_980 ();
 sg13g2_decap_8 FILLER_86_987 ();
 sg13g2_decap_8 FILLER_86_994 ();
 sg13g2_decap_8 FILLER_86_1001 ();
 sg13g2_decap_8 FILLER_86_1008 ();
 sg13g2_decap_8 FILLER_86_1015 ();
 sg13g2_fill_2 FILLER_86_1022 ();
 sg13g2_decap_8 FILLER_86_1034 ();
 sg13g2_decap_8 FILLER_86_1041 ();
 sg13g2_decap_4 FILLER_86_1048 ();
 sg13g2_decap_8 FILLER_86_1062 ();
 sg13g2_decap_8 FILLER_86_1069 ();
 sg13g2_decap_8 FILLER_86_1076 ();
 sg13g2_decap_8 FILLER_86_1083 ();
 sg13g2_decap_8 FILLER_86_1090 ();
 sg13g2_fill_1 FILLER_86_1097 ();
 sg13g2_fill_2 FILLER_86_1112 ();
 sg13g2_fill_1 FILLER_86_1114 ();
 sg13g2_decap_4 FILLER_86_1130 ();
 sg13g2_fill_1 FILLER_86_1145 ();
 sg13g2_decap_8 FILLER_86_1165 ();
 sg13g2_decap_8 FILLER_86_1172 ();
 sg13g2_decap_4 FILLER_86_1179 ();
 sg13g2_fill_2 FILLER_86_1206 ();
 sg13g2_decap_8 FILLER_86_1213 ();
 sg13g2_decap_4 FILLER_86_1220 ();
 sg13g2_fill_2 FILLER_86_1224 ();
 sg13g2_decap_8 FILLER_86_1258 ();
 sg13g2_decap_8 FILLER_86_1265 ();
 sg13g2_decap_4 FILLER_86_1272 ();
 sg13g2_decap_8 FILLER_86_1306 ();
 sg13g2_decap_8 FILLER_86_1313 ();
 sg13g2_decap_8 FILLER_86_1320 ();
 sg13g2_decap_8 FILLER_86_1327 ();
 sg13g2_fill_1 FILLER_86_1334 ();
 sg13g2_fill_2 FILLER_86_1344 ();
 sg13g2_fill_1 FILLER_86_1346 ();
 sg13g2_decap_4 FILLER_86_1351 ();
 sg13g2_fill_1 FILLER_86_1355 ();
 sg13g2_decap_8 FILLER_86_1360 ();
 sg13g2_fill_1 FILLER_86_1367 ();
 sg13g2_fill_2 FILLER_86_1389 ();
 sg13g2_decap_8 FILLER_86_1400 ();
 sg13g2_fill_2 FILLER_86_1407 ();
 sg13g2_decap_4 FILLER_86_1413 ();
 sg13g2_fill_2 FILLER_86_1417 ();
 sg13g2_decap_8 FILLER_86_1424 ();
 sg13g2_fill_1 FILLER_86_1431 ();
 sg13g2_decap_4 FILLER_86_1437 ();
 sg13g2_fill_2 FILLER_86_1441 ();
 sg13g2_fill_2 FILLER_86_1453 ();
 sg13g2_fill_1 FILLER_86_1505 ();
 sg13g2_fill_2 FILLER_86_1591 ();
 sg13g2_fill_1 FILLER_86_1593 ();
 sg13g2_fill_1 FILLER_86_1598 ();
 sg13g2_decap_8 FILLER_87_0 ();
 sg13g2_decap_8 FILLER_87_7 ();
 sg13g2_decap_8 FILLER_87_14 ();
 sg13g2_decap_8 FILLER_87_21 ();
 sg13g2_decap_8 FILLER_87_28 ();
 sg13g2_decap_8 FILLER_87_35 ();
 sg13g2_decap_8 FILLER_87_42 ();
 sg13g2_decap_8 FILLER_87_49 ();
 sg13g2_decap_8 FILLER_87_56 ();
 sg13g2_decap_8 FILLER_87_63 ();
 sg13g2_decap_8 FILLER_87_70 ();
 sg13g2_decap_8 FILLER_87_77 ();
 sg13g2_decap_8 FILLER_87_88 ();
 sg13g2_decap_4 FILLER_87_95 ();
 sg13g2_fill_2 FILLER_87_133 ();
 sg13g2_fill_2 FILLER_87_161 ();
 sg13g2_fill_2 FILLER_87_197 ();
 sg13g2_fill_1 FILLER_87_199 ();
 sg13g2_fill_2 FILLER_87_230 ();
 sg13g2_fill_1 FILLER_87_257 ();
 sg13g2_decap_8 FILLER_87_292 ();
 sg13g2_decap_8 FILLER_87_299 ();
 sg13g2_decap_4 FILLER_87_306 ();
 sg13g2_fill_2 FILLER_87_310 ();
 sg13g2_decap_4 FILLER_87_363 ();
 sg13g2_fill_1 FILLER_87_367 ();
 sg13g2_decap_8 FILLER_87_397 ();
 sg13g2_decap_4 FILLER_87_404 ();
 sg13g2_fill_2 FILLER_87_408 ();
 sg13g2_decap_8 FILLER_87_414 ();
 sg13g2_decap_8 FILLER_87_449 ();
 sg13g2_decap_8 FILLER_87_456 ();
 sg13g2_decap_8 FILLER_87_463 ();
 sg13g2_decap_8 FILLER_87_470 ();
 sg13g2_decap_8 FILLER_87_477 ();
 sg13g2_fill_2 FILLER_87_484 ();
 sg13g2_decap_8 FILLER_87_490 ();
 sg13g2_decap_8 FILLER_87_497 ();
 sg13g2_decap_8 FILLER_87_504 ();
 sg13g2_decap_8 FILLER_87_511 ();
 sg13g2_fill_2 FILLER_87_518 ();
 sg13g2_fill_1 FILLER_87_520 ();
 sg13g2_decap_8 FILLER_87_525 ();
 sg13g2_decap_8 FILLER_87_532 ();
 sg13g2_decap_4 FILLER_87_539 ();
 sg13g2_fill_1 FILLER_87_543 ();
 sg13g2_fill_1 FILLER_87_547 ();
 sg13g2_fill_1 FILLER_87_555 ();
 sg13g2_decap_4 FILLER_87_574 ();
 sg13g2_fill_1 FILLER_87_583 ();
 sg13g2_fill_2 FILLER_87_590 ();
 sg13g2_decap_4 FILLER_87_602 ();
 sg13g2_fill_2 FILLER_87_606 ();
 sg13g2_decap_8 FILLER_87_613 ();
 sg13g2_decap_8 FILLER_87_620 ();
 sg13g2_decap_8 FILLER_87_634 ();
 sg13g2_decap_8 FILLER_87_641 ();
 sg13g2_fill_1 FILLER_87_648 ();
 sg13g2_decap_8 FILLER_87_653 ();
 sg13g2_decap_4 FILLER_87_660 ();
 sg13g2_decap_8 FILLER_87_671 ();
 sg13g2_decap_8 FILLER_87_678 ();
 sg13g2_decap_8 FILLER_87_685 ();
 sg13g2_decap_8 FILLER_87_692 ();
 sg13g2_decap_8 FILLER_87_699 ();
 sg13g2_decap_4 FILLER_87_706 ();
 sg13g2_fill_2 FILLER_87_710 ();
 sg13g2_decap_8 FILLER_87_716 ();
 sg13g2_decap_8 FILLER_87_723 ();
 sg13g2_decap_8 FILLER_87_730 ();
 sg13g2_decap_8 FILLER_87_737 ();
 sg13g2_decap_8 FILLER_87_744 ();
 sg13g2_decap_8 FILLER_87_751 ();
 sg13g2_decap_4 FILLER_87_758 ();
 sg13g2_fill_1 FILLER_87_762 ();
 sg13g2_decap_8 FILLER_87_773 ();
 sg13g2_decap_8 FILLER_87_780 ();
 sg13g2_fill_2 FILLER_87_802 ();
 sg13g2_fill_1 FILLER_87_804 ();
 sg13g2_fill_2 FILLER_87_810 ();
 sg13g2_fill_2 FILLER_87_860 ();
 sg13g2_decap_8 FILLER_87_866 ();
 sg13g2_decap_8 FILLER_87_873 ();
 sg13g2_decap_8 FILLER_87_880 ();
 sg13g2_decap_8 FILLER_87_887 ();
 sg13g2_fill_2 FILLER_87_894 ();
 sg13g2_fill_1 FILLER_87_896 ();
 sg13g2_fill_2 FILLER_87_908 ();
 sg13g2_fill_1 FILLER_87_910 ();
 sg13g2_fill_2 FILLER_87_940 ();
 sg13g2_decap_4 FILLER_87_968 ();
 sg13g2_fill_1 FILLER_87_972 ();
 sg13g2_decap_8 FILLER_87_986 ();
 sg13g2_fill_1 FILLER_87_993 ();
 sg13g2_decap_4 FILLER_87_998 ();
 sg13g2_fill_2 FILLER_87_1002 ();
 sg13g2_fill_2 FILLER_87_1012 ();
 sg13g2_fill_1 FILLER_87_1014 ();
 sg13g2_decap_8 FILLER_87_1054 ();
 sg13g2_decap_8 FILLER_87_1065 ();
 sg13g2_fill_2 FILLER_87_1072 ();
 sg13g2_decap_8 FILLER_87_1082 ();
 sg13g2_decap_8 FILLER_87_1089 ();
 sg13g2_decap_8 FILLER_87_1106 ();
 sg13g2_decap_8 FILLER_87_1118 ();
 sg13g2_decap_8 FILLER_87_1125 ();
 sg13g2_decap_8 FILLER_87_1132 ();
 sg13g2_decap_8 FILLER_87_1139 ();
 sg13g2_fill_1 FILLER_87_1146 ();
 sg13g2_fill_1 FILLER_87_1174 ();
 sg13g2_decap_4 FILLER_87_1180 ();
 sg13g2_fill_1 FILLER_87_1184 ();
 sg13g2_fill_1 FILLER_87_1197 ();
 sg13g2_decap_8 FILLER_87_1209 ();
 sg13g2_fill_1 FILLER_87_1221 ();
 sg13g2_decap_4 FILLER_87_1252 ();
 sg13g2_fill_1 FILLER_87_1256 ();
 sg13g2_decap_8 FILLER_87_1272 ();
 sg13g2_fill_1 FILLER_87_1279 ();
 sg13g2_decap_8 FILLER_87_1326 ();
 sg13g2_fill_1 FILLER_87_1333 ();
 sg13g2_decap_8 FILLER_87_1360 ();
 sg13g2_decap_8 FILLER_87_1367 ();
 sg13g2_decap_8 FILLER_87_1374 ();
 sg13g2_decap_8 FILLER_87_1381 ();
 sg13g2_decap_8 FILLER_87_1388 ();
 sg13g2_fill_1 FILLER_87_1395 ();
 sg13g2_fill_1 FILLER_87_1427 ();
 sg13g2_fill_2 FILLER_87_1491 ();
 sg13g2_fill_2 FILLER_87_1514 ();
 sg13g2_decap_4 FILLER_87_1542 ();
 sg13g2_decap_8 FILLER_87_1555 ();
 sg13g2_decap_8 FILLER_87_1562 ();
 sg13g2_decap_8 FILLER_87_1569 ();
 sg13g2_decap_8 FILLER_87_1576 ();
 sg13g2_decap_8 FILLER_87_1583 ();
 sg13g2_decap_4 FILLER_87_1590 ();
 sg13g2_decap_8 FILLER_87_1599 ();
 sg13g2_decap_8 FILLER_87_1610 ();
 sg13g2_decap_8 FILLER_87_1617 ();
 sg13g2_fill_1 FILLER_87_1624 ();
 sg13g2_decap_8 FILLER_88_0 ();
 sg13g2_decap_8 FILLER_88_7 ();
 sg13g2_decap_8 FILLER_88_14 ();
 sg13g2_decap_8 FILLER_88_21 ();
 sg13g2_decap_8 FILLER_88_28 ();
 sg13g2_decap_8 FILLER_88_35 ();
 sg13g2_decap_8 FILLER_88_42 ();
 sg13g2_decap_8 FILLER_88_49 ();
 sg13g2_decap_8 FILLER_88_56 ();
 sg13g2_decap_8 FILLER_88_63 ();
 sg13g2_decap_8 FILLER_88_70 ();
 sg13g2_decap_8 FILLER_88_128 ();
 sg13g2_fill_2 FILLER_88_135 ();
 sg13g2_decap_8 FILLER_88_149 ();
 sg13g2_fill_2 FILLER_88_156 ();
 sg13g2_decap_4 FILLER_88_191 ();
 sg13g2_fill_2 FILLER_88_220 ();
 sg13g2_fill_1 FILLER_88_222 ();
 sg13g2_fill_2 FILLER_88_253 ();
 sg13g2_decap_8 FILLER_88_293 ();
 sg13g2_decap_8 FILLER_88_300 ();
 sg13g2_decap_4 FILLER_88_307 ();
 sg13g2_decap_8 FILLER_88_337 ();
 sg13g2_decap_8 FILLER_88_344 ();
 sg13g2_fill_2 FILLER_88_351 ();
 sg13g2_fill_1 FILLER_88_353 ();
 sg13g2_decap_8 FILLER_88_401 ();
 sg13g2_decap_8 FILLER_88_408 ();
 sg13g2_decap_4 FILLER_88_415 ();
 sg13g2_fill_1 FILLER_88_419 ();
 sg13g2_decap_8 FILLER_88_425 ();
 sg13g2_fill_2 FILLER_88_432 ();
 sg13g2_fill_1 FILLER_88_434 ();
 sg13g2_decap_4 FILLER_88_443 ();
 sg13g2_fill_1 FILLER_88_447 ();
 sg13g2_fill_1 FILLER_88_473 ();
 sg13g2_decap_4 FILLER_88_509 ();
 sg13g2_fill_1 FILLER_88_513 ();
 sg13g2_decap_4 FILLER_88_540 ();
 sg13g2_decap_8 FILLER_88_558 ();
 sg13g2_fill_2 FILLER_88_565 ();
 sg13g2_fill_1 FILLER_88_567 ();
 sg13g2_decap_8 FILLER_88_575 ();
 sg13g2_decap_8 FILLER_88_582 ();
 sg13g2_decap_8 FILLER_88_589 ();
 sg13g2_fill_1 FILLER_88_596 ();
 sg13g2_decap_4 FILLER_88_602 ();
 sg13g2_fill_1 FILLER_88_606 ();
 sg13g2_fill_2 FILLER_88_612 ();
 sg13g2_fill_1 FILLER_88_614 ();
 sg13g2_fill_2 FILLER_88_634 ();
 sg13g2_fill_1 FILLER_88_636 ();
 sg13g2_fill_2 FILLER_88_673 ();
 sg13g2_fill_2 FILLER_88_680 ();
 sg13g2_fill_1 FILLER_88_682 ();
 sg13g2_fill_2 FILLER_88_704 ();
 sg13g2_decap_8 FILLER_88_732 ();
 sg13g2_decap_4 FILLER_88_739 ();
 sg13g2_fill_2 FILLER_88_743 ();
 sg13g2_decap_8 FILLER_88_750 ();
 sg13g2_decap_8 FILLER_88_757 ();
 sg13g2_fill_1 FILLER_88_769 ();
 sg13g2_decap_8 FILLER_88_775 ();
 sg13g2_fill_2 FILLER_88_782 ();
 sg13g2_fill_1 FILLER_88_784 ();
 sg13g2_decap_8 FILLER_88_790 ();
 sg13g2_decap_8 FILLER_88_801 ();
 sg13g2_decap_8 FILLER_88_808 ();
 sg13g2_fill_1 FILLER_88_815 ();
 sg13g2_decap_8 FILLER_88_821 ();
 sg13g2_decap_8 FILLER_88_828 ();
 sg13g2_decap_4 FILLER_88_876 ();
 sg13g2_fill_2 FILLER_88_880 ();
 sg13g2_fill_2 FILLER_88_887 ();
 sg13g2_fill_1 FILLER_88_889 ();
 sg13g2_decap_4 FILLER_88_899 ();
 sg13g2_fill_2 FILLER_88_903 ();
 sg13g2_decap_4 FILLER_88_956 ();
 sg13g2_decap_8 FILLER_88_970 ();
 sg13g2_fill_1 FILLER_88_977 ();
 sg13g2_decap_4 FILLER_88_982 ();
 sg13g2_fill_2 FILLER_88_986 ();
 sg13g2_decap_8 FILLER_88_1019 ();
 sg13g2_fill_2 FILLER_88_1030 ();
 sg13g2_fill_2 FILLER_88_1058 ();
 sg13g2_fill_1 FILLER_88_1060 ();
 sg13g2_decap_8 FILLER_88_1090 ();
 sg13g2_decap_4 FILLER_88_1097 ();
 sg13g2_fill_2 FILLER_88_1101 ();
 sg13g2_decap_8 FILLER_88_1117 ();
 sg13g2_decap_8 FILLER_88_1124 ();
 sg13g2_decap_8 FILLER_88_1131 ();
 sg13g2_decap_8 FILLER_88_1138 ();
 sg13g2_fill_2 FILLER_88_1145 ();
 sg13g2_decap_8 FILLER_88_1168 ();
 sg13g2_decap_8 FILLER_88_1175 ();
 sg13g2_decap_4 FILLER_88_1182 ();
 sg13g2_decap_4 FILLER_88_1192 ();
 sg13g2_fill_1 FILLER_88_1196 ();
 sg13g2_decap_8 FILLER_88_1202 ();
 sg13g2_decap_8 FILLER_88_1209 ();
 sg13g2_decap_8 FILLER_88_1228 ();
 sg13g2_decap_8 FILLER_88_1235 ();
 sg13g2_decap_8 FILLER_88_1242 ();
 sg13g2_fill_2 FILLER_88_1249 ();
 sg13g2_fill_1 FILLER_88_1251 ();
 sg13g2_decap_4 FILLER_88_1278 ();
 sg13g2_fill_1 FILLER_88_1282 ();
 sg13g2_decap_8 FILLER_88_1304 ();
 sg13g2_decap_8 FILLER_88_1311 ();
 sg13g2_fill_2 FILLER_88_1318 ();
 sg13g2_decap_8 FILLER_88_1354 ();
 sg13g2_decap_4 FILLER_88_1361 ();
 sg13g2_decap_8 FILLER_88_1396 ();
 sg13g2_decap_8 FILLER_88_1474 ();
 sg13g2_decap_8 FILLER_88_1481 ();
 sg13g2_fill_1 FILLER_88_1488 ();
 sg13g2_fill_1 FILLER_88_1510 ();
 sg13g2_fill_2 FILLER_88_1532 ();
 sg13g2_fill_1 FILLER_88_1534 ();
 sg13g2_fill_2 FILLER_88_1540 ();
 sg13g2_decap_8 FILLER_88_1546 ();
 sg13g2_decap_8 FILLER_88_1553 ();
 sg13g2_fill_2 FILLER_88_1560 ();
 sg13g2_fill_1 FILLER_88_1562 ();
 sg13g2_fill_2 FILLER_88_1568 ();
 sg13g2_decap_4 FILLER_88_1574 ();
 sg13g2_fill_2 FILLER_88_1578 ();
 sg13g2_decap_8 FILLER_88_1589 ();
 sg13g2_decap_8 FILLER_88_1596 ();
 sg13g2_decap_8 FILLER_88_1603 ();
 sg13g2_decap_8 FILLER_88_1610 ();
 sg13g2_decap_8 FILLER_88_1617 ();
 sg13g2_fill_1 FILLER_88_1624 ();
 sg13g2_decap_8 FILLER_89_0 ();
 sg13g2_decap_8 FILLER_89_7 ();
 sg13g2_decap_8 FILLER_89_14 ();
 sg13g2_decap_8 FILLER_89_21 ();
 sg13g2_decap_8 FILLER_89_28 ();
 sg13g2_decap_8 FILLER_89_35 ();
 sg13g2_decap_8 FILLER_89_42 ();
 sg13g2_decap_8 FILLER_89_49 ();
 sg13g2_decap_8 FILLER_89_56 ();
 sg13g2_decap_8 FILLER_89_63 ();
 sg13g2_decap_8 FILLER_89_70 ();
 sg13g2_decap_8 FILLER_89_77 ();
 sg13g2_decap_8 FILLER_89_84 ();
 sg13g2_decap_8 FILLER_89_91 ();
 sg13g2_decap_4 FILLER_89_114 ();
 sg13g2_decap_8 FILLER_89_122 ();
 sg13g2_fill_2 FILLER_89_129 ();
 sg13g2_fill_1 FILLER_89_139 ();
 sg13g2_decap_8 FILLER_89_145 ();
 sg13g2_fill_2 FILLER_89_152 ();
 sg13g2_fill_1 FILLER_89_154 ();
 sg13g2_decap_8 FILLER_89_184 ();
 sg13g2_decap_8 FILLER_89_191 ();
 sg13g2_decap_4 FILLER_89_198 ();
 sg13g2_decap_4 FILLER_89_226 ();
 sg13g2_fill_2 FILLER_89_230 ();
 sg13g2_fill_1 FILLER_89_257 ();
 sg13g2_fill_2 FILLER_89_262 ();
 sg13g2_decap_8 FILLER_89_268 ();
 sg13g2_decap_8 FILLER_89_275 ();
 sg13g2_decap_8 FILLER_89_282 ();
 sg13g2_decap_4 FILLER_89_289 ();
 sg13g2_fill_1 FILLER_89_293 ();
 sg13g2_decap_8 FILLER_89_303 ();
 sg13g2_decap_8 FILLER_89_310 ();
 sg13g2_fill_1 FILLER_89_317 ();
 sg13g2_decap_8 FILLER_89_322 ();
 sg13g2_fill_2 FILLER_89_329 ();
 sg13g2_decap_4 FILLER_89_345 ();
 sg13g2_fill_2 FILLER_89_353 ();
 sg13g2_decap_8 FILLER_89_376 ();
 sg13g2_decap_8 FILLER_89_387 ();
 sg13g2_fill_2 FILLER_89_394 ();
 sg13g2_fill_1 FILLER_89_396 ();
 sg13g2_fill_2 FILLER_89_418 ();
 sg13g2_fill_1 FILLER_89_420 ();
 sg13g2_decap_8 FILLER_89_473 ();
 sg13g2_decap_4 FILLER_89_480 ();
 sg13g2_fill_1 FILLER_89_493 ();
 sg13g2_decap_8 FILLER_89_520 ();
 sg13g2_decap_8 FILLER_89_527 ();
 sg13g2_decap_8 FILLER_89_534 ();
 sg13g2_decap_4 FILLER_89_541 ();
 sg13g2_decap_4 FILLER_89_578 ();
 sg13g2_fill_1 FILLER_89_582 ();
 sg13g2_decap_4 FILLER_89_588 ();
 sg13g2_fill_1 FILLER_89_592 ();
 sg13g2_decap_4 FILLER_89_613 ();
 sg13g2_fill_2 FILLER_89_617 ();
 sg13g2_decap_8 FILLER_89_633 ();
 sg13g2_decap_8 FILLER_89_640 ();
 sg13g2_decap_8 FILLER_89_647 ();
 sg13g2_fill_2 FILLER_89_654 ();
 sg13g2_fill_1 FILLER_89_656 ();
 sg13g2_decap_4 FILLER_89_661 ();
 sg13g2_decap_8 FILLER_89_673 ();
 sg13g2_fill_2 FILLER_89_680 ();
 sg13g2_fill_2 FILLER_89_687 ();
 sg13g2_decap_8 FILLER_89_701 ();
 sg13g2_fill_2 FILLER_89_708 ();
 sg13g2_decap_8 FILLER_89_762 ();
 sg13g2_decap_8 FILLER_89_769 ();
 sg13g2_decap_8 FILLER_89_780 ();
 sg13g2_fill_2 FILLER_89_787 ();
 sg13g2_decap_8 FILLER_89_820 ();
 sg13g2_decap_8 FILLER_89_827 ();
 sg13g2_decap_8 FILLER_89_834 ();
 sg13g2_decap_4 FILLER_89_841 ();
 sg13g2_decap_8 FILLER_89_881 ();
 sg13g2_decap_4 FILLER_89_888 ();
 sg13g2_fill_1 FILLER_89_892 ();
 sg13g2_fill_2 FILLER_89_903 ();
 sg13g2_fill_1 FILLER_89_905 ();
 sg13g2_fill_2 FILLER_89_914 ();
 sg13g2_decap_8 FILLER_89_951 ();
 sg13g2_decap_8 FILLER_89_958 ();
 sg13g2_decap_4 FILLER_89_965 ();
 sg13g2_fill_2 FILLER_89_969 ();
 sg13g2_decap_8 FILLER_89_997 ();
 sg13g2_decap_8 FILLER_89_1004 ();
 sg13g2_decap_8 FILLER_89_1011 ();
 sg13g2_fill_2 FILLER_89_1018 ();
 sg13g2_decap_4 FILLER_89_1024 ();
 sg13g2_decap_8 FILLER_89_1033 ();
 sg13g2_decap_8 FILLER_89_1044 ();
 sg13g2_fill_1 FILLER_89_1051 ();
 sg13g2_decap_8 FILLER_89_1083 ();
 sg13g2_decap_8 FILLER_89_1090 ();
 sg13g2_decap_4 FILLER_89_1097 ();
 sg13g2_fill_1 FILLER_89_1101 ();
 sg13g2_fill_1 FILLER_89_1107 ();
 sg13g2_decap_8 FILLER_89_1113 ();
 sg13g2_decap_8 FILLER_89_1120 ();
 sg13g2_decap_4 FILLER_89_1127 ();
 sg13g2_fill_2 FILLER_89_1131 ();
 sg13g2_decap_8 FILLER_89_1143 ();
 sg13g2_decap_4 FILLER_89_1150 ();
 sg13g2_decap_8 FILLER_89_1159 ();
 sg13g2_fill_2 FILLER_89_1166 ();
 sg13g2_decap_4 FILLER_89_1172 ();
 sg13g2_decap_8 FILLER_89_1210 ();
 sg13g2_fill_1 FILLER_89_1241 ();
 sg13g2_decap_4 FILLER_89_1246 ();
 sg13g2_fill_1 FILLER_89_1250 ();
 sg13g2_decap_8 FILLER_89_1306 ();
 sg13g2_fill_1 FILLER_89_1313 ();
 sg13g2_decap_8 FILLER_89_1344 ();
 sg13g2_decap_8 FILLER_89_1351 ();
 sg13g2_decap_8 FILLER_89_1358 ();
 sg13g2_decap_8 FILLER_89_1365 ();
 sg13g2_decap_8 FILLER_89_1372 ();
 sg13g2_decap_8 FILLER_89_1379 ();
 sg13g2_fill_1 FILLER_89_1395 ();
 sg13g2_decap_8 FILLER_89_1400 ();
 sg13g2_decap_8 FILLER_89_1407 ();
 sg13g2_fill_1 FILLER_89_1414 ();
 sg13g2_decap_8 FILLER_89_1436 ();
 sg13g2_decap_8 FILLER_89_1443 ();
 sg13g2_decap_8 FILLER_89_1450 ();
 sg13g2_decap_8 FILLER_89_1457 ();
 sg13g2_decap_8 FILLER_89_1464 ();
 sg13g2_decap_8 FILLER_89_1471 ();
 sg13g2_decap_8 FILLER_89_1478 ();
 sg13g2_decap_8 FILLER_89_1485 ();
 sg13g2_decap_4 FILLER_89_1492 ();
 sg13g2_decap_8 FILLER_89_1500 ();
 sg13g2_decap_4 FILLER_89_1507 ();
 sg13g2_fill_1 FILLER_89_1511 ();
 sg13g2_fill_2 FILLER_89_1533 ();
 sg13g2_fill_1 FILLER_89_1535 ();
 sg13g2_decap_8 FILLER_89_1588 ();
 sg13g2_decap_8 FILLER_89_1595 ();
 sg13g2_decap_8 FILLER_89_1602 ();
 sg13g2_decap_8 FILLER_89_1609 ();
 sg13g2_decap_8 FILLER_89_1616 ();
 sg13g2_fill_2 FILLER_89_1623 ();
 sg13g2_decap_8 FILLER_90_0 ();
 sg13g2_decap_8 FILLER_90_7 ();
 sg13g2_decap_8 FILLER_90_14 ();
 sg13g2_decap_8 FILLER_90_21 ();
 sg13g2_decap_8 FILLER_90_28 ();
 sg13g2_decap_8 FILLER_90_35 ();
 sg13g2_decap_8 FILLER_90_42 ();
 sg13g2_decap_8 FILLER_90_49 ();
 sg13g2_decap_8 FILLER_90_56 ();
 sg13g2_decap_8 FILLER_90_63 ();
 sg13g2_decap_8 FILLER_90_70 ();
 sg13g2_decap_8 FILLER_90_77 ();
 sg13g2_fill_1 FILLER_90_84 ();
 sg13g2_decap_8 FILLER_90_89 ();
 sg13g2_decap_8 FILLER_90_96 ();
 sg13g2_decap_8 FILLER_90_103 ();
 sg13g2_decap_4 FILLER_90_110 ();
 sg13g2_fill_2 FILLER_90_114 ();
 sg13g2_fill_1 FILLER_90_122 ();
 sg13g2_decap_4 FILLER_90_127 ();
 sg13g2_fill_2 FILLER_90_131 ();
 sg13g2_decap_8 FILLER_90_138 ();
 sg13g2_fill_2 FILLER_90_192 ();
 sg13g2_fill_1 FILLER_90_194 ();
 sg13g2_decap_4 FILLER_90_200 ();
 sg13g2_fill_1 FILLER_90_216 ();
 sg13g2_decap_8 FILLER_90_222 ();
 sg13g2_decap_8 FILLER_90_229 ();
 sg13g2_decap_8 FILLER_90_236 ();
 sg13g2_decap_8 FILLER_90_243 ();
 sg13g2_fill_1 FILLER_90_250 ();
 sg13g2_decap_4 FILLER_90_277 ();
 sg13g2_fill_2 FILLER_90_281 ();
 sg13g2_fill_2 FILLER_90_287 ();
 sg13g2_fill_1 FILLER_90_289 ();
 sg13g2_decap_8 FILLER_90_316 ();
 sg13g2_decap_4 FILLER_90_323 ();
 sg13g2_fill_2 FILLER_90_327 ();
 sg13g2_decap_8 FILLER_90_355 ();
 sg13g2_decap_8 FILLER_90_362 ();
 sg13g2_decap_8 FILLER_90_369 ();
 sg13g2_decap_8 FILLER_90_376 ();
 sg13g2_decap_8 FILLER_90_383 ();
 sg13g2_decap_8 FILLER_90_390 ();
 sg13g2_decap_8 FILLER_90_418 ();
 sg13g2_fill_2 FILLER_90_425 ();
 sg13g2_fill_1 FILLER_90_427 ();
 sg13g2_decap_8 FILLER_90_432 ();
 sg13g2_decap_8 FILLER_90_439 ();
 sg13g2_decap_8 FILLER_90_446 ();
 sg13g2_decap_4 FILLER_90_453 ();
 sg13g2_decap_8 FILLER_90_517 ();
 sg13g2_decap_8 FILLER_90_524 ();
 sg13g2_decap_8 FILLER_90_531 ();
 sg13g2_decap_4 FILLER_90_538 ();
 sg13g2_fill_1 FILLER_90_554 ();
 sg13g2_decap_8 FILLER_90_563 ();
 sg13g2_decap_8 FILLER_90_570 ();
 sg13g2_fill_2 FILLER_90_577 ();
 sg13g2_decap_8 FILLER_90_584 ();
 sg13g2_decap_8 FILLER_90_591 ();
 sg13g2_fill_1 FILLER_90_598 ();
 sg13g2_decap_8 FILLER_90_615 ();
 sg13g2_decap_8 FILLER_90_622 ();
 sg13g2_fill_1 FILLER_90_629 ();
 sg13g2_fill_2 FILLER_90_665 ();
 sg13g2_fill_2 FILLER_90_672 ();
 sg13g2_decap_4 FILLER_90_679 ();
 sg13g2_fill_2 FILLER_90_683 ();
 sg13g2_decap_8 FILLER_90_693 ();
 sg13g2_decap_8 FILLER_90_700 ();
 sg13g2_decap_8 FILLER_90_707 ();
 sg13g2_fill_2 FILLER_90_714 ();
 sg13g2_fill_1 FILLER_90_716 ();
 sg13g2_decap_8 FILLER_90_721 ();
 sg13g2_decap_8 FILLER_90_728 ();
 sg13g2_fill_2 FILLER_90_735 ();
 sg13g2_fill_1 FILLER_90_737 ();
 sg13g2_decap_8 FILLER_90_751 ();
 sg13g2_decap_8 FILLER_90_758 ();
 sg13g2_decap_4 FILLER_90_765 ();
 sg13g2_fill_2 FILLER_90_795 ();
 sg13g2_decap_4 FILLER_90_802 ();
 sg13g2_fill_2 FILLER_90_806 ();
 sg13g2_decap_8 FILLER_90_813 ();
 sg13g2_fill_1 FILLER_90_820 ();
 sg13g2_fill_1 FILLER_90_830 ();
 sg13g2_fill_1 FILLER_90_839 ();
 sg13g2_fill_2 FILLER_90_869 ();
 sg13g2_decap_4 FILLER_90_879 ();
 sg13g2_fill_2 FILLER_90_883 ();
 sg13g2_fill_1 FILLER_90_922 ();
 sg13g2_fill_1 FILLER_90_927 ();
 sg13g2_fill_1 FILLER_90_944 ();
 sg13g2_decap_4 FILLER_90_970 ();
 sg13g2_decap_4 FILLER_90_979 ();
 sg13g2_fill_1 FILLER_90_983 ();
 sg13g2_decap_8 FILLER_90_994 ();
 sg13g2_fill_1 FILLER_90_1001 ();
 sg13g2_decap_4 FILLER_90_1012 ();
 sg13g2_fill_1 FILLER_90_1016 ();
 sg13g2_decap_4 FILLER_90_1032 ();
 sg13g2_fill_1 FILLER_90_1036 ();
 sg13g2_decap_8 FILLER_90_1041 ();
 sg13g2_decap_8 FILLER_90_1048 ();
 sg13g2_decap_8 FILLER_90_1055 ();
 sg13g2_decap_8 FILLER_90_1062 ();
 sg13g2_decap_8 FILLER_90_1069 ();
 sg13g2_decap_8 FILLER_90_1126 ();
 sg13g2_fill_2 FILLER_90_1133 ();
 sg13g2_decap_8 FILLER_90_1152 ();
 sg13g2_fill_2 FILLER_90_1159 ();
 sg13g2_decap_8 FILLER_90_1218 ();
 sg13g2_fill_2 FILLER_90_1225 ();
 sg13g2_fill_1 FILLER_90_1227 ();
 sg13g2_fill_2 FILLER_90_1254 ();
 sg13g2_decap_8 FILLER_90_1285 ();
 sg13g2_decap_4 FILLER_90_1292 ();
 sg13g2_decap_8 FILLER_90_1317 ();
 sg13g2_decap_4 FILLER_90_1324 ();
 sg13g2_fill_1 FILLER_90_1328 ();
 sg13g2_fill_1 FILLER_90_1332 ();
 sg13g2_fill_2 FILLER_90_1338 ();
 sg13g2_fill_1 FILLER_90_1340 ();
 sg13g2_decap_4 FILLER_90_1383 ();
 sg13g2_fill_1 FILLER_90_1387 ();
 sg13g2_decap_8 FILLER_90_1414 ();
 sg13g2_fill_2 FILLER_90_1421 ();
 sg13g2_fill_1 FILLER_90_1423 ();
 sg13g2_decap_8 FILLER_90_1453 ();
 sg13g2_decap_8 FILLER_90_1460 ();
 sg13g2_fill_1 FILLER_90_1467 ();
 sg13g2_decap_4 FILLER_90_1473 ();
 sg13g2_fill_1 FILLER_90_1477 ();
 sg13g2_decap_8 FILLER_90_1482 ();
 sg13g2_decap_8 FILLER_90_1515 ();
 sg13g2_decap_8 FILLER_90_1522 ();
 sg13g2_decap_8 FILLER_90_1529 ();
 sg13g2_decap_8 FILLER_90_1540 ();
 sg13g2_decap_8 FILLER_90_1547 ();
 sg13g2_decap_4 FILLER_90_1554 ();
 sg13g2_fill_2 FILLER_90_1558 ();
 sg13g2_decap_4 FILLER_90_1564 ();
 sg13g2_decap_8 FILLER_90_1572 ();
 sg13g2_decap_4 FILLER_90_1579 ();
 sg13g2_fill_1 FILLER_90_1583 ();
 sg13g2_decap_8 FILLER_90_1610 ();
 sg13g2_decap_8 FILLER_90_1617 ();
 sg13g2_fill_1 FILLER_90_1624 ();
 sg13g2_decap_8 FILLER_91_0 ();
 sg13g2_decap_8 FILLER_91_7 ();
 sg13g2_decap_8 FILLER_91_14 ();
 sg13g2_decap_8 FILLER_91_21 ();
 sg13g2_decap_8 FILLER_91_28 ();
 sg13g2_decap_8 FILLER_91_35 ();
 sg13g2_decap_8 FILLER_91_42 ();
 sg13g2_decap_8 FILLER_91_49 ();
 sg13g2_decap_4 FILLER_91_56 ();
 sg13g2_fill_2 FILLER_91_60 ();
 sg13g2_decap_8 FILLER_91_66 ();
 sg13g2_decap_4 FILLER_91_73 ();
 sg13g2_fill_2 FILLER_91_77 ();
 sg13g2_fill_2 FILLER_91_110 ();
 sg13g2_decap_8 FILLER_91_138 ();
 sg13g2_decap_4 FILLER_91_145 ();
 sg13g2_fill_1 FILLER_91_160 ();
 sg13g2_decap_8 FILLER_91_199 ();
 sg13g2_decap_4 FILLER_91_206 ();
 sg13g2_fill_2 FILLER_91_219 ();
 sg13g2_decap_8 FILLER_91_255 ();
 sg13g2_decap_8 FILLER_91_262 ();
 sg13g2_decap_8 FILLER_91_269 ();
 sg13g2_fill_1 FILLER_91_276 ();
 sg13g2_decap_4 FILLER_91_306 ();
 sg13g2_fill_2 FILLER_91_310 ();
 sg13g2_decap_8 FILLER_91_325 ();
 sg13g2_decap_8 FILLER_91_332 ();
 sg13g2_decap_8 FILLER_91_339 ();
 sg13g2_decap_8 FILLER_91_346 ();
 sg13g2_decap_8 FILLER_91_353 ();
 sg13g2_fill_2 FILLER_91_360 ();
 sg13g2_fill_2 FILLER_91_371 ();
 sg13g2_decap_4 FILLER_91_377 ();
 sg13g2_fill_2 FILLER_91_381 ();
 sg13g2_decap_8 FILLER_91_388 ();
 sg13g2_fill_2 FILLER_91_395 ();
 sg13g2_fill_1 FILLER_91_406 ();
 sg13g2_decap_8 FILLER_91_411 ();
 sg13g2_decap_8 FILLER_91_418 ();
 sg13g2_fill_2 FILLER_91_425 ();
 sg13g2_fill_1 FILLER_91_427 ();
 sg13g2_decap_8 FILLER_91_433 ();
 sg13g2_decap_8 FILLER_91_440 ();
 sg13g2_fill_2 FILLER_91_447 ();
 sg13g2_fill_1 FILLER_91_449 ();
 sg13g2_decap_8 FILLER_91_454 ();
 sg13g2_decap_8 FILLER_91_461 ();
 sg13g2_decap_4 FILLER_91_468 ();
 sg13g2_fill_2 FILLER_91_472 ();
 sg13g2_decap_8 FILLER_91_478 ();
 sg13g2_decap_8 FILLER_91_485 ();
 sg13g2_decap_8 FILLER_91_492 ();
 sg13g2_decap_8 FILLER_91_503 ();
 sg13g2_decap_8 FILLER_91_510 ();
 sg13g2_decap_8 FILLER_91_517 ();
 sg13g2_decap_8 FILLER_91_524 ();
 sg13g2_decap_8 FILLER_91_531 ();
 sg13g2_decap_8 FILLER_91_538 ();
 sg13g2_decap_8 FILLER_91_545 ();
 sg13g2_fill_2 FILLER_91_552 ();
 sg13g2_fill_1 FILLER_91_554 ();
 sg13g2_decap_4 FILLER_91_564 ();
 sg13g2_fill_2 FILLER_91_568 ();
 sg13g2_decap_4 FILLER_91_575 ();
 sg13g2_fill_2 FILLER_91_579 ();
 sg13g2_fill_1 FILLER_91_589 ();
 sg13g2_fill_1 FILLER_91_599 ();
 sg13g2_decap_8 FILLER_91_610 ();
 sg13g2_decap_8 FILLER_91_617 ();
 sg13g2_fill_2 FILLER_91_624 ();
 sg13g2_decap_8 FILLER_91_631 ();
 sg13g2_decap_8 FILLER_91_638 ();
 sg13g2_decap_8 FILLER_91_645 ();
 sg13g2_fill_1 FILLER_91_652 ();
 sg13g2_decap_8 FILLER_91_664 ();
 sg13g2_decap_4 FILLER_91_671 ();
 sg13g2_decap_4 FILLER_91_690 ();
 sg13g2_fill_1 FILLER_91_694 ();
 sg13g2_decap_4 FILLER_91_701 ();
 sg13g2_decap_8 FILLER_91_716 ();
 sg13g2_decap_8 FILLER_91_723 ();
 sg13g2_decap_4 FILLER_91_730 ();
 sg13g2_fill_1 FILLER_91_734 ();
 sg13g2_decap_8 FILLER_91_740 ();
 sg13g2_fill_2 FILLER_91_751 ();
 sg13g2_decap_4 FILLER_91_759 ();
 sg13g2_fill_1 FILLER_91_763 ();
 sg13g2_fill_1 FILLER_91_769 ();
 sg13g2_fill_2 FILLER_91_865 ();
 sg13g2_fill_1 FILLER_91_902 ();
 sg13g2_fill_1 FILLER_91_908 ();
 sg13g2_decap_8 FILLER_91_946 ();
 sg13g2_decap_4 FILLER_91_953 ();
 sg13g2_fill_1 FILLER_91_957 ();
 sg13g2_decap_8 FILLER_91_963 ();
 sg13g2_decap_8 FILLER_91_970 ();
 sg13g2_decap_8 FILLER_91_977 ();
 sg13g2_decap_8 FILLER_91_984 ();
 sg13g2_decap_8 FILLER_91_991 ();
 sg13g2_decap_4 FILLER_91_998 ();
 sg13g2_fill_1 FILLER_91_1028 ();
 sg13g2_fill_2 FILLER_91_1060 ();
 sg13g2_fill_1 FILLER_91_1062 ();
 sg13g2_fill_2 FILLER_91_1075 ();
 sg13g2_decap_4 FILLER_91_1102 ();
 sg13g2_decap_8 FILLER_91_1116 ();
 sg13g2_decap_8 FILLER_91_1123 ();
 sg13g2_decap_4 FILLER_91_1130 ();
 sg13g2_fill_2 FILLER_91_1134 ();
 sg13g2_fill_2 FILLER_91_1145 ();
 sg13g2_decap_8 FILLER_91_1156 ();
 sg13g2_decap_8 FILLER_91_1163 ();
 sg13g2_decap_4 FILLER_91_1170 ();
 sg13g2_fill_1 FILLER_91_1174 ();
 sg13g2_decap_4 FILLER_91_1180 ();
 sg13g2_fill_2 FILLER_91_1184 ();
 sg13g2_decap_4 FILLER_91_1195 ();
 sg13g2_fill_1 FILLER_91_1199 ();
 sg13g2_decap_8 FILLER_91_1204 ();
 sg13g2_decap_8 FILLER_91_1211 ();
 sg13g2_fill_1 FILLER_91_1232 ();
 sg13g2_decap_8 FILLER_91_1258 ();
 sg13g2_fill_1 FILLER_91_1265 ();
 sg13g2_decap_8 FILLER_91_1274 ();
 sg13g2_fill_2 FILLER_91_1281 ();
 sg13g2_fill_1 FILLER_91_1283 ();
 sg13g2_decap_8 FILLER_91_1309 ();
 sg13g2_decap_8 FILLER_91_1316 ();
 sg13g2_decap_8 FILLER_91_1323 ();
 sg13g2_fill_2 FILLER_91_1330 ();
 sg13g2_fill_2 FILLER_91_1337 ();
 sg13g2_fill_1 FILLER_91_1339 ();
 sg13g2_decap_8 FILLER_91_1366 ();
 sg13g2_decap_8 FILLER_91_1373 ();
 sg13g2_fill_2 FILLER_91_1380 ();
 sg13g2_fill_1 FILLER_91_1382 ();
 sg13g2_fill_2 FILLER_91_1387 ();
 sg13g2_fill_1 FILLER_91_1389 ();
 sg13g2_decap_8 FILLER_91_1419 ();
 sg13g2_fill_2 FILLER_91_1426 ();
 sg13g2_fill_1 FILLER_91_1489 ();
 sg13g2_decap_8 FILLER_91_1499 ();
 sg13g2_decap_8 FILLER_91_1506 ();
 sg13g2_decap_4 FILLER_91_1513 ();
 sg13g2_fill_2 FILLER_91_1517 ();
 sg13g2_decap_8 FILLER_91_1540 ();
 sg13g2_decap_8 FILLER_91_1572 ();
 sg13g2_decap_8 FILLER_91_1579 ();
 sg13g2_decap_4 FILLER_91_1586 ();
 sg13g2_fill_2 FILLER_91_1590 ();
 sg13g2_decap_8 FILLER_91_1596 ();
 sg13g2_decap_8 FILLER_91_1603 ();
 sg13g2_decap_8 FILLER_91_1610 ();
 sg13g2_decap_8 FILLER_91_1617 ();
 sg13g2_fill_1 FILLER_91_1624 ();
 sg13g2_decap_8 FILLER_92_0 ();
 sg13g2_decap_8 FILLER_92_7 ();
 sg13g2_decap_8 FILLER_92_14 ();
 sg13g2_decap_8 FILLER_92_21 ();
 sg13g2_decap_8 FILLER_92_28 ();
 sg13g2_decap_8 FILLER_92_35 ();
 sg13g2_decap_8 FILLER_92_42 ();
 sg13g2_decap_4 FILLER_92_49 ();
 sg13g2_fill_2 FILLER_92_53 ();
 sg13g2_fill_2 FILLER_92_81 ();
 sg13g2_fill_2 FILLER_92_98 ();
 sg13g2_fill_1 FILLER_92_100 ();
 sg13g2_decap_4 FILLER_92_111 ();
 sg13g2_decap_8 FILLER_92_125 ();
 sg13g2_decap_8 FILLER_92_132 ();
 sg13g2_decap_4 FILLER_92_184 ();
 sg13g2_decap_4 FILLER_92_214 ();
 sg13g2_fill_2 FILLER_92_218 ();
 sg13g2_decap_8 FILLER_92_224 ();
 sg13g2_fill_1 FILLER_92_231 ();
 sg13g2_decap_8 FILLER_92_236 ();
 sg13g2_fill_2 FILLER_92_243 ();
 sg13g2_fill_1 FILLER_92_245 ();
 sg13g2_decap_8 FILLER_92_300 ();
 sg13g2_fill_2 FILLER_92_307 ();
 sg13g2_fill_1 FILLER_92_309 ();
 sg13g2_decap_8 FILLER_92_336 ();
 sg13g2_decap_4 FILLER_92_343 ();
 sg13g2_fill_2 FILLER_92_347 ();
 sg13g2_decap_4 FILLER_92_358 ();
 sg13g2_fill_2 FILLER_92_362 ();
 sg13g2_decap_4 FILLER_92_390 ();
 sg13g2_decap_4 FILLER_92_424 ();
 sg13g2_fill_2 FILLER_92_428 ();
 sg13g2_decap_8 FILLER_92_456 ();
 sg13g2_decap_4 FILLER_92_463 ();
 sg13g2_fill_1 FILLER_92_467 ();
 sg13g2_decap_4 FILLER_92_472 ();
 sg13g2_decap_8 FILLER_92_485 ();
 sg13g2_decap_4 FILLER_92_527 ();
 sg13g2_decap_8 FILLER_92_546 ();
 sg13g2_fill_1 FILLER_92_553 ();
 sg13g2_decap_8 FILLER_92_562 ();
 sg13g2_decap_8 FILLER_92_569 ();
 sg13g2_decap_8 FILLER_92_576 ();
 sg13g2_decap_8 FILLER_92_583 ();
 sg13g2_decap_8 FILLER_92_590 ();
 sg13g2_decap_4 FILLER_92_597 ();
 sg13g2_fill_2 FILLER_92_601 ();
 sg13g2_decap_4 FILLER_92_613 ();
 sg13g2_fill_2 FILLER_92_631 ();
 sg13g2_fill_2 FILLER_92_642 ();
 sg13g2_fill_1 FILLER_92_644 ();
 sg13g2_fill_1 FILLER_92_648 ();
 sg13g2_fill_2 FILLER_92_654 ();
 sg13g2_fill_1 FILLER_92_656 ();
 sg13g2_decap_8 FILLER_92_672 ();
 sg13g2_decap_4 FILLER_92_679 ();
 sg13g2_decap_4 FILLER_92_703 ();
 sg13g2_decap_4 FILLER_92_734 ();
 sg13g2_fill_2 FILLER_92_738 ();
 sg13g2_decap_4 FILLER_92_772 ();
 sg13g2_fill_2 FILLER_92_786 ();
 sg13g2_decap_4 FILLER_92_801 ();
 sg13g2_fill_1 FILLER_92_805 ();
 sg13g2_fill_2 FILLER_92_823 ();
 sg13g2_fill_2 FILLER_92_846 ();
 sg13g2_fill_1 FILLER_92_848 ();
 sg13g2_fill_1 FILLER_92_853 ();
 sg13g2_fill_2 FILLER_92_862 ();
 sg13g2_decap_8 FILLER_92_923 ();
 sg13g2_decap_4 FILLER_92_930 ();
 sg13g2_decap_8 FILLER_92_938 ();
 sg13g2_decap_8 FILLER_92_945 ();
 sg13g2_decap_8 FILLER_92_952 ();
 sg13g2_decap_8 FILLER_92_999 ();
 sg13g2_fill_2 FILLER_92_1006 ();
 sg13g2_fill_1 FILLER_92_1008 ();
 sg13g2_decap_8 FILLER_92_1013 ();
 sg13g2_decap_8 FILLER_92_1045 ();
 sg13g2_decap_8 FILLER_92_1052 ();
 sg13g2_fill_2 FILLER_92_1059 ();
 sg13g2_decap_4 FILLER_92_1069 ();
 sg13g2_fill_1 FILLER_92_1073 ();
 sg13g2_fill_2 FILLER_92_1094 ();
 sg13g2_fill_2 FILLER_92_1101 ();
 sg13g2_fill_1 FILLER_92_1103 ();
 sg13g2_decap_8 FILLER_92_1116 ();
 sg13g2_decap_8 FILLER_92_1123 ();
 sg13g2_decap_4 FILLER_92_1130 ();
 sg13g2_decap_8 FILLER_92_1149 ();
 sg13g2_decap_8 FILLER_92_1156 ();
 sg13g2_decap_8 FILLER_92_1163 ();
 sg13g2_decap_8 FILLER_92_1170 ();
 sg13g2_decap_8 FILLER_92_1177 ();
 sg13g2_decap_4 FILLER_92_1184 ();
 sg13g2_decap_8 FILLER_92_1196 ();
 sg13g2_decap_8 FILLER_92_1203 ();
 sg13g2_decap_8 FILLER_92_1210 ();
 sg13g2_decap_8 FILLER_92_1217 ();
 sg13g2_fill_2 FILLER_92_1224 ();
 sg13g2_fill_2 FILLER_92_1230 ();
 sg13g2_fill_1 FILLER_92_1232 ();
 sg13g2_decap_8 FILLER_92_1259 ();
 sg13g2_decap_8 FILLER_92_1266 ();
 sg13g2_fill_2 FILLER_92_1273 ();
 sg13g2_fill_1 FILLER_92_1279 ();
 sg13g2_decap_4 FILLER_92_1289 ();
 sg13g2_fill_2 FILLER_92_1293 ();
 sg13g2_decap_8 FILLER_92_1316 ();
 sg13g2_decap_4 FILLER_92_1323 ();
 sg13g2_decap_4 FILLER_92_1336 ();
 sg13g2_decap_4 FILLER_92_1344 ();
 sg13g2_fill_1 FILLER_92_1353 ();
 sg13g2_fill_1 FILLER_92_1358 ();
 sg13g2_decap_8 FILLER_92_1363 ();
 sg13g2_decap_8 FILLER_92_1370 ();
 sg13g2_decap_4 FILLER_92_1377 ();
 sg13g2_fill_2 FILLER_92_1381 ();
 sg13g2_decap_8 FILLER_92_1414 ();
 sg13g2_decap_8 FILLER_92_1421 ();
 sg13g2_decap_8 FILLER_92_1428 ();
 sg13g2_decap_8 FILLER_92_1435 ();
 sg13g2_decap_8 FILLER_92_1442 ();
 sg13g2_fill_1 FILLER_92_1449 ();
 sg13g2_decap_4 FILLER_92_1455 ();
 sg13g2_decap_4 FILLER_92_1463 ();
 sg13g2_decap_4 FILLER_92_1475 ();
 sg13g2_fill_2 FILLER_92_1479 ();
 sg13g2_decap_4 FILLER_92_1510 ();
 sg13g2_fill_2 FILLER_92_1540 ();
 sg13g2_fill_1 FILLER_92_1542 ();
 sg13g2_decap_8 FILLER_92_1578 ();
 sg13g2_fill_1 FILLER_92_1585 ();
 sg13g2_decap_8 FILLER_92_1590 ();
 sg13g2_decap_8 FILLER_92_1597 ();
 sg13g2_decap_8 FILLER_92_1604 ();
 sg13g2_decap_8 FILLER_92_1611 ();
 sg13g2_decap_8 FILLER_92_1618 ();
 sg13g2_decap_8 FILLER_93_0 ();
 sg13g2_decap_8 FILLER_93_7 ();
 sg13g2_decap_8 FILLER_93_14 ();
 sg13g2_decap_8 FILLER_93_21 ();
 sg13g2_decap_8 FILLER_93_28 ();
 sg13g2_decap_8 FILLER_93_35 ();
 sg13g2_decap_8 FILLER_93_42 ();
 sg13g2_decap_8 FILLER_93_49 ();
 sg13g2_decap_4 FILLER_93_56 ();
 sg13g2_decap_8 FILLER_93_64 ();
 sg13g2_fill_1 FILLER_93_71 ();
 sg13g2_decap_4 FILLER_93_97 ();
 sg13g2_fill_1 FILLER_93_101 ();
 sg13g2_decap_8 FILLER_93_131 ();
 sg13g2_decap_8 FILLER_93_150 ();
 sg13g2_fill_1 FILLER_93_157 ();
 sg13g2_fill_1 FILLER_93_165 ();
 sg13g2_decap_8 FILLER_93_191 ();
 sg13g2_fill_2 FILLER_93_198 ();
 sg13g2_decap_4 FILLER_93_204 ();
 sg13g2_fill_2 FILLER_93_208 ();
 sg13g2_decap_4 FILLER_93_227 ();
 sg13g2_fill_2 FILLER_93_231 ();
 sg13g2_fill_1 FILLER_93_246 ();
 sg13g2_fill_2 FILLER_93_253 ();
 sg13g2_fill_1 FILLER_93_255 ();
 sg13g2_decap_8 FILLER_93_297 ();
 sg13g2_decap_8 FILLER_93_304 ();
 sg13g2_decap_8 FILLER_93_311 ();
 sg13g2_fill_2 FILLER_93_318 ();
 sg13g2_fill_1 FILLER_93_320 ();
 sg13g2_decap_8 FILLER_93_325 ();
 sg13g2_fill_2 FILLER_93_332 ();
 sg13g2_fill_1 FILLER_93_334 ();
 sg13g2_fill_2 FILLER_93_361 ();
 sg13g2_decap_8 FILLER_93_367 ();
 sg13g2_decap_4 FILLER_93_374 ();
 sg13g2_decap_4 FILLER_93_420 ();
 sg13g2_fill_2 FILLER_93_424 ();
 sg13g2_fill_2 FILLER_93_459 ();
 sg13g2_fill_1 FILLER_93_461 ();
 sg13g2_fill_2 FILLER_93_488 ();
 sg13g2_decap_8 FILLER_93_499 ();
 sg13g2_decap_4 FILLER_93_506 ();
 sg13g2_fill_1 FILLER_93_510 ();
 sg13g2_fill_1 FILLER_93_515 ();
 sg13g2_fill_1 FILLER_93_521 ();
 sg13g2_fill_1 FILLER_93_527 ();
 sg13g2_fill_2 FILLER_93_532 ();
 sg13g2_fill_2 FILLER_93_539 ();
 sg13g2_decap_4 FILLER_93_551 ();
 sg13g2_fill_1 FILLER_93_555 ();
 sg13g2_fill_1 FILLER_93_568 ();
 sg13g2_fill_2 FILLER_93_574 ();
 sg13g2_decap_8 FILLER_93_590 ();
 sg13g2_decap_4 FILLER_93_597 ();
 sg13g2_fill_2 FILLER_93_615 ();
 sg13g2_fill_1 FILLER_93_617 ();
 sg13g2_fill_1 FILLER_93_626 ();
 sg13g2_decap_8 FILLER_93_634 ();
 sg13g2_decap_8 FILLER_93_641 ();
 sg13g2_decap_4 FILLER_93_648 ();
 sg13g2_fill_2 FILLER_93_652 ();
 sg13g2_decap_4 FILLER_93_667 ();
 sg13g2_decap_8 FILLER_93_679 ();
 sg13g2_fill_2 FILLER_93_686 ();
 sg13g2_fill_1 FILLER_93_688 ();
 sg13g2_decap_8 FILLER_93_698 ();
 sg13g2_decap_4 FILLER_93_705 ();
 sg13g2_fill_2 FILLER_93_709 ();
 sg13g2_decap_8 FILLER_93_715 ();
 sg13g2_decap_8 FILLER_93_722 ();
 sg13g2_decap_8 FILLER_93_729 ();
 sg13g2_decap_8 FILLER_93_736 ();
 sg13g2_decap_8 FILLER_93_743 ();
 sg13g2_decap_8 FILLER_93_750 ();
 sg13g2_decap_8 FILLER_93_757 ();
 sg13g2_decap_8 FILLER_93_764 ();
 sg13g2_fill_2 FILLER_93_771 ();
 sg13g2_fill_1 FILLER_93_773 ();
 sg13g2_decap_8 FILLER_93_785 ();
 sg13g2_decap_4 FILLER_93_792 ();
 sg13g2_decap_8 FILLER_93_801 ();
 sg13g2_decap_4 FILLER_93_808 ();
 sg13g2_fill_2 FILLER_93_812 ();
 sg13g2_decap_4 FILLER_93_819 ();
 sg13g2_decap_8 FILLER_93_828 ();
 sg13g2_fill_2 FILLER_93_841 ();
 sg13g2_fill_1 FILLER_93_843 ();
 sg13g2_decap_8 FILLER_93_848 ();
 sg13g2_decap_4 FILLER_93_855 ();
 sg13g2_fill_1 FILLER_93_859 ();
 sg13g2_decap_8 FILLER_93_872 ();
 sg13g2_fill_2 FILLER_93_879 ();
 sg13g2_fill_1 FILLER_93_881 ();
 sg13g2_decap_8 FILLER_93_887 ();
 sg13g2_decap_8 FILLER_93_894 ();
 sg13g2_decap_8 FILLER_93_901 ();
 sg13g2_fill_1 FILLER_93_920 ();
 sg13g2_fill_1 FILLER_93_968 ();
 sg13g2_decap_4 FILLER_93_976 ();
 sg13g2_fill_1 FILLER_93_980 ();
 sg13g2_fill_2 FILLER_93_985 ();
 sg13g2_fill_1 FILLER_93_987 ();
 sg13g2_fill_1 FILLER_93_997 ();
 sg13g2_decap_8 FILLER_93_1029 ();
 sg13g2_decap_4 FILLER_93_1036 ();
 sg13g2_fill_1 FILLER_93_1040 ();
 sg13g2_fill_2 FILLER_93_1057 ();
 sg13g2_fill_1 FILLER_93_1059 ();
 sg13g2_decap_8 FILLER_93_1064 ();
 sg13g2_decap_8 FILLER_93_1076 ();
 sg13g2_fill_1 FILLER_93_1083 ();
 sg13g2_fill_1 FILLER_93_1088 ();
 sg13g2_fill_2 FILLER_93_1094 ();
 sg13g2_fill_1 FILLER_93_1096 ();
 sg13g2_fill_2 FILLER_93_1102 ();
 sg13g2_fill_1 FILLER_93_1104 ();
 sg13g2_decap_4 FILLER_93_1126 ();
 sg13g2_fill_2 FILLER_93_1147 ();
 sg13g2_fill_1 FILLER_93_1149 ();
 sg13g2_fill_1 FILLER_93_1189 ();
 sg13g2_decap_8 FILLER_93_1207 ();
 sg13g2_fill_2 FILLER_93_1221 ();
 sg13g2_fill_1 FILLER_93_1223 ();
 sg13g2_decap_8 FILLER_93_1250 ();
 sg13g2_decap_8 FILLER_93_1257 ();
 sg13g2_decap_4 FILLER_93_1264 ();
 sg13g2_fill_2 FILLER_93_1294 ();
 sg13g2_decap_8 FILLER_93_1300 ();
 sg13g2_decap_8 FILLER_93_1307 ();
 sg13g2_decap_4 FILLER_93_1314 ();
 sg13g2_fill_1 FILLER_93_1318 ();
 sg13g2_decap_4 FILLER_93_1345 ();
 sg13g2_fill_1 FILLER_93_1349 ();
 sg13g2_decap_8 FILLER_93_1376 ();
 sg13g2_decap_8 FILLER_93_1383 ();
 sg13g2_fill_1 FILLER_93_1437 ();
 sg13g2_decap_8 FILLER_93_1514 ();
 sg13g2_decap_8 FILLER_93_1521 ();
 sg13g2_decap_8 FILLER_93_1528 ();
 sg13g2_fill_2 FILLER_93_1544 ();
 sg13g2_decap_8 FILLER_93_1550 ();
 sg13g2_decap_8 FILLER_93_1557 ();
 sg13g2_decap_4 FILLER_93_1564 ();
 sg13g2_fill_1 FILLER_93_1568 ();
 sg13g2_decap_8 FILLER_93_1604 ();
 sg13g2_decap_8 FILLER_93_1611 ();
 sg13g2_decap_8 FILLER_93_1618 ();
 sg13g2_decap_8 FILLER_94_0 ();
 sg13g2_decap_8 FILLER_94_7 ();
 sg13g2_decap_8 FILLER_94_14 ();
 sg13g2_decap_8 FILLER_94_21 ();
 sg13g2_decap_8 FILLER_94_28 ();
 sg13g2_decap_8 FILLER_94_35 ();
 sg13g2_decap_8 FILLER_94_42 ();
 sg13g2_decap_4 FILLER_94_49 ();
 sg13g2_fill_1 FILLER_94_53 ();
 sg13g2_fill_2 FILLER_94_80 ();
 sg13g2_fill_1 FILLER_94_82 ();
 sg13g2_decap_4 FILLER_94_93 ();
 sg13g2_fill_1 FILLER_94_97 ();
 sg13g2_decap_4 FILLER_94_106 ();
 sg13g2_fill_1 FILLER_94_110 ();
 sg13g2_fill_2 FILLER_94_120 ();
 sg13g2_fill_1 FILLER_94_122 ();
 sg13g2_fill_2 FILLER_94_129 ();
 sg13g2_decap_8 FILLER_94_153 ();
 sg13g2_decap_4 FILLER_94_160 ();
 sg13g2_fill_1 FILLER_94_164 ();
 sg13g2_decap_8 FILLER_94_185 ();
 sg13g2_fill_1 FILLER_94_192 ();
 sg13g2_decap_8 FILLER_94_226 ();
 sg13g2_decap_4 FILLER_94_233 ();
 sg13g2_fill_2 FILLER_94_237 ();
 sg13g2_decap_8 FILLER_94_243 ();
 sg13g2_decap_8 FILLER_94_250 ();
 sg13g2_decap_4 FILLER_94_257 ();
 sg13g2_fill_2 FILLER_94_261 ();
 sg13g2_decap_8 FILLER_94_302 ();
 sg13g2_decap_8 FILLER_94_309 ();
 sg13g2_fill_1 FILLER_94_316 ();
 sg13g2_fill_2 FILLER_94_346 ();
 sg13g2_fill_1 FILLER_94_348 ();
 sg13g2_fill_1 FILLER_94_353 ();
 sg13g2_fill_1 FILLER_94_406 ();
 sg13g2_fill_1 FILLER_94_433 ();
 sg13g2_decap_8 FILLER_94_465 ();
 sg13g2_fill_2 FILLER_94_472 ();
 sg13g2_fill_1 FILLER_94_474 ();
 sg13g2_fill_1 FILLER_94_487 ();
 sg13g2_decap_8 FILLER_94_531 ();
 sg13g2_decap_4 FILLER_94_538 ();
 sg13g2_fill_1 FILLER_94_542 ();
 sg13g2_decap_4 FILLER_94_561 ();
 sg13g2_fill_1 FILLER_94_573 ();
 sg13g2_fill_2 FILLER_94_595 ();
 sg13g2_fill_1 FILLER_94_597 ();
 sg13g2_decap_8 FILLER_94_615 ();
 sg13g2_fill_1 FILLER_94_632 ();
 sg13g2_decap_8 FILLER_94_637 ();
 sg13g2_decap_8 FILLER_94_649 ();
 sg13g2_decap_8 FILLER_94_656 ();
 sg13g2_fill_2 FILLER_94_663 ();
 sg13g2_decap_8 FILLER_94_677 ();
 sg13g2_fill_2 FILLER_94_684 ();
 sg13g2_fill_1 FILLER_94_686 ();
 sg13g2_decap_8 FILLER_94_692 ();
 sg13g2_decap_4 FILLER_94_699 ();
 sg13g2_fill_1 FILLER_94_703 ();
 sg13g2_fill_2 FILLER_94_718 ();
 sg13g2_decap_8 FILLER_94_725 ();
 sg13g2_decap_4 FILLER_94_732 ();
 sg13g2_fill_2 FILLER_94_736 ();
 sg13g2_decap_4 FILLER_94_744 ();
 sg13g2_decap_8 FILLER_94_752 ();
 sg13g2_decap_8 FILLER_94_759 ();
 sg13g2_fill_2 FILLER_94_766 ();
 sg13g2_fill_1 FILLER_94_768 ();
 sg13g2_decap_8 FILLER_94_787 ();
 sg13g2_decap_8 FILLER_94_794 ();
 sg13g2_decap_8 FILLER_94_801 ();
 sg13g2_decap_8 FILLER_94_823 ();
 sg13g2_decap_8 FILLER_94_830 ();
 sg13g2_decap_4 FILLER_94_837 ();
 sg13g2_decap_8 FILLER_94_847 ();
 sg13g2_decap_4 FILLER_94_854 ();
 sg13g2_fill_1 FILLER_94_858 ();
 sg13g2_decap_4 FILLER_94_864 ();
 sg13g2_fill_1 FILLER_94_868 ();
 sg13g2_fill_1 FILLER_94_877 ();
 sg13g2_fill_1 FILLER_94_889 ();
 sg13g2_decap_8 FILLER_94_894 ();
 sg13g2_decap_8 FILLER_94_901 ();
 sg13g2_decap_8 FILLER_94_908 ();
 sg13g2_decap_4 FILLER_94_923 ();
 sg13g2_decap_8 FILLER_94_930 ();
 sg13g2_decap_8 FILLER_94_937 ();
 sg13g2_fill_2 FILLER_94_944 ();
 sg13g2_fill_2 FILLER_94_959 ();
 sg13g2_fill_1 FILLER_94_971 ();
 sg13g2_decap_8 FILLER_94_985 ();
 sg13g2_decap_8 FILLER_94_992 ();
 sg13g2_fill_2 FILLER_94_999 ();
 sg13g2_fill_2 FILLER_94_1006 ();
 sg13g2_fill_1 FILLER_94_1008 ();
 sg13g2_decap_8 FILLER_94_1017 ();
 sg13g2_decap_8 FILLER_94_1024 ();
 sg13g2_fill_1 FILLER_94_1043 ();
 sg13g2_fill_1 FILLER_94_1052 ();
 sg13g2_fill_1 FILLER_94_1068 ();
 sg13g2_decap_8 FILLER_94_1144 ();
 sg13g2_decap_8 FILLER_94_1151 ();
 sg13g2_decap_4 FILLER_94_1162 ();
 sg13g2_fill_2 FILLER_94_1166 ();
 sg13g2_decap_8 FILLER_94_1178 ();
 sg13g2_decap_8 FILLER_94_1185 ();
 sg13g2_decap_8 FILLER_94_1192 ();
 sg13g2_fill_2 FILLER_94_1199 ();
 sg13g2_fill_1 FILLER_94_1201 ();
 sg13g2_decap_8 FILLER_94_1212 ();
 sg13g2_decap_8 FILLER_94_1219 ();
 sg13g2_decap_8 FILLER_94_1226 ();
 sg13g2_decap_8 FILLER_94_1237 ();
 sg13g2_decap_8 FILLER_94_1244 ();
 sg13g2_decap_8 FILLER_94_1251 ();
 sg13g2_fill_1 FILLER_94_1267 ();
 sg13g2_decap_4 FILLER_94_1272 ();
 sg13g2_decap_4 FILLER_94_1279 ();
 sg13g2_decap_8 FILLER_94_1314 ();
 sg13g2_decap_8 FILLER_94_1321 ();
 sg13g2_fill_2 FILLER_94_1328 ();
 sg13g2_fill_1 FILLER_94_1330 ();
 sg13g2_decap_8 FILLER_94_1340 ();
 sg13g2_decap_8 FILLER_94_1347 ();
 sg13g2_decap_8 FILLER_94_1354 ();
 sg13g2_decap_8 FILLER_94_1361 ();
 sg13g2_decap_8 FILLER_94_1368 ();
 sg13g2_decap_8 FILLER_94_1375 ();
 sg13g2_decap_8 FILLER_94_1382 ();
 sg13g2_decap_4 FILLER_94_1389 ();
 sg13g2_fill_2 FILLER_94_1393 ();
 sg13g2_decap_4 FILLER_94_1399 ();
 sg13g2_decap_4 FILLER_94_1408 ();
 sg13g2_fill_1 FILLER_94_1412 ();
 sg13g2_decap_8 FILLER_94_1439 ();
 sg13g2_decap_4 FILLER_94_1446 ();
 sg13g2_fill_2 FILLER_94_1450 ();
 sg13g2_fill_2 FILLER_94_1478 ();
 sg13g2_decap_4 FILLER_94_1532 ();
 sg13g2_fill_2 FILLER_94_1536 ();
 sg13g2_decap_8 FILLER_94_1564 ();
 sg13g2_decap_8 FILLER_94_1571 ();
 sg13g2_fill_2 FILLER_94_1578 ();
 sg13g2_fill_1 FILLER_94_1580 ();
 sg13g2_decap_8 FILLER_94_1610 ();
 sg13g2_decap_8 FILLER_94_1617 ();
 sg13g2_fill_1 FILLER_94_1624 ();
 sg13g2_decap_8 FILLER_95_0 ();
 sg13g2_decap_8 FILLER_95_7 ();
 sg13g2_decap_8 FILLER_95_14 ();
 sg13g2_decap_8 FILLER_95_21 ();
 sg13g2_decap_8 FILLER_95_28 ();
 sg13g2_decap_8 FILLER_95_35 ();
 sg13g2_decap_4 FILLER_95_42 ();
 sg13g2_fill_1 FILLER_95_46 ();
 sg13g2_fill_2 FILLER_95_79 ();
 sg13g2_decap_4 FILLER_95_86 ();
 sg13g2_decap_8 FILLER_95_94 ();
 sg13g2_decap_8 FILLER_95_101 ();
 sg13g2_decap_4 FILLER_95_108 ();
 sg13g2_fill_2 FILLER_95_112 ();
 sg13g2_decap_8 FILLER_95_119 ();
 sg13g2_decap_8 FILLER_95_126 ();
 sg13g2_decap_4 FILLER_95_133 ();
 sg13g2_fill_1 FILLER_95_137 ();
 sg13g2_decap_4 FILLER_95_144 ();
 sg13g2_fill_1 FILLER_95_148 ();
 sg13g2_decap_8 FILLER_95_157 ();
 sg13g2_fill_1 FILLER_95_164 ();
 sg13g2_fill_2 FILLER_95_179 ();
 sg13g2_decap_4 FILLER_95_189 ();
 sg13g2_fill_1 FILLER_95_193 ();
 sg13g2_decap_8 FILLER_95_224 ();
 sg13g2_decap_8 FILLER_95_231 ();
 sg13g2_decap_4 FILLER_95_238 ();
 sg13g2_fill_2 FILLER_95_242 ();
 sg13g2_fill_1 FILLER_95_252 ();
 sg13g2_fill_2 FILLER_95_261 ();
 sg13g2_fill_1 FILLER_95_276 ();
 sg13g2_decap_8 FILLER_95_282 ();
 sg13g2_decap_8 FILLER_95_289 ();
 sg13g2_decap_8 FILLER_95_296 ();
 sg13g2_decap_4 FILLER_95_303 ();
 sg13g2_fill_2 FILLER_95_307 ();
 sg13g2_decap_4 FILLER_95_340 ();
 sg13g2_fill_1 FILLER_95_348 ();
 sg13g2_fill_1 FILLER_95_382 ();
 sg13g2_decap_8 FILLER_95_397 ();
 sg13g2_decap_4 FILLER_95_404 ();
 sg13g2_fill_1 FILLER_95_408 ();
 sg13g2_decap_4 FILLER_95_413 ();
 sg13g2_fill_1 FILLER_95_447 ();
 sg13g2_decap_4 FILLER_95_533 ();
 sg13g2_decap_8 FILLER_95_542 ();
 sg13g2_fill_1 FILLER_95_549 ();
 sg13g2_fill_2 FILLER_95_566 ();
 sg13g2_fill_1 FILLER_95_568 ();
 sg13g2_decap_4 FILLER_95_583 ();
 sg13g2_fill_1 FILLER_95_587 ();
 sg13g2_decap_8 FILLER_95_606 ();
 sg13g2_decap_8 FILLER_95_613 ();
 sg13g2_fill_1 FILLER_95_620 ();
 sg13g2_decap_4 FILLER_95_636 ();
 sg13g2_fill_2 FILLER_95_653 ();
 sg13g2_fill_1 FILLER_95_655 ();
 sg13g2_fill_1 FILLER_95_662 ();
 sg13g2_decap_8 FILLER_95_671 ();
 sg13g2_decap_8 FILLER_95_678 ();
 sg13g2_fill_1 FILLER_95_685 ();
 sg13g2_decap_4 FILLER_95_694 ();
 sg13g2_fill_1 FILLER_95_714 ();
 sg13g2_fill_1 FILLER_95_721 ();
 sg13g2_fill_1 FILLER_95_728 ();
 sg13g2_fill_1 FILLER_95_735 ();
 sg13g2_fill_1 FILLER_95_740 ();
 sg13g2_decap_8 FILLER_95_767 ();
 sg13g2_fill_2 FILLER_95_774 ();
 sg13g2_fill_2 FILLER_95_789 ();
 sg13g2_decap_4 FILLER_95_804 ();
 sg13g2_fill_2 FILLER_95_808 ();
 sg13g2_fill_2 FILLER_95_822 ();
 sg13g2_fill_2 FILLER_95_828 ();
 sg13g2_fill_1 FILLER_95_836 ();
 sg13g2_fill_1 FILLER_95_846 ();
 sg13g2_fill_1 FILLER_95_852 ();
 sg13g2_decap_4 FILLER_95_858 ();
 sg13g2_fill_2 FILLER_95_884 ();
 sg13g2_fill_1 FILLER_95_886 ();
 sg13g2_decap_8 FILLER_95_914 ();
 sg13g2_decap_4 FILLER_95_921 ();
 sg13g2_fill_1 FILLER_95_925 ();
 sg13g2_decap_4 FILLER_95_935 ();
 sg13g2_fill_2 FILLER_95_939 ();
 sg13g2_fill_2 FILLER_95_972 ();
 sg13g2_fill_1 FILLER_95_974 ();
 sg13g2_decap_4 FILLER_95_987 ();
 sg13g2_decap_8 FILLER_95_1004 ();
 sg13g2_decap_8 FILLER_95_1011 ();
 sg13g2_decap_8 FILLER_95_1018 ();
 sg13g2_decap_8 FILLER_95_1025 ();
 sg13g2_decap_8 FILLER_95_1032 ();
 sg13g2_fill_2 FILLER_95_1039 ();
 sg13g2_fill_1 FILLER_95_1041 ();
 sg13g2_decap_8 FILLER_95_1053 ();
 sg13g2_decap_8 FILLER_95_1060 ();
 sg13g2_decap_4 FILLER_95_1067 ();
 sg13g2_decap_8 FILLER_95_1076 ();
 sg13g2_fill_2 FILLER_95_1083 ();
 sg13g2_fill_2 FILLER_95_1103 ();
 sg13g2_fill_1 FILLER_95_1105 ();
 sg13g2_fill_1 FILLER_95_1115 ();
 sg13g2_fill_1 FILLER_95_1124 ();
 sg13g2_fill_2 FILLER_95_1133 ();
 sg13g2_fill_1 FILLER_95_1135 ();
 sg13g2_decap_4 FILLER_95_1192 ();
 sg13g2_decap_4 FILLER_95_1206 ();
 sg13g2_decap_8 FILLER_95_1231 ();
 sg13g2_decap_8 FILLER_95_1238 ();
 sg13g2_decap_8 FILLER_95_1245 ();
 sg13g2_fill_2 FILLER_95_1252 ();
 sg13g2_fill_1 FILLER_95_1254 ();
 sg13g2_fill_2 FILLER_95_1306 ();
 sg13g2_decap_8 FILLER_95_1312 ();
 sg13g2_fill_2 FILLER_95_1319 ();
 sg13g2_fill_1 FILLER_95_1350 ();
 sg13g2_decap_8 FILLER_95_1372 ();
 sg13g2_fill_2 FILLER_95_1379 ();
 sg13g2_fill_1 FILLER_95_1381 ();
 sg13g2_fill_2 FILLER_95_1392 ();
 sg13g2_fill_1 FILLER_95_1402 ();
 sg13g2_fill_2 FILLER_95_1407 ();
 sg13g2_fill_1 FILLER_95_1414 ();
 sg13g2_fill_2 FILLER_95_1470 ();
 sg13g2_fill_1 FILLER_95_1472 ();
 sg13g2_fill_2 FILLER_95_1510 ();
 sg13g2_fill_1 FILLER_95_1512 ();
 sg13g2_decap_4 FILLER_95_1521 ();
 sg13g2_fill_1 FILLER_95_1525 ();
 sg13g2_decap_8 FILLER_95_1530 ();
 sg13g2_decap_8 FILLER_95_1537 ();
 sg13g2_decap_8 FILLER_95_1544 ();
 sg13g2_decap_8 FILLER_95_1551 ();
 sg13g2_decap_8 FILLER_95_1558 ();
 sg13g2_decap_8 FILLER_95_1565 ();
 sg13g2_decap_8 FILLER_95_1572 ();
 sg13g2_decap_8 FILLER_95_1608 ();
 sg13g2_decap_8 FILLER_95_1615 ();
 sg13g2_fill_2 FILLER_95_1622 ();
 sg13g2_fill_1 FILLER_95_1624 ();
 sg13g2_decap_8 FILLER_96_0 ();
 sg13g2_decap_8 FILLER_96_7 ();
 sg13g2_decap_8 FILLER_96_14 ();
 sg13g2_decap_8 FILLER_96_21 ();
 sg13g2_decap_8 FILLER_96_28 ();
 sg13g2_decap_8 FILLER_96_35 ();
 sg13g2_fill_2 FILLER_96_42 ();
 sg13g2_decap_8 FILLER_96_70 ();
 sg13g2_fill_1 FILLER_96_77 ();
 sg13g2_fill_2 FILLER_96_132 ();
 sg13g2_decap_4 FILLER_96_154 ();
 sg13g2_decap_8 FILLER_96_162 ();
 sg13g2_decap_4 FILLER_96_169 ();
 sg13g2_fill_1 FILLER_96_173 ();
 sg13g2_decap_8 FILLER_96_179 ();
 sg13g2_fill_2 FILLER_96_186 ();
 sg13g2_decap_8 FILLER_96_202 ();
 sg13g2_fill_1 FILLER_96_209 ();
 sg13g2_decap_4 FILLER_96_236 ();
 sg13g2_fill_1 FILLER_96_240 ();
 sg13g2_decap_4 FILLER_96_255 ();
 sg13g2_fill_1 FILLER_96_259 ();
 sg13g2_fill_2 FILLER_96_284 ();
 sg13g2_fill_1 FILLER_96_286 ();
 sg13g2_fill_2 FILLER_96_292 ();
 sg13g2_fill_1 FILLER_96_302 ();
 sg13g2_fill_2 FILLER_96_313 ();
 sg13g2_decap_8 FILLER_96_319 ();
 sg13g2_decap_8 FILLER_96_326 ();
 sg13g2_fill_2 FILLER_96_333 ();
 sg13g2_fill_1 FILLER_96_335 ();
 sg13g2_fill_2 FILLER_96_367 ();
 sg13g2_fill_1 FILLER_96_369 ();
 sg13g2_decap_4 FILLER_96_395 ();
 sg13g2_fill_1 FILLER_96_399 ();
 sg13g2_decap_8 FILLER_96_404 ();
 sg13g2_decap_8 FILLER_96_411 ();
 sg13g2_decap_8 FILLER_96_452 ();
 sg13g2_decap_8 FILLER_96_459 ();
 sg13g2_decap_8 FILLER_96_466 ();
 sg13g2_decap_4 FILLER_96_473 ();
 sg13g2_fill_1 FILLER_96_477 ();
 sg13g2_fill_1 FILLER_96_504 ();
 sg13g2_fill_2 FILLER_96_531 ();
 sg13g2_fill_2 FILLER_96_537 ();
 sg13g2_fill_2 FILLER_96_544 ();
 sg13g2_fill_1 FILLER_96_558 ();
 sg13g2_fill_2 FILLER_96_564 ();
 sg13g2_fill_1 FILLER_96_566 ();
 sg13g2_fill_2 FILLER_96_572 ();
 sg13g2_fill_1 FILLER_96_574 ();
 sg13g2_decap_8 FILLER_96_583 ();
 sg13g2_decap_8 FILLER_96_590 ();
 sg13g2_fill_2 FILLER_96_597 ();
 sg13g2_decap_4 FILLER_96_604 ();
 sg13g2_fill_2 FILLER_96_608 ();
 sg13g2_decap_8 FILLER_96_614 ();
 sg13g2_decap_8 FILLER_96_621 ();
 sg13g2_decap_4 FILLER_96_628 ();
 sg13g2_decap_4 FILLER_96_640 ();
 sg13g2_fill_1 FILLER_96_644 ();
 sg13g2_decap_8 FILLER_96_653 ();
 sg13g2_decap_8 FILLER_96_660 ();
 sg13g2_decap_8 FILLER_96_667 ();
 sg13g2_decap_8 FILLER_96_674 ();
 sg13g2_decap_8 FILLER_96_681 ();
 sg13g2_decap_4 FILLER_96_688 ();
 sg13g2_fill_1 FILLER_96_692 ();
 sg13g2_decap_4 FILLER_96_706 ();
 sg13g2_fill_1 FILLER_96_713 ();
 sg13g2_decap_8 FILLER_96_719 ();
 sg13g2_decap_8 FILLER_96_726 ();
 sg13g2_decap_8 FILLER_96_738 ();
 sg13g2_decap_8 FILLER_96_745 ();
 sg13g2_decap_8 FILLER_96_752 ();
 sg13g2_decap_8 FILLER_96_759 ();
 sg13g2_decap_8 FILLER_96_766 ();
 sg13g2_fill_1 FILLER_96_773 ();
 sg13g2_decap_8 FILLER_96_780 ();
 sg13g2_decap_8 FILLER_96_787 ();
 sg13g2_fill_1 FILLER_96_794 ();
 sg13g2_decap_4 FILLER_96_800 ();
 sg13g2_fill_1 FILLER_96_804 ();
 sg13g2_decap_8 FILLER_96_842 ();
 sg13g2_fill_1 FILLER_96_849 ();
 sg13g2_fill_1 FILLER_96_865 ();
 sg13g2_decap_4 FILLER_96_877 ();
 sg13g2_decap_8 FILLER_96_897 ();
 sg13g2_fill_1 FILLER_96_904 ();
 sg13g2_decap_8 FILLER_96_909 ();
 sg13g2_decap_4 FILLER_96_916 ();
 sg13g2_fill_1 FILLER_96_920 ();
 sg13g2_decap_8 FILLER_96_930 ();
 sg13g2_decap_8 FILLER_96_937 ();
 sg13g2_decap_4 FILLER_96_944 ();
 sg13g2_fill_1 FILLER_96_948 ();
 sg13g2_fill_2 FILLER_96_966 ();
 sg13g2_decap_8 FILLER_96_981 ();
 sg13g2_decap_8 FILLER_96_988 ();
 sg13g2_fill_2 FILLER_96_995 ();
 sg13g2_fill_1 FILLER_96_997 ();
 sg13g2_decap_4 FILLER_96_1012 ();
 sg13g2_fill_2 FILLER_96_1027 ();
 sg13g2_fill_1 FILLER_96_1033 ();
 sg13g2_decap_8 FILLER_96_1042 ();
 sg13g2_decap_8 FILLER_96_1049 ();
 sg13g2_decap_4 FILLER_96_1061 ();
 sg13g2_fill_2 FILLER_96_1065 ();
 sg13g2_decap_8 FILLER_96_1074 ();
 sg13g2_fill_2 FILLER_96_1081 ();
 sg13g2_fill_1 FILLER_96_1083 ();
 sg13g2_decap_4 FILLER_96_1099 ();
 sg13g2_fill_1 FILLER_96_1103 ();
 sg13g2_fill_1 FILLER_96_1173 ();
 sg13g2_decap_4 FILLER_96_1184 ();
 sg13g2_fill_2 FILLER_96_1188 ();
 sg13g2_fill_1 FILLER_96_1195 ();
 sg13g2_decap_8 FILLER_96_1209 ();
 sg13g2_decap_4 FILLER_96_1216 ();
 sg13g2_fill_1 FILLER_96_1220 ();
 sg13g2_decap_4 FILLER_96_1229 ();
 sg13g2_fill_2 FILLER_96_1233 ();
 sg13g2_decap_8 FILLER_96_1240 ();
 sg13g2_decap_8 FILLER_96_1247 ();
 sg13g2_decap_4 FILLER_96_1254 ();
 sg13g2_fill_2 FILLER_96_1263 ();
 sg13g2_fill_1 FILLER_96_1265 ();
 sg13g2_fill_2 FILLER_96_1271 ();
 sg13g2_fill_1 FILLER_96_1273 ();
 sg13g2_decap_4 FILLER_96_1278 ();
 sg13g2_fill_1 FILLER_96_1282 ();
 sg13g2_decap_4 FILLER_96_1288 ();
 sg13g2_fill_1 FILLER_96_1292 ();
 sg13g2_decap_8 FILLER_96_1374 ();
 sg13g2_fill_1 FILLER_96_1381 ();
 sg13g2_decap_8 FILLER_96_1411 ();
 sg13g2_decap_4 FILLER_96_1418 ();
 sg13g2_decap_8 FILLER_96_1426 ();
 sg13g2_decap_4 FILLER_96_1433 ();
 sg13g2_fill_1 FILLER_96_1437 ();
 sg13g2_decap_8 FILLER_96_1541 ();
 sg13g2_decap_8 FILLER_96_1548 ();
 sg13g2_decap_8 FILLER_96_1555 ();
 sg13g2_decap_8 FILLER_96_1562 ();
 sg13g2_decap_8 FILLER_96_1569 ();
 sg13g2_decap_8 FILLER_96_1576 ();
 sg13g2_decap_8 FILLER_96_1583 ();
 sg13g2_decap_8 FILLER_96_1590 ();
 sg13g2_decap_8 FILLER_96_1597 ();
 sg13g2_decap_8 FILLER_96_1604 ();
 sg13g2_decap_8 FILLER_96_1611 ();
 sg13g2_decap_8 FILLER_96_1618 ();
 sg13g2_decap_8 FILLER_97_0 ();
 sg13g2_decap_8 FILLER_97_7 ();
 sg13g2_decap_8 FILLER_97_14 ();
 sg13g2_decap_8 FILLER_97_21 ();
 sg13g2_decap_4 FILLER_97_28 ();
 sg13g2_decap_8 FILLER_97_36 ();
 sg13g2_decap_4 FILLER_97_43 ();
 sg13g2_decap_4 FILLER_97_51 ();
 sg13g2_decap_8 FILLER_97_59 ();
 sg13g2_decap_8 FILLER_97_66 ();
 sg13g2_decap_8 FILLER_97_77 ();
 sg13g2_decap_8 FILLER_97_84 ();
 sg13g2_decap_8 FILLER_97_91 ();
 sg13g2_decap_8 FILLER_97_98 ();
 sg13g2_decap_8 FILLER_97_105 ();
 sg13g2_fill_1 FILLER_97_112 ();
 sg13g2_decap_8 FILLER_97_121 ();
 sg13g2_decap_4 FILLER_97_128 ();
 sg13g2_fill_1 FILLER_97_140 ();
 sg13g2_decap_4 FILLER_97_147 ();
 sg13g2_decap_4 FILLER_97_177 ();
 sg13g2_decap_4 FILLER_97_185 ();
 sg13g2_fill_2 FILLER_97_189 ();
 sg13g2_decap_8 FILLER_97_199 ();
 sg13g2_decap_4 FILLER_97_206 ();
 sg13g2_fill_1 FILLER_97_222 ();
 sg13g2_fill_2 FILLER_97_227 ();
 sg13g2_fill_1 FILLER_97_234 ();
 sg13g2_fill_2 FILLER_97_240 ();
 sg13g2_fill_2 FILLER_97_259 ();
 sg13g2_decap_8 FILLER_97_269 ();
 sg13g2_decap_4 FILLER_97_276 ();
 sg13g2_fill_1 FILLER_97_280 ();
 sg13g2_decap_4 FILLER_97_286 ();
 sg13g2_fill_2 FILLER_97_290 ();
 sg13g2_fill_2 FILLER_97_333 ();
 sg13g2_decap_8 FILLER_97_340 ();
 sg13g2_decap_8 FILLER_97_347 ();
 sg13g2_decap_8 FILLER_97_354 ();
 sg13g2_fill_1 FILLER_97_361 ();
 sg13g2_decap_4 FILLER_97_388 ();
 sg13g2_fill_1 FILLER_97_392 ();
 sg13g2_decap_8 FILLER_97_423 ();
 sg13g2_fill_1 FILLER_97_430 ();
 sg13g2_decap_8 FILLER_97_435 ();
 sg13g2_fill_1 FILLER_97_442 ();
 sg13g2_fill_2 FILLER_97_451 ();
 sg13g2_decap_8 FILLER_97_458 ();
 sg13g2_decap_4 FILLER_97_465 ();
 sg13g2_decap_8 FILLER_97_473 ();
 sg13g2_decap_8 FILLER_97_522 ();
 sg13g2_decap_8 FILLER_97_529 ();
 sg13g2_decap_8 FILLER_97_536 ();
 sg13g2_decap_8 FILLER_97_543 ();
 sg13g2_decap_8 FILLER_97_550 ();
 sg13g2_decap_4 FILLER_97_557 ();
 sg13g2_decap_8 FILLER_97_566 ();
 sg13g2_decap_4 FILLER_97_573 ();
 sg13g2_fill_2 FILLER_97_577 ();
 sg13g2_decap_8 FILLER_97_589 ();
 sg13g2_decap_4 FILLER_97_596 ();
 sg13g2_decap_4 FILLER_97_604 ();
 sg13g2_fill_2 FILLER_97_608 ();
 sg13g2_fill_1 FILLER_97_615 ();
 sg13g2_fill_1 FILLER_97_621 ();
 sg13g2_decap_8 FILLER_97_632 ();
 sg13g2_fill_2 FILLER_97_639 ();
 sg13g2_decap_8 FILLER_97_652 ();
 sg13g2_decap_4 FILLER_97_659 ();
 sg13g2_fill_1 FILLER_97_663 ();
 sg13g2_decap_8 FILLER_97_669 ();
 sg13g2_decap_8 FILLER_97_676 ();
 sg13g2_fill_2 FILLER_97_683 ();
 sg13g2_fill_1 FILLER_97_685 ();
 sg13g2_fill_2 FILLER_97_693 ();
 sg13g2_fill_2 FILLER_97_701 ();
 sg13g2_fill_1 FILLER_97_707 ();
 sg13g2_fill_2 FILLER_97_721 ();
 sg13g2_fill_1 FILLER_97_723 ();
 sg13g2_fill_1 FILLER_97_729 ();
 sg13g2_fill_2 FILLER_97_735 ();
 sg13g2_fill_1 FILLER_97_747 ();
 sg13g2_decap_4 FILLER_97_758 ();
 sg13g2_fill_1 FILLER_97_762 ();
 sg13g2_decap_8 FILLER_97_768 ();
 sg13g2_decap_4 FILLER_97_775 ();
 sg13g2_fill_2 FILLER_97_790 ();
 sg13g2_decap_8 FILLER_97_798 ();
 sg13g2_decap_8 FILLER_97_805 ();
 sg13g2_decap_4 FILLER_97_812 ();
 sg13g2_fill_1 FILLER_97_816 ();
 sg13g2_decap_8 FILLER_97_822 ();
 sg13g2_decap_4 FILLER_97_829 ();
 sg13g2_fill_2 FILLER_97_833 ();
 sg13g2_decap_8 FILLER_97_840 ();
 sg13g2_decap_8 FILLER_97_847 ();
 sg13g2_decap_4 FILLER_97_854 ();
 sg13g2_decap_4 FILLER_97_866 ();
 sg13g2_fill_1 FILLER_97_870 ();
 sg13g2_decap_8 FILLER_97_891 ();
 sg13g2_fill_2 FILLER_97_898 ();
 sg13g2_fill_1 FILLER_97_912 ();
 sg13g2_decap_8 FILLER_97_917 ();
 sg13g2_decap_8 FILLER_97_924 ();
 sg13g2_decap_8 FILLER_97_931 ();
 sg13g2_fill_2 FILLER_97_938 ();
 sg13g2_fill_1 FILLER_97_940 ();
 sg13g2_decap_8 FILLER_97_967 ();
 sg13g2_decap_8 FILLER_97_974 ();
 sg13g2_decap_8 FILLER_97_981 ();
 sg13g2_decap_4 FILLER_97_988 ();
 sg13g2_fill_1 FILLER_97_992 ();
 sg13g2_fill_1 FILLER_97_1032 ();
 sg13g2_fill_1 FILLER_97_1038 ();
 sg13g2_fill_2 FILLER_97_1064 ();
 sg13g2_fill_1 FILLER_97_1066 ();
 sg13g2_decap_8 FILLER_97_1074 ();
 sg13g2_decap_4 FILLER_97_1081 ();
 sg13g2_fill_2 FILLER_97_1085 ();
 sg13g2_fill_2 FILLER_97_1122 ();
 sg13g2_decap_8 FILLER_97_1176 ();
 sg13g2_decap_4 FILLER_97_1183 ();
 sg13g2_fill_2 FILLER_97_1187 ();
 sg13g2_fill_2 FILLER_97_1194 ();
 sg13g2_fill_2 FILLER_97_1202 ();
 sg13g2_fill_2 FILLER_97_1227 ();
 sg13g2_decap_8 FILLER_97_1246 ();
 sg13g2_decap_8 FILLER_97_1253 ();
 sg13g2_decap_8 FILLER_97_1312 ();
 sg13g2_decap_4 FILLER_97_1319 ();
 sg13g2_decap_8 FILLER_97_1327 ();
 sg13g2_fill_1 FILLER_97_1334 ();
 sg13g2_fill_1 FILLER_97_1340 ();
 sg13g2_fill_2 FILLER_97_1346 ();
 sg13g2_fill_1 FILLER_97_1348 ();
 sg13g2_fill_1 FILLER_97_1375 ();
 sg13g2_decap_8 FILLER_97_1410 ();
 sg13g2_decap_8 FILLER_97_1417 ();
 sg13g2_fill_2 FILLER_97_1424 ();
 sg13g2_fill_2 FILLER_97_1472 ();
 sg13g2_fill_2 FILLER_97_1489 ();
 sg13g2_decap_8 FILLER_97_1543 ();
 sg13g2_decap_8 FILLER_97_1550 ();
 sg13g2_decap_8 FILLER_97_1557 ();
 sg13g2_decap_8 FILLER_97_1564 ();
 sg13g2_decap_8 FILLER_97_1571 ();
 sg13g2_decap_8 FILLER_97_1578 ();
 sg13g2_decap_8 FILLER_97_1585 ();
 sg13g2_decap_8 FILLER_97_1592 ();
 sg13g2_decap_8 FILLER_97_1599 ();
 sg13g2_decap_8 FILLER_97_1606 ();
 sg13g2_decap_8 FILLER_97_1613 ();
 sg13g2_decap_4 FILLER_97_1620 ();
 sg13g2_fill_1 FILLER_97_1624 ();
 sg13g2_decap_8 FILLER_98_0 ();
 sg13g2_decap_8 FILLER_98_7 ();
 sg13g2_decap_8 FILLER_98_14 ();
 sg13g2_decap_4 FILLER_98_21 ();
 sg13g2_fill_1 FILLER_98_25 ();
 sg13g2_decap_8 FILLER_98_60 ();
 sg13g2_fill_2 FILLER_98_93 ();
 sg13g2_fill_1 FILLER_98_95 ();
 sg13g2_decap_8 FILLER_98_100 ();
 sg13g2_decap_8 FILLER_98_107 ();
 sg13g2_decap_8 FILLER_98_114 ();
 sg13g2_decap_8 FILLER_98_121 ();
 sg13g2_decap_4 FILLER_98_128 ();
 sg13g2_decap_4 FILLER_98_136 ();
 sg13g2_fill_1 FILLER_98_140 ();
 sg13g2_decap_4 FILLER_98_146 ();
 sg13g2_fill_1 FILLER_98_150 ();
 sg13g2_decap_8 FILLER_98_161 ();
 sg13g2_decap_8 FILLER_98_199 ();
 sg13g2_decap_8 FILLER_98_206 ();
 sg13g2_decap_8 FILLER_98_213 ();
 sg13g2_decap_8 FILLER_98_220 ();
 sg13g2_decap_8 FILLER_98_227 ();
 sg13g2_decap_4 FILLER_98_234 ();
 sg13g2_fill_2 FILLER_98_238 ();
 sg13g2_fill_2 FILLER_98_245 ();
 sg13g2_decap_8 FILLER_98_269 ();
 sg13g2_decap_8 FILLER_98_276 ();
 sg13g2_decap_8 FILLER_98_283 ();
 sg13g2_decap_8 FILLER_98_290 ();
 sg13g2_decap_8 FILLER_98_297 ();
 sg13g2_decap_8 FILLER_98_304 ();
 sg13g2_decap_8 FILLER_98_311 ();
 sg13g2_decap_8 FILLER_98_318 ();
 sg13g2_decap_8 FILLER_98_335 ();
 sg13g2_fill_1 FILLER_98_342 ();
 sg13g2_decap_4 FILLER_98_348 ();
 sg13g2_fill_1 FILLER_98_352 ();
 sg13g2_decap_8 FILLER_98_357 ();
 sg13g2_decap_4 FILLER_98_364 ();
 sg13g2_fill_2 FILLER_98_368 ();
 sg13g2_decap_4 FILLER_98_374 ();
 sg13g2_decap_8 FILLER_98_388 ();
 sg13g2_decap_4 FILLER_98_395 ();
 sg13g2_fill_1 FILLER_98_409 ();
 sg13g2_fill_2 FILLER_98_436 ();
 sg13g2_fill_2 FILLER_98_493 ();
 sg13g2_fill_2 FILLER_98_524 ();
 sg13g2_fill_1 FILLER_98_526 ();
 sg13g2_decap_4 FILLER_98_537 ();
 sg13g2_fill_2 FILLER_98_550 ();
 sg13g2_fill_1 FILLER_98_552 ();
 sg13g2_fill_2 FILLER_98_577 ();
 sg13g2_decap_8 FILLER_98_589 ();
 sg13g2_decap_4 FILLER_98_596 ();
 sg13g2_fill_2 FILLER_98_617 ();
 sg13g2_fill_1 FILLER_98_619 ();
 sg13g2_fill_2 FILLER_98_633 ();
 sg13g2_fill_1 FILLER_98_646 ();
 sg13g2_fill_2 FILLER_98_652 ();
 sg13g2_decap_8 FILLER_98_659 ();
 sg13g2_decap_8 FILLER_98_666 ();
 sg13g2_fill_2 FILLER_98_673 ();
 sg13g2_decap_8 FILLER_98_689 ();
 sg13g2_fill_1 FILLER_98_696 ();
 sg13g2_decap_8 FILLER_98_703 ();
 sg13g2_decap_4 FILLER_98_716 ();
 sg13g2_fill_1 FILLER_98_720 ();
 sg13g2_decap_4 FILLER_98_735 ();
 sg13g2_fill_1 FILLER_98_765 ();
 sg13g2_fill_1 FILLER_98_772 ();
 sg13g2_fill_1 FILLER_98_778 ();
 sg13g2_fill_1 FILLER_98_789 ();
 sg13g2_fill_2 FILLER_98_795 ();
 sg13g2_fill_2 FILLER_98_802 ();
 sg13g2_fill_1 FILLER_98_809 ();
 sg13g2_fill_2 FILLER_98_825 ();
 sg13g2_fill_2 FILLER_98_834 ();
 sg13g2_decap_8 FILLER_98_840 ();
 sg13g2_decap_4 FILLER_98_847 ();
 sg13g2_fill_2 FILLER_98_851 ();
 sg13g2_decap_8 FILLER_98_880 ();
 sg13g2_decap_8 FILLER_98_887 ();
 sg13g2_fill_2 FILLER_98_894 ();
 sg13g2_fill_1 FILLER_98_896 ();
 sg13g2_decap_8 FILLER_98_902 ();
 sg13g2_decap_4 FILLER_98_909 ();
 sg13g2_fill_2 FILLER_98_913 ();
 sg13g2_fill_2 FILLER_98_938 ();
 sg13g2_fill_1 FILLER_98_940 ();
 sg13g2_decap_4 FILLER_98_954 ();
 sg13g2_fill_2 FILLER_98_958 ();
 sg13g2_fill_2 FILLER_98_965 ();
 sg13g2_fill_2 FILLER_98_976 ();
 sg13g2_fill_1 FILLER_98_991 ();
 sg13g2_decap_8 FILLER_98_1001 ();
 sg13g2_fill_1 FILLER_98_1008 ();
 sg13g2_fill_1 FILLER_98_1024 ();
 sg13g2_decap_8 FILLER_98_1033 ();
 sg13g2_fill_2 FILLER_98_1040 ();
 sg13g2_fill_1 FILLER_98_1042 ();
 sg13g2_fill_2 FILLER_98_1048 ();
 sg13g2_decap_8 FILLER_98_1058 ();
 sg13g2_decap_4 FILLER_98_1071 ();
 sg13g2_fill_1 FILLER_98_1091 ();
 sg13g2_fill_1 FILLER_98_1104 ();
 sg13g2_fill_2 FILLER_98_1136 ();
 sg13g2_fill_1 FILLER_98_1138 ();
 sg13g2_fill_1 FILLER_98_1171 ();
 sg13g2_fill_2 FILLER_98_1177 ();
 sg13g2_decap_4 FILLER_98_1182 ();
 sg13g2_decap_8 FILLER_98_1199 ();
 sg13g2_fill_1 FILLER_98_1206 ();
 sg13g2_fill_1 FILLER_98_1211 ();
 sg13g2_fill_2 FILLER_98_1217 ();
 sg13g2_decap_8 FILLER_98_1224 ();
 sg13g2_decap_8 FILLER_98_1231 ();
 sg13g2_decap_8 FILLER_98_1238 ();
 sg13g2_decap_8 FILLER_98_1245 ();
 sg13g2_decap_8 FILLER_98_1252 ();
 sg13g2_decap_8 FILLER_98_1259 ();
 sg13g2_fill_1 FILLER_98_1266 ();
 sg13g2_decap_4 FILLER_98_1271 ();
 sg13g2_decap_8 FILLER_98_1307 ();
 sg13g2_fill_2 FILLER_98_1314 ();
 sg13g2_decap_4 FILLER_98_1342 ();
 sg13g2_decap_4 FILLER_98_1350 ();
 sg13g2_decap_8 FILLER_98_1358 ();
 sg13g2_decap_8 FILLER_98_1365 ();
 sg13g2_fill_2 FILLER_98_1372 ();
 sg13g2_fill_1 FILLER_98_1374 ();
 sg13g2_decap_4 FILLER_98_1401 ();
 sg13g2_fill_2 FILLER_98_1405 ();
 sg13g2_decap_4 FILLER_98_1420 ();
 sg13g2_fill_2 FILLER_98_1424 ();
 sg13g2_fill_1 FILLER_98_1431 ();
 sg13g2_fill_1 FILLER_98_1457 ();
 sg13g2_decap_8 FILLER_98_1512 ();
 sg13g2_decap_8 FILLER_98_1519 ();
 sg13g2_decap_8 FILLER_98_1526 ();
 sg13g2_decap_8 FILLER_98_1533 ();
 sg13g2_decap_8 FILLER_98_1540 ();
 sg13g2_decap_8 FILLER_98_1547 ();
 sg13g2_decap_8 FILLER_98_1554 ();
 sg13g2_decap_8 FILLER_98_1561 ();
 sg13g2_decap_8 FILLER_98_1568 ();
 sg13g2_decap_8 FILLER_98_1575 ();
 sg13g2_decap_8 FILLER_98_1582 ();
 sg13g2_decap_8 FILLER_98_1589 ();
 sg13g2_decap_8 FILLER_98_1596 ();
 sg13g2_decap_8 FILLER_98_1603 ();
 sg13g2_decap_8 FILLER_98_1610 ();
 sg13g2_decap_8 FILLER_98_1617 ();
 sg13g2_fill_1 FILLER_98_1624 ();
 sg13g2_decap_8 FILLER_99_0 ();
 sg13g2_decap_8 FILLER_99_7 ();
 sg13g2_decap_8 FILLER_99_14 ();
 sg13g2_decap_8 FILLER_99_21 ();
 sg13g2_decap_8 FILLER_99_28 ();
 sg13g2_decap_4 FILLER_99_35 ();
 sg13g2_fill_2 FILLER_99_39 ();
 sg13g2_decap_8 FILLER_99_53 ();
 sg13g2_fill_1 FILLER_99_60 ();
 sg13g2_fill_2 FILLER_99_69 ();
 sg13g2_fill_1 FILLER_99_78 ();
 sg13g2_decap_4 FILLER_99_108 ();
 sg13g2_decap_8 FILLER_99_157 ();
 sg13g2_fill_2 FILLER_99_164 ();
 sg13g2_fill_1 FILLER_99_166 ();
 sg13g2_fill_1 FILLER_99_177 ();
 sg13g2_decap_8 FILLER_99_219 ();
 sg13g2_decap_4 FILLER_99_226 ();
 sg13g2_decap_8 FILLER_99_234 ();
 sg13g2_decap_8 FILLER_99_241 ();
 sg13g2_decap_8 FILLER_99_248 ();
 sg13g2_decap_4 FILLER_99_255 ();
 sg13g2_fill_2 FILLER_99_259 ();
 sg13g2_decap_8 FILLER_99_269 ();
 sg13g2_decap_8 FILLER_99_276 ();
 sg13g2_decap_4 FILLER_99_319 ();
 sg13g2_fill_2 FILLER_99_323 ();
 sg13g2_decap_4 FILLER_99_329 ();
 sg13g2_fill_2 FILLER_99_333 ();
 sg13g2_decap_8 FILLER_99_371 ();
 sg13g2_decap_8 FILLER_99_378 ();
 sg13g2_decap_8 FILLER_99_385 ();
 sg13g2_fill_1 FILLER_99_397 ();
 sg13g2_fill_2 FILLER_99_402 ();
 sg13g2_fill_2 FILLER_99_488 ();
 sg13g2_fill_2 FILLER_99_495 ();
 sg13g2_decap_4 FILLER_99_523 ();
 sg13g2_fill_1 FILLER_99_527 ();
 sg13g2_fill_1 FILLER_99_562 ();
 sg13g2_fill_2 FILLER_99_568 ();
 sg13g2_fill_2 FILLER_99_574 ();
 sg13g2_fill_2 FILLER_99_582 ();
 sg13g2_fill_1 FILLER_99_584 ();
 sg13g2_decap_4 FILLER_99_590 ();
 sg13g2_fill_1 FILLER_99_594 ();
 sg13g2_decap_8 FILLER_99_605 ();
 sg13g2_decap_8 FILLER_99_612 ();
 sg13g2_decap_8 FILLER_99_619 ();
 sg13g2_decap_4 FILLER_99_626 ();
 sg13g2_fill_2 FILLER_99_630 ();
 sg13g2_fill_2 FILLER_99_652 ();
 sg13g2_fill_1 FILLER_99_654 ();
 sg13g2_fill_2 FILLER_99_659 ();
 sg13g2_fill_2 FILLER_99_666 ();
 sg13g2_decap_4 FILLER_99_694 ();
 sg13g2_decap_4 FILLER_99_703 ();
 sg13g2_fill_2 FILLER_99_712 ();
 sg13g2_fill_1 FILLER_99_714 ();
 sg13g2_decap_4 FILLER_99_725 ();
 sg13g2_decap_8 FILLER_99_739 ();
 sg13g2_decap_8 FILLER_99_746 ();
 sg13g2_decap_8 FILLER_99_753 ();
 sg13g2_decap_8 FILLER_99_760 ();
 sg13g2_decap_8 FILLER_99_767 ();
 sg13g2_decap_4 FILLER_99_774 ();
 sg13g2_fill_1 FILLER_99_778 ();
 sg13g2_fill_2 FILLER_99_787 ();
 sg13g2_decap_4 FILLER_99_794 ();
 sg13g2_fill_1 FILLER_99_798 ();
 sg13g2_fill_1 FILLER_99_804 ();
 sg13g2_decap_4 FILLER_99_823 ();
 sg13g2_fill_2 FILLER_99_827 ();
 sg13g2_decap_8 FILLER_99_855 ();
 sg13g2_decap_8 FILLER_99_862 ();
 sg13g2_fill_2 FILLER_99_869 ();
 sg13g2_decap_8 FILLER_99_876 ();
 sg13g2_fill_1 FILLER_99_888 ();
 sg13g2_decap_4 FILLER_99_899 ();
 sg13g2_decap_8 FILLER_99_909 ();
 sg13g2_decap_8 FILLER_99_916 ();
 sg13g2_decap_8 FILLER_99_923 ();
 sg13g2_decap_8 FILLER_99_930 ();
 sg13g2_decap_8 FILLER_99_937 ();
 sg13g2_decap_8 FILLER_99_944 ();
 sg13g2_fill_2 FILLER_99_967 ();
 sg13g2_fill_1 FILLER_99_969 ();
 sg13g2_fill_2 FILLER_99_974 ();
 sg13g2_fill_1 FILLER_99_976 ();
 sg13g2_decap_8 FILLER_99_986 ();
 sg13g2_decap_4 FILLER_99_993 ();
 sg13g2_fill_2 FILLER_99_997 ();
 sg13g2_decap_8 FILLER_99_1017 ();
 sg13g2_fill_1 FILLER_99_1029 ();
 sg13g2_fill_1 FILLER_99_1038 ();
 sg13g2_decap_4 FILLER_99_1044 ();
 sg13g2_fill_2 FILLER_99_1052 ();
 sg13g2_fill_1 FILLER_99_1058 ();
 sg13g2_decap_8 FILLER_99_1064 ();
 sg13g2_fill_1 FILLER_99_1136 ();
 sg13g2_decap_4 FILLER_99_1161 ();
 sg13g2_fill_2 FILLER_99_1165 ();
 sg13g2_decap_4 FILLER_99_1185 ();
 sg13g2_fill_1 FILLER_99_1189 ();
 sg13g2_fill_1 FILLER_99_1195 ();
 sg13g2_fill_2 FILLER_99_1200 ();
 sg13g2_fill_1 FILLER_99_1202 ();
 sg13g2_fill_1 FILLER_99_1226 ();
 sg13g2_fill_1 FILLER_99_1231 ();
 sg13g2_fill_2 FILLER_99_1241 ();
 sg13g2_decap_4 FILLER_99_1263 ();
 sg13g2_fill_2 FILLER_99_1267 ();
 sg13g2_fill_1 FILLER_99_1277 ();
 sg13g2_fill_1 FILLER_99_1283 ();
 sg13g2_decap_8 FILLER_99_1367 ();
 sg13g2_decap_8 FILLER_99_1374 ();
 sg13g2_fill_1 FILLER_99_1381 ();
 sg13g2_decap_8 FILLER_99_1386 ();
 sg13g2_decap_8 FILLER_99_1393 ();
 sg13g2_decap_4 FILLER_99_1400 ();
 sg13g2_decap_4 FILLER_99_1430 ();
 sg13g2_fill_1 FILLER_99_1434 ();
 sg13g2_decap_8 FILLER_99_1465 ();
 sg13g2_decap_4 FILLER_99_1472 ();
 sg13g2_fill_1 FILLER_99_1476 ();
 sg13g2_decap_8 FILLER_99_1503 ();
 sg13g2_decap_8 FILLER_99_1510 ();
 sg13g2_decap_8 FILLER_99_1517 ();
 sg13g2_decap_8 FILLER_99_1524 ();
 sg13g2_decap_8 FILLER_99_1531 ();
 sg13g2_decap_8 FILLER_99_1538 ();
 sg13g2_decap_8 FILLER_99_1545 ();
 sg13g2_decap_8 FILLER_99_1552 ();
 sg13g2_decap_8 FILLER_99_1559 ();
 sg13g2_decap_8 FILLER_99_1566 ();
 sg13g2_decap_8 FILLER_99_1573 ();
 sg13g2_decap_8 FILLER_99_1580 ();
 sg13g2_decap_8 FILLER_99_1587 ();
 sg13g2_decap_8 FILLER_99_1594 ();
 sg13g2_decap_8 FILLER_99_1601 ();
 sg13g2_decap_8 FILLER_99_1608 ();
 sg13g2_decap_8 FILLER_99_1615 ();
 sg13g2_fill_2 FILLER_99_1622 ();
 sg13g2_fill_1 FILLER_99_1624 ();
 sg13g2_decap_8 FILLER_100_0 ();
 sg13g2_decap_8 FILLER_100_7 ();
 sg13g2_decap_8 FILLER_100_14 ();
 sg13g2_decap_4 FILLER_100_21 ();
 sg13g2_fill_2 FILLER_100_25 ();
 sg13g2_fill_1 FILLER_100_98 ();
 sg13g2_decap_8 FILLER_100_104 ();
 sg13g2_fill_2 FILLER_100_111 ();
 sg13g2_decap_8 FILLER_100_121 ();
 sg13g2_decap_8 FILLER_100_128 ();
 sg13g2_decap_8 FILLER_100_135 ();
 sg13g2_decap_8 FILLER_100_142 ();
 sg13g2_fill_2 FILLER_100_149 ();
 sg13g2_fill_1 FILLER_100_151 ();
 sg13g2_decap_4 FILLER_100_181 ();
 sg13g2_fill_1 FILLER_100_185 ();
 sg13g2_fill_2 FILLER_100_220 ();
 sg13g2_decap_8 FILLER_100_255 ();
 sg13g2_decap_4 FILLER_100_262 ();
 sg13g2_fill_1 FILLER_100_266 ();
 sg13g2_fill_1 FILLER_100_275 ();
 sg13g2_decap_8 FILLER_100_286 ();
 sg13g2_fill_2 FILLER_100_293 ();
 sg13g2_fill_1 FILLER_100_295 ();
 sg13g2_decap_4 FILLER_100_300 ();
 sg13g2_decap_4 FILLER_100_344 ();
 sg13g2_fill_2 FILLER_100_348 ();
 sg13g2_fill_2 FILLER_100_385 ();
 sg13g2_fill_2 FILLER_100_413 ();
 sg13g2_fill_1 FILLER_100_415 ();
 sg13g2_fill_1 FILLER_100_442 ();
 sg13g2_fill_2 FILLER_100_476 ();
 sg13g2_fill_1 FILLER_100_478 ();
 sg13g2_decap_8 FILLER_100_513 ();
 sg13g2_decap_8 FILLER_100_520 ();
 sg13g2_decap_4 FILLER_100_527 ();
 sg13g2_fill_1 FILLER_100_531 ();
 sg13g2_decap_8 FILLER_100_545 ();
 sg13g2_decap_4 FILLER_100_552 ();
 sg13g2_fill_1 FILLER_100_556 ();
 sg13g2_fill_1 FILLER_100_562 ();
 sg13g2_decap_4 FILLER_100_570 ();
 sg13g2_fill_1 FILLER_100_574 ();
 sg13g2_decap_8 FILLER_100_587 ();
 sg13g2_fill_1 FILLER_100_594 ();
 sg13g2_decap_8 FILLER_100_602 ();
 sg13g2_decap_8 FILLER_100_609 ();
 sg13g2_fill_2 FILLER_100_616 ();
 sg13g2_fill_1 FILLER_100_618 ();
 sg13g2_decap_8 FILLER_100_623 ();
 sg13g2_decap_8 FILLER_100_630 ();
 sg13g2_decap_8 FILLER_100_637 ();
 sg13g2_decap_4 FILLER_100_644 ();
 sg13g2_fill_1 FILLER_100_648 ();
 sg13g2_decap_8 FILLER_100_675 ();
 sg13g2_fill_2 FILLER_100_682 ();
 sg13g2_fill_1 FILLER_100_684 ();
 sg13g2_decap_8 FILLER_100_689 ();
 sg13g2_decap_8 FILLER_100_696 ();
 sg13g2_fill_1 FILLER_100_703 ();
 sg13g2_fill_2 FILLER_100_728 ();
 sg13g2_fill_1 FILLER_100_730 ();
 sg13g2_decap_4 FILLER_100_735 ();
 sg13g2_fill_1 FILLER_100_739 ();
 sg13g2_fill_2 FILLER_100_744 ();
 sg13g2_decap_4 FILLER_100_750 ();
 sg13g2_fill_1 FILLER_100_754 ();
 sg13g2_decap_8 FILLER_100_759 ();
 sg13g2_decap_8 FILLER_100_766 ();
 sg13g2_decap_8 FILLER_100_773 ();
 sg13g2_fill_2 FILLER_100_780 ();
 sg13g2_decap_8 FILLER_100_786 ();
 sg13g2_decap_8 FILLER_100_793 ();
 sg13g2_decap_8 FILLER_100_800 ();
 sg13g2_decap_8 FILLER_100_807 ();
 sg13g2_fill_1 FILLER_100_814 ();
 sg13g2_decap_8 FILLER_100_820 ();
 sg13g2_decap_8 FILLER_100_827 ();
 sg13g2_decap_8 FILLER_100_834 ();
 sg13g2_decap_8 FILLER_100_841 ();
 sg13g2_decap_8 FILLER_100_848 ();
 sg13g2_fill_2 FILLER_100_855 ();
 sg13g2_fill_2 FILLER_100_883 ();
 sg13g2_fill_1 FILLER_100_885 ();
 sg13g2_decap_4 FILLER_100_912 ();
 sg13g2_fill_1 FILLER_100_916 ();
 sg13g2_decap_4 FILLER_100_945 ();
 sg13g2_fill_1 FILLER_100_949 ();
 sg13g2_fill_1 FILLER_100_963 ();
 sg13g2_fill_2 FILLER_100_970 ();
 sg13g2_decap_8 FILLER_100_980 ();
 sg13g2_fill_1 FILLER_100_987 ();
 sg13g2_decap_4 FILLER_100_996 ();
 sg13g2_fill_2 FILLER_100_1000 ();
 sg13g2_decap_8 FILLER_100_1007 ();
 sg13g2_decap_4 FILLER_100_1014 ();
 sg13g2_fill_1 FILLER_100_1018 ();
 sg13g2_decap_4 FILLER_100_1040 ();
 sg13g2_fill_1 FILLER_100_1044 ();
 sg13g2_decap_8 FILLER_100_1049 ();
 sg13g2_decap_8 FILLER_100_1056 ();
 sg13g2_decap_8 FILLER_100_1063 ();
 sg13g2_fill_2 FILLER_100_1070 ();
 sg13g2_fill_2 FILLER_100_1103 ();
 sg13g2_decap_8 FILLER_100_1136 ();
 sg13g2_decap_4 FILLER_100_1162 ();
 sg13g2_fill_1 FILLER_100_1179 ();
 sg13g2_fill_1 FILLER_100_1185 ();
 sg13g2_fill_2 FILLER_100_1203 ();
 sg13g2_fill_1 FILLER_100_1205 ();
 sg13g2_fill_2 FILLER_100_1214 ();
 sg13g2_decap_8 FILLER_100_1221 ();
 sg13g2_decap_4 FILLER_100_1228 ();
 sg13g2_fill_2 FILLER_100_1232 ();
 sg13g2_fill_2 FILLER_100_1238 ();
 sg13g2_fill_2 FILLER_100_1304 ();
 sg13g2_fill_2 FILLER_100_1310 ();
 sg13g2_decap_8 FILLER_100_1380 ();
 sg13g2_decap_4 FILLER_100_1387 ();
 sg13g2_fill_2 FILLER_100_1391 ();
 sg13g2_decap_4 FILLER_100_1414 ();
 sg13g2_fill_2 FILLER_100_1418 ();
 sg13g2_fill_2 FILLER_100_1425 ();
 sg13g2_fill_1 FILLER_100_1453 ();
 sg13g2_decap_8 FILLER_100_1480 ();
 sg13g2_decap_8 FILLER_100_1487 ();
 sg13g2_decap_8 FILLER_100_1494 ();
 sg13g2_decap_8 FILLER_100_1501 ();
 sg13g2_decap_8 FILLER_100_1508 ();
 sg13g2_decap_8 FILLER_100_1515 ();
 sg13g2_decap_8 FILLER_100_1522 ();
 sg13g2_decap_8 FILLER_100_1529 ();
 sg13g2_decap_8 FILLER_100_1536 ();
 sg13g2_decap_8 FILLER_100_1543 ();
 sg13g2_decap_8 FILLER_100_1550 ();
 sg13g2_decap_8 FILLER_100_1557 ();
 sg13g2_decap_8 FILLER_100_1564 ();
 sg13g2_decap_8 FILLER_100_1571 ();
 sg13g2_decap_8 FILLER_100_1578 ();
 sg13g2_decap_8 FILLER_100_1585 ();
 sg13g2_decap_8 FILLER_100_1592 ();
 sg13g2_decap_8 FILLER_100_1599 ();
 sg13g2_decap_8 FILLER_100_1606 ();
 sg13g2_decap_8 FILLER_100_1613 ();
 sg13g2_decap_4 FILLER_100_1620 ();
 sg13g2_fill_1 FILLER_100_1624 ();
 sg13g2_decap_8 FILLER_101_0 ();
 sg13g2_decap_8 FILLER_101_7 ();
 sg13g2_decap_8 FILLER_101_14 ();
 sg13g2_decap_4 FILLER_101_21 ();
 sg13g2_fill_2 FILLER_101_25 ();
 sg13g2_decap_4 FILLER_101_53 ();
 sg13g2_fill_1 FILLER_101_57 ();
 sg13g2_decap_4 FILLER_101_96 ();
 sg13g2_decap_4 FILLER_101_108 ();
 sg13g2_fill_1 FILLER_101_112 ();
 sg13g2_decap_8 FILLER_101_128 ();
 sg13g2_fill_2 FILLER_101_135 ();
 sg13g2_fill_1 FILLER_101_137 ();
 sg13g2_decap_8 FILLER_101_142 ();
 sg13g2_fill_1 FILLER_101_149 ();
 sg13g2_decap_4 FILLER_101_160 ();
 sg13g2_fill_1 FILLER_101_164 ();
 sg13g2_decap_8 FILLER_101_191 ();
 sg13g2_decap_8 FILLER_101_198 ();
 sg13g2_decap_8 FILLER_101_205 ();
 sg13g2_fill_2 FILLER_101_212 ();
 sg13g2_fill_1 FILLER_101_214 ();
 sg13g2_decap_8 FILLER_101_230 ();
 sg13g2_fill_2 FILLER_101_237 ();
 sg13g2_decap_4 FILLER_101_270 ();
 sg13g2_fill_1 FILLER_101_274 ();
 sg13g2_decap_8 FILLER_101_285 ();
 sg13g2_decap_4 FILLER_101_292 ();
 sg13g2_decap_8 FILLER_101_300 ();
 sg13g2_fill_2 FILLER_101_307 ();
 sg13g2_fill_1 FILLER_101_309 ();
 sg13g2_decap_4 FILLER_101_335 ();
 sg13g2_decap_8 FILLER_101_377 ();
 sg13g2_decap_4 FILLER_101_384 ();
 sg13g2_fill_1 FILLER_101_388 ();
 sg13g2_decap_8 FILLER_101_393 ();
 sg13g2_decap_8 FILLER_101_400 ();
 sg13g2_decap_8 FILLER_101_407 ();
 sg13g2_decap_8 FILLER_101_414 ();
 sg13g2_decap_8 FILLER_101_421 ();
 sg13g2_decap_8 FILLER_101_467 ();
 sg13g2_decap_4 FILLER_101_474 ();
 sg13g2_fill_1 FILLER_101_478 ();
 sg13g2_decap_8 FILLER_101_509 ();
 sg13g2_fill_2 FILLER_101_516 ();
 sg13g2_fill_1 FILLER_101_518 ();
 sg13g2_decap_4 FILLER_101_523 ();
 sg13g2_fill_2 FILLER_101_527 ();
 sg13g2_decap_8 FILLER_101_566 ();
 sg13g2_decap_8 FILLER_101_573 ();
 sg13g2_decap_8 FILLER_101_580 ();
 sg13g2_decap_8 FILLER_101_587 ();
 sg13g2_fill_2 FILLER_101_594 ();
 sg13g2_fill_1 FILLER_101_596 ();
 sg13g2_decap_8 FILLER_101_601 ();
 sg13g2_decap_4 FILLER_101_608 ();
 sg13g2_decap_8 FILLER_101_638 ();
 sg13g2_fill_2 FILLER_101_645 ();
 sg13g2_decap_8 FILLER_101_703 ();
 sg13g2_decap_4 FILLER_101_718 ();
 sg13g2_fill_1 FILLER_101_722 ();
 sg13g2_decap_8 FILLER_101_805 ();
 sg13g2_fill_2 FILLER_101_812 ();
 sg13g2_fill_1 FILLER_101_814 ();
 sg13g2_decap_8 FILLER_101_819 ();
 sg13g2_decap_8 FILLER_101_826 ();
 sg13g2_decap_8 FILLER_101_833 ();
 sg13g2_fill_2 FILLER_101_846 ();
 sg13g2_decap_4 FILLER_101_877 ();
 sg13g2_fill_2 FILLER_101_881 ();
 sg13g2_decap_4 FILLER_101_921 ();
 sg13g2_fill_2 FILLER_101_925 ();
 sg13g2_decap_8 FILLER_101_970 ();
 sg13g2_decap_8 FILLER_101_977 ();
 sg13g2_decap_4 FILLER_101_984 ();
 sg13g2_decap_8 FILLER_101_993 ();
 sg13g2_decap_8 FILLER_101_1000 ();
 sg13g2_decap_8 FILLER_101_1007 ();
 sg13g2_decap_8 FILLER_101_1014 ();
 sg13g2_fill_1 FILLER_101_1027 ();
 sg13g2_fill_2 FILLER_101_1032 ();
 sg13g2_fill_1 FILLER_101_1034 ();
 sg13g2_fill_2 FILLER_101_1039 ();
 sg13g2_decap_4 FILLER_101_1051 ();
 sg13g2_fill_2 FILLER_101_1055 ();
 sg13g2_fill_2 FILLER_101_1066 ();
 sg13g2_fill_2 FILLER_101_1081 ();
 sg13g2_fill_1 FILLER_101_1083 ();
 sg13g2_fill_1 FILLER_101_1126 ();
 sg13g2_decap_8 FILLER_101_1137 ();
 sg13g2_fill_2 FILLER_101_1144 ();
 sg13g2_fill_1 FILLER_101_1146 ();
 sg13g2_fill_2 FILLER_101_1161 ();
 sg13g2_decap_8 FILLER_101_1168 ();
 sg13g2_decap_8 FILLER_101_1175 ();
 sg13g2_fill_1 FILLER_101_1182 ();
 sg13g2_decap_8 FILLER_101_1207 ();
 sg13g2_decap_8 FILLER_101_1214 ();
 sg13g2_decap_8 FILLER_101_1221 ();
 sg13g2_decap_8 FILLER_101_1228 ();
 sg13g2_decap_8 FILLER_101_1235 ();
 sg13g2_fill_1 FILLER_101_1242 ();
 sg13g2_decap_8 FILLER_101_1248 ();
 sg13g2_decap_4 FILLER_101_1255 ();
 sg13g2_fill_1 FILLER_101_1268 ();
 sg13g2_fill_2 FILLER_101_1327 ();
 sg13g2_decap_4 FILLER_101_1363 ();
 sg13g2_decap_8 FILLER_101_1393 ();
 sg13g2_decap_8 FILLER_101_1400 ();
 sg13g2_fill_2 FILLER_101_1407 ();
 sg13g2_decap_8 FILLER_101_1459 ();
 sg13g2_decap_4 FILLER_101_1466 ();
 sg13g2_decap_8 FILLER_101_1495 ();
 sg13g2_decap_8 FILLER_101_1502 ();
 sg13g2_decap_8 FILLER_101_1509 ();
 sg13g2_decap_8 FILLER_101_1516 ();
 sg13g2_decap_8 FILLER_101_1523 ();
 sg13g2_decap_8 FILLER_101_1530 ();
 sg13g2_decap_8 FILLER_101_1537 ();
 sg13g2_decap_8 FILLER_101_1544 ();
 sg13g2_decap_8 FILLER_101_1551 ();
 sg13g2_decap_8 FILLER_101_1558 ();
 sg13g2_decap_8 FILLER_101_1565 ();
 sg13g2_decap_8 FILLER_101_1572 ();
 sg13g2_decap_8 FILLER_101_1579 ();
 sg13g2_decap_8 FILLER_101_1586 ();
 sg13g2_decap_8 FILLER_101_1593 ();
 sg13g2_decap_8 FILLER_101_1600 ();
 sg13g2_decap_8 FILLER_101_1607 ();
 sg13g2_decap_8 FILLER_101_1614 ();
 sg13g2_decap_4 FILLER_101_1621 ();
 sg13g2_decap_8 FILLER_102_0 ();
 sg13g2_decap_8 FILLER_102_7 ();
 sg13g2_decap_8 FILLER_102_14 ();
 sg13g2_decap_8 FILLER_102_21 ();
 sg13g2_fill_2 FILLER_102_28 ();
 sg13g2_fill_1 FILLER_102_30 ();
 sg13g2_decap_8 FILLER_102_35 ();
 sg13g2_decap_8 FILLER_102_42 ();
 sg13g2_fill_2 FILLER_102_49 ();
 sg13g2_decap_8 FILLER_102_55 ();
 sg13g2_fill_1 FILLER_102_62 ();
 sg13g2_decap_8 FILLER_102_67 ();
 sg13g2_decap_8 FILLER_102_74 ();
 sg13g2_decap_8 FILLER_102_81 ();
 sg13g2_decap_8 FILLER_102_88 ();
 sg13g2_fill_2 FILLER_102_95 ();
 sg13g2_fill_1 FILLER_102_97 ();
 sg13g2_fill_2 FILLER_102_110 ();
 sg13g2_fill_2 FILLER_102_120 ();
 sg13g2_fill_1 FILLER_102_122 ();
 sg13g2_fill_1 FILLER_102_131 ();
 sg13g2_fill_2 FILLER_102_158 ();
 sg13g2_fill_1 FILLER_102_160 ();
 sg13g2_decap_8 FILLER_102_176 ();
 sg13g2_decap_8 FILLER_102_183 ();
 sg13g2_decap_8 FILLER_102_190 ();
 sg13g2_decap_8 FILLER_102_197 ();
 sg13g2_decap_8 FILLER_102_204 ();
 sg13g2_decap_4 FILLER_102_211 ();
 sg13g2_fill_1 FILLER_102_215 ();
 sg13g2_decap_4 FILLER_102_222 ();
 sg13g2_fill_2 FILLER_102_226 ();
 sg13g2_decap_8 FILLER_102_232 ();
 sg13g2_decap_8 FILLER_102_239 ();
 sg13g2_fill_2 FILLER_102_271 ();
 sg13g2_fill_1 FILLER_102_273 ();
 sg13g2_decap_4 FILLER_102_282 ();
 sg13g2_fill_2 FILLER_102_286 ();
 sg13g2_decap_4 FILLER_102_314 ();
 sg13g2_fill_1 FILLER_102_318 ();
 sg13g2_decap_4 FILLER_102_329 ();
 sg13g2_fill_1 FILLER_102_333 ();
 sg13g2_decap_8 FILLER_102_370 ();
 sg13g2_fill_2 FILLER_102_377 ();
 sg13g2_fill_1 FILLER_102_379 ();
 sg13g2_fill_2 FILLER_102_385 ();
 sg13g2_fill_1 FILLER_102_387 ();
 sg13g2_fill_1 FILLER_102_397 ();
 sg13g2_decap_8 FILLER_102_402 ();
 sg13g2_decap_4 FILLER_102_409 ();
 sg13g2_decap_8 FILLER_102_418 ();
 sg13g2_decap_8 FILLER_102_425 ();
 sg13g2_decap_4 FILLER_102_507 ();
 sg13g2_fill_2 FILLER_102_537 ();
 sg13g2_fill_1 FILLER_102_539 ();
 sg13g2_decap_8 FILLER_102_545 ();
 sg13g2_fill_2 FILLER_102_552 ();
 sg13g2_fill_1 FILLER_102_554 ();
 sg13g2_decap_4 FILLER_102_576 ();
 sg13g2_fill_2 FILLER_102_580 ();
 sg13g2_decap_4 FILLER_102_586 ();
 sg13g2_decap_8 FILLER_102_624 ();
 sg13g2_decap_4 FILLER_102_631 ();
 sg13g2_fill_2 FILLER_102_635 ();
 sg13g2_decap_8 FILLER_102_642 ();
 sg13g2_decap_8 FILLER_102_649 ();
 sg13g2_decap_4 FILLER_102_656 ();
 sg13g2_fill_2 FILLER_102_660 ();
 sg13g2_decap_8 FILLER_102_700 ();
 sg13g2_decap_8 FILLER_102_707 ();
 sg13g2_decap_8 FILLER_102_714 ();
 sg13g2_decap_8 FILLER_102_721 ();
 sg13g2_decap_4 FILLER_102_728 ();
 sg13g2_fill_1 FILLER_102_732 ();
 sg13g2_decap_8 FILLER_102_742 ();
 sg13g2_decap_8 FILLER_102_749 ();
 sg13g2_decap_4 FILLER_102_756 ();
 sg13g2_fill_2 FILLER_102_760 ();
 sg13g2_fill_2 FILLER_102_805 ();
 sg13g2_fill_1 FILLER_102_846 ();
 sg13g2_fill_1 FILLER_102_864 ();
 sg13g2_fill_2 FILLER_102_873 ();
 sg13g2_fill_1 FILLER_102_875 ();
 sg13g2_fill_1 FILLER_102_937 ();
 sg13g2_decap_4 FILLER_102_972 ();
 sg13g2_fill_2 FILLER_102_976 ();
 sg13g2_fill_2 FILLER_102_998 ();
 sg13g2_fill_2 FILLER_102_1005 ();
 sg13g2_fill_1 FILLER_102_1007 ();
 sg13g2_decap_8 FILLER_102_1013 ();
 sg13g2_decap_8 FILLER_102_1020 ();
 sg13g2_fill_2 FILLER_102_1027 ();
 sg13g2_decap_8 FILLER_102_1034 ();
 sg13g2_decap_4 FILLER_102_1053 ();
 sg13g2_decap_8 FILLER_102_1065 ();
 sg13g2_decap_8 FILLER_102_1077 ();
 sg13g2_fill_1 FILLER_102_1084 ();
 sg13g2_fill_2 FILLER_102_1090 ();
 sg13g2_fill_1 FILLER_102_1110 ();
 sg13g2_decap_4 FILLER_102_1123 ();
 sg13g2_fill_2 FILLER_102_1127 ();
 sg13g2_decap_8 FILLER_102_1142 ();
 sg13g2_decap_8 FILLER_102_1183 ();
 sg13g2_fill_2 FILLER_102_1190 ();
 sg13g2_fill_1 FILLER_102_1192 ();
 sg13g2_decap_8 FILLER_102_1201 ();
 sg13g2_decap_8 FILLER_102_1208 ();
 sg13g2_fill_1 FILLER_102_1215 ();
 sg13g2_decap_8 FILLER_102_1220 ();
 sg13g2_decap_8 FILLER_102_1227 ();
 sg13g2_decap_8 FILLER_102_1234 ();
 sg13g2_decap_8 FILLER_102_1241 ();
 sg13g2_decap_8 FILLER_102_1248 ();
 sg13g2_fill_2 FILLER_102_1255 ();
 sg13g2_fill_1 FILLER_102_1257 ();
 sg13g2_fill_1 FILLER_102_1263 ();
 sg13g2_decap_4 FILLER_102_1270 ();
 sg13g2_decap_4 FILLER_102_1282 ();
 sg13g2_fill_2 FILLER_102_1286 ();
 sg13g2_fill_2 FILLER_102_1318 ();
 sg13g2_fill_1 FILLER_102_1320 ();
 sg13g2_decap_4 FILLER_102_1368 ();
 sg13g2_fill_2 FILLER_102_1372 ();
 sg13g2_decap_8 FILLER_102_1378 ();
 sg13g2_decap_8 FILLER_102_1385 ();
 sg13g2_decap_8 FILLER_102_1444 ();
 sg13g2_decap_4 FILLER_102_1451 ();
 sg13g2_fill_1 FILLER_102_1455 ();
 sg13g2_decap_8 FILLER_102_1460 ();
 sg13g2_decap_8 FILLER_102_1467 ();
 sg13g2_decap_8 FILLER_102_1474 ();
 sg13g2_decap_8 FILLER_102_1481 ();
 sg13g2_decap_8 FILLER_102_1488 ();
 sg13g2_decap_8 FILLER_102_1495 ();
 sg13g2_decap_8 FILLER_102_1502 ();
 sg13g2_decap_8 FILLER_102_1509 ();
 sg13g2_decap_8 FILLER_102_1516 ();
 sg13g2_decap_8 FILLER_102_1523 ();
 sg13g2_decap_8 FILLER_102_1530 ();
 sg13g2_decap_8 FILLER_102_1537 ();
 sg13g2_decap_8 FILLER_102_1544 ();
 sg13g2_decap_8 FILLER_102_1551 ();
 sg13g2_decap_8 FILLER_102_1558 ();
 sg13g2_decap_8 FILLER_102_1565 ();
 sg13g2_decap_8 FILLER_102_1572 ();
 sg13g2_decap_8 FILLER_102_1579 ();
 sg13g2_decap_8 FILLER_102_1586 ();
 sg13g2_decap_8 FILLER_102_1593 ();
 sg13g2_decap_8 FILLER_102_1600 ();
 sg13g2_decap_8 FILLER_102_1607 ();
 sg13g2_decap_8 FILLER_102_1614 ();
 sg13g2_decap_4 FILLER_102_1621 ();
 sg13g2_decap_8 FILLER_103_0 ();
 sg13g2_decap_8 FILLER_103_7 ();
 sg13g2_decap_8 FILLER_103_14 ();
 sg13g2_decap_4 FILLER_103_21 ();
 sg13g2_fill_1 FILLER_103_51 ();
 sg13g2_decap_8 FILLER_103_82 ();
 sg13g2_decap_4 FILLER_103_89 ();
 sg13g2_decap_8 FILLER_103_101 ();
 sg13g2_decap_8 FILLER_103_108 ();
 sg13g2_decap_4 FILLER_103_115 ();
 sg13g2_fill_1 FILLER_103_119 ();
 sg13g2_decap_8 FILLER_103_130 ();
 sg13g2_decap_8 FILLER_103_137 ();
 sg13g2_decap_8 FILLER_103_144 ();
 sg13g2_decap_4 FILLER_103_151 ();
 sg13g2_fill_1 FILLER_103_155 ();
 sg13g2_decap_8 FILLER_103_161 ();
 sg13g2_decap_8 FILLER_103_168 ();
 sg13g2_decap_8 FILLER_103_175 ();
 sg13g2_fill_2 FILLER_103_182 ();
 sg13g2_fill_1 FILLER_103_184 ();
 sg13g2_fill_1 FILLER_103_211 ();
 sg13g2_decap_4 FILLER_103_246 ();
 sg13g2_fill_2 FILLER_103_250 ();
 sg13g2_decap_8 FILLER_103_274 ();
 sg13g2_decap_8 FILLER_103_281 ();
 sg13g2_fill_2 FILLER_103_288 ();
 sg13g2_fill_1 FILLER_103_290 ();
 sg13g2_decap_4 FILLER_103_295 ();
 sg13g2_fill_2 FILLER_103_299 ();
 sg13g2_decap_4 FILLER_103_313 ();
 sg13g2_fill_2 FILLER_103_317 ();
 sg13g2_decap_8 FILLER_103_323 ();
 sg13g2_fill_2 FILLER_103_330 ();
 sg13g2_decap_4 FILLER_103_357 ();
 sg13g2_fill_2 FILLER_103_361 ();
 sg13g2_decap_8 FILLER_103_367 ();
 sg13g2_decap_8 FILLER_103_374 ();
 sg13g2_decap_8 FILLER_103_381 ();
 sg13g2_fill_2 FILLER_103_388 ();
 sg13g2_fill_1 FILLER_103_416 ();
 sg13g2_decap_8 FILLER_103_468 ();
 sg13g2_decap_4 FILLER_103_475 ();
 sg13g2_decap_8 FILLER_103_482 ();
 sg13g2_fill_2 FILLER_103_489 ();
 sg13g2_fill_2 FILLER_103_495 ();
 sg13g2_fill_1 FILLER_103_497 ();
 sg13g2_decap_4 FILLER_103_516 ();
 sg13g2_fill_2 FILLER_103_520 ();
 sg13g2_decap_4 FILLER_103_527 ();
 sg13g2_decap_8 FILLER_103_560 ();
 sg13g2_decap_8 FILLER_103_567 ();
 sg13g2_decap_4 FILLER_103_604 ();
 sg13g2_fill_2 FILLER_103_616 ();
 sg13g2_fill_1 FILLER_103_618 ();
 sg13g2_decap_8 FILLER_103_628 ();
 sg13g2_decap_4 FILLER_103_648 ();
 sg13g2_fill_1 FILLER_103_652 ();
 sg13g2_decap_4 FILLER_103_657 ();
 sg13g2_fill_2 FILLER_103_661 ();
 sg13g2_fill_2 FILLER_103_673 ();
 sg13g2_fill_1 FILLER_103_675 ();
 sg13g2_fill_2 FILLER_103_684 ();
 sg13g2_fill_1 FILLER_103_686 ();
 sg13g2_decap_4 FILLER_103_705 ();
 sg13g2_fill_2 FILLER_103_718 ();
 sg13g2_fill_2 FILLER_103_724 ();
 sg13g2_decap_8 FILLER_103_763 ();
 sg13g2_fill_1 FILLER_103_770 ();
 sg13g2_decap_4 FILLER_103_779 ();
 sg13g2_fill_1 FILLER_103_783 ();
 sg13g2_fill_2 FILLER_103_790 ();
 sg13g2_fill_2 FILLER_103_802 ();
 sg13g2_decap_4 FILLER_103_838 ();
 sg13g2_decap_8 FILLER_103_846 ();
 sg13g2_fill_2 FILLER_103_853 ();
 sg13g2_fill_1 FILLER_103_855 ();
 sg13g2_decap_8 FILLER_103_865 ();
 sg13g2_fill_1 FILLER_103_872 ();
 sg13g2_decap_8 FILLER_103_877 ();
 sg13g2_fill_1 FILLER_103_884 ();
 sg13g2_decap_8 FILLER_103_914 ();
 sg13g2_fill_1 FILLER_103_921 ();
 sg13g2_fill_2 FILLER_103_948 ();
 sg13g2_fill_1 FILLER_103_950 ();
 sg13g2_decap_4 FILLER_103_977 ();
 sg13g2_decap_4 FILLER_103_988 ();
 sg13g2_fill_2 FILLER_103_992 ();
 sg13g2_fill_2 FILLER_103_999 ();
 sg13g2_fill_1 FILLER_103_1001 ();
 sg13g2_fill_2 FILLER_103_1031 ();
 sg13g2_fill_2 FILLER_103_1041 ();
 sg13g2_fill_2 FILLER_103_1048 ();
 sg13g2_fill_1 FILLER_103_1050 ();
 sg13g2_decap_8 FILLER_103_1061 ();
 sg13g2_fill_2 FILLER_103_1068 ();
 sg13g2_fill_1 FILLER_103_1070 ();
 sg13g2_decap_8 FILLER_103_1081 ();
 sg13g2_decap_4 FILLER_103_1088 ();
 sg13g2_fill_1 FILLER_103_1092 ();
 sg13g2_fill_1 FILLER_103_1111 ();
 sg13g2_decap_4 FILLER_103_1120 ();
 sg13g2_decap_8 FILLER_103_1140 ();
 sg13g2_decap_4 FILLER_103_1147 ();
 sg13g2_fill_1 FILLER_103_1159 ();
 sg13g2_decap_8 FILLER_103_1170 ();
 sg13g2_decap_8 FILLER_103_1177 ();
 sg13g2_decap_8 FILLER_103_1184 ();
 sg13g2_decap_8 FILLER_103_1191 ();
 sg13g2_decap_8 FILLER_103_1198 ();
 sg13g2_decap_4 FILLER_103_1205 ();
 sg13g2_fill_1 FILLER_103_1209 ();
 sg13g2_fill_1 FILLER_103_1236 ();
 sg13g2_decap_8 FILLER_103_1241 ();
 sg13g2_decap_8 FILLER_103_1248 ();
 sg13g2_decap_4 FILLER_103_1255 ();
 sg13g2_fill_2 FILLER_103_1259 ();
 sg13g2_fill_1 FILLER_103_1273 ();
 sg13g2_fill_2 FILLER_103_1279 ();
 sg13g2_fill_1 FILLER_103_1281 ();
 sg13g2_decap_4 FILLER_103_1290 ();
 sg13g2_fill_2 FILLER_103_1294 ();
 sg13g2_fill_1 FILLER_103_1310 ();
 sg13g2_decap_8 FILLER_103_1316 ();
 sg13g2_decap_4 FILLER_103_1323 ();
 sg13g2_decap_4 FILLER_103_1331 ();
 sg13g2_fill_1 FILLER_103_1335 ();
 sg13g2_decap_4 FILLER_103_1348 ();
 sg13g2_fill_2 FILLER_103_1352 ();
 sg13g2_decap_8 FILLER_103_1358 ();
 sg13g2_decap_8 FILLER_103_1365 ();
 sg13g2_decap_8 FILLER_103_1372 ();
 sg13g2_decap_8 FILLER_103_1379 ();
 sg13g2_decap_8 FILLER_103_1386 ();
 sg13g2_decap_8 FILLER_103_1393 ();
 sg13g2_decap_8 FILLER_103_1400 ();
 sg13g2_decap_4 FILLER_103_1407 ();
 sg13g2_fill_2 FILLER_103_1411 ();
 sg13g2_decap_8 FILLER_103_1471 ();
 sg13g2_decap_8 FILLER_103_1478 ();
 sg13g2_decap_8 FILLER_103_1485 ();
 sg13g2_decap_8 FILLER_103_1492 ();
 sg13g2_decap_8 FILLER_103_1499 ();
 sg13g2_decap_8 FILLER_103_1506 ();
 sg13g2_decap_8 FILLER_103_1513 ();
 sg13g2_decap_8 FILLER_103_1520 ();
 sg13g2_decap_8 FILLER_103_1527 ();
 sg13g2_decap_8 FILLER_103_1534 ();
 sg13g2_decap_8 FILLER_103_1541 ();
 sg13g2_decap_8 FILLER_103_1548 ();
 sg13g2_decap_8 FILLER_103_1555 ();
 sg13g2_decap_8 FILLER_103_1562 ();
 sg13g2_decap_8 FILLER_103_1569 ();
 sg13g2_decap_8 FILLER_103_1576 ();
 sg13g2_decap_8 FILLER_103_1583 ();
 sg13g2_decap_8 FILLER_103_1590 ();
 sg13g2_decap_8 FILLER_103_1597 ();
 sg13g2_decap_8 FILLER_103_1604 ();
 sg13g2_decap_8 FILLER_103_1611 ();
 sg13g2_decap_8 FILLER_103_1618 ();
 sg13g2_decap_8 FILLER_104_0 ();
 sg13g2_decap_8 FILLER_104_7 ();
 sg13g2_decap_8 FILLER_104_14 ();
 sg13g2_decap_8 FILLER_104_21 ();
 sg13g2_decap_8 FILLER_104_28 ();
 sg13g2_decap_8 FILLER_104_35 ();
 sg13g2_fill_2 FILLER_104_42 ();
 sg13g2_fill_1 FILLER_104_44 ();
 sg13g2_decap_4 FILLER_104_70 ();
 sg13g2_decap_8 FILLER_104_77 ();
 sg13g2_decap_8 FILLER_104_84 ();
 sg13g2_decap_4 FILLER_104_91 ();
 sg13g2_fill_2 FILLER_104_95 ();
 sg13g2_decap_8 FILLER_104_105 ();
 sg13g2_decap_4 FILLER_104_112 ();
 sg13g2_decap_8 FILLER_104_121 ();
 sg13g2_decap_8 FILLER_104_128 ();
 sg13g2_decap_8 FILLER_104_135 ();
 sg13g2_decap_8 FILLER_104_142 ();
 sg13g2_decap_8 FILLER_104_149 ();
 sg13g2_fill_2 FILLER_104_169 ();
 sg13g2_fill_1 FILLER_104_171 ();
 sg13g2_decap_8 FILLER_104_176 ();
 sg13g2_decap_8 FILLER_104_183 ();
 sg13g2_decap_4 FILLER_104_190 ();
 sg13g2_decap_8 FILLER_104_199 ();
 sg13g2_fill_2 FILLER_104_206 ();
 sg13g2_fill_1 FILLER_104_208 ();
 sg13g2_decap_8 FILLER_104_224 ();
 sg13g2_decap_8 FILLER_104_231 ();
 sg13g2_decap_8 FILLER_104_238 ();
 sg13g2_fill_1 FILLER_104_245 ();
 sg13g2_fill_1 FILLER_104_251 ();
 sg13g2_fill_2 FILLER_104_256 ();
 sg13g2_fill_1 FILLER_104_258 ();
 sg13g2_decap_4 FILLER_104_267 ();
 sg13g2_fill_1 FILLER_104_271 ();
 sg13g2_decap_8 FILLER_104_280 ();
 sg13g2_fill_2 FILLER_104_299 ();
 sg13g2_fill_1 FILLER_104_305 ();
 sg13g2_fill_2 FILLER_104_337 ();
 sg13g2_fill_1 FILLER_104_339 ();
 sg13g2_decap_8 FILLER_104_344 ();
 sg13g2_decap_4 FILLER_104_351 ();
 sg13g2_fill_1 FILLER_104_355 ();
 sg13g2_fill_1 FILLER_104_382 ();
 sg13g2_decap_4 FILLER_104_387 ();
 sg13g2_decap_4 FILLER_104_396 ();
 sg13g2_fill_1 FILLER_104_400 ();
 sg13g2_decap_8 FILLER_104_411 ();
 sg13g2_decap_4 FILLER_104_418 ();
 sg13g2_fill_2 FILLER_104_422 ();
 sg13g2_fill_2 FILLER_104_428 ();
 sg13g2_decap_4 FILLER_104_477 ();
 sg13g2_fill_2 FILLER_104_486 ();
 sg13g2_fill_1 FILLER_104_488 ();
 sg13g2_decap_8 FILLER_104_494 ();
 sg13g2_decap_4 FILLER_104_501 ();
 sg13g2_fill_2 FILLER_104_505 ();
 sg13g2_decap_8 FILLER_104_511 ();
 sg13g2_decap_8 FILLER_104_568 ();
 sg13g2_decap_8 FILLER_104_575 ();
 sg13g2_decap_4 FILLER_104_582 ();
 sg13g2_fill_2 FILLER_104_586 ();
 sg13g2_decap_8 FILLER_104_613 ();
 sg13g2_fill_1 FILLER_104_620 ();
 sg13g2_fill_1 FILLER_104_629 ();
 sg13g2_decap_8 FILLER_104_635 ();
 sg13g2_fill_2 FILLER_104_642 ();
 sg13g2_fill_2 FILLER_104_670 ();
 sg13g2_fill_1 FILLER_104_672 ();
 sg13g2_fill_1 FILLER_104_678 ();
 sg13g2_fill_2 FILLER_104_685 ();
 sg13g2_decap_8 FILLER_104_697 ();
 sg13g2_decap_8 FILLER_104_704 ();
 sg13g2_decap_8 FILLER_104_711 ();
 sg13g2_fill_2 FILLER_104_718 ();
 sg13g2_fill_1 FILLER_104_720 ();
 sg13g2_decap_4 FILLER_104_745 ();
 sg13g2_decap_8 FILLER_104_753 ();
 sg13g2_decap_4 FILLER_104_760 ();
 sg13g2_fill_2 FILLER_104_764 ();
 sg13g2_fill_1 FILLER_104_780 ();
 sg13g2_decap_8 FILLER_104_797 ();
 sg13g2_decap_8 FILLER_104_804 ();
 sg13g2_decap_8 FILLER_104_811 ();
 sg13g2_fill_2 FILLER_104_818 ();
 sg13g2_fill_2 FILLER_104_828 ();
 sg13g2_fill_1 FILLER_104_838 ();
 sg13g2_fill_2 FILLER_104_848 ();
 sg13g2_decap_8 FILLER_104_858 ();
 sg13g2_fill_1 FILLER_104_865 ();
 sg13g2_fill_2 FILLER_104_918 ();
 sg13g2_decap_8 FILLER_104_924 ();
 sg13g2_fill_2 FILLER_104_931 ();
 sg13g2_fill_2 FILLER_104_966 ();
 sg13g2_fill_1 FILLER_104_968 ();
 sg13g2_decap_8 FILLER_104_980 ();
 sg13g2_decap_8 FILLER_104_987 ();
 sg13g2_fill_1 FILLER_104_994 ();
 sg13g2_decap_8 FILLER_104_999 ();
 sg13g2_decap_8 FILLER_104_1006 ();
 sg13g2_decap_8 FILLER_104_1013 ();
 sg13g2_decap_8 FILLER_104_1020 ();
 sg13g2_fill_1 FILLER_104_1031 ();
 sg13g2_decap_4 FILLER_104_1037 ();
 sg13g2_fill_2 FILLER_104_1041 ();
 sg13g2_decap_8 FILLER_104_1053 ();
 sg13g2_decap_4 FILLER_104_1060 ();
 sg13g2_fill_1 FILLER_104_1064 ();
 sg13g2_fill_1 FILLER_104_1082 ();
 sg13g2_decap_8 FILLER_104_1098 ();
 sg13g2_fill_1 FILLER_104_1105 ();
 sg13g2_decap_8 FILLER_104_1124 ();
 sg13g2_decap_8 FILLER_104_1131 ();
 sg13g2_decap_8 FILLER_104_1138 ();
 sg13g2_decap_8 FILLER_104_1145 ();
 sg13g2_decap_8 FILLER_104_1152 ();
 sg13g2_fill_2 FILLER_104_1159 ();
 sg13g2_fill_1 FILLER_104_1161 ();
 sg13g2_decap_4 FILLER_104_1172 ();
 sg13g2_fill_2 FILLER_104_1176 ();
 sg13g2_decap_4 FILLER_104_1188 ();
 sg13g2_decap_8 FILLER_104_1197 ();
 sg13g2_fill_1 FILLER_104_1204 ();
 sg13g2_fill_2 FILLER_104_1219 ();
 sg13g2_fill_2 FILLER_104_1225 ();
 sg13g2_fill_1 FILLER_104_1227 ();
 sg13g2_fill_2 FILLER_104_1254 ();
 sg13g2_fill_2 FILLER_104_1260 ();
 sg13g2_fill_1 FILLER_104_1262 ();
 sg13g2_fill_1 FILLER_104_1300 ();
 sg13g2_fill_1 FILLER_104_1309 ();
 sg13g2_fill_1 FILLER_104_1318 ();
 sg13g2_decap_4 FILLER_104_1331 ();
 sg13g2_fill_2 FILLER_104_1335 ();
 sg13g2_decap_8 FILLER_104_1363 ();
 sg13g2_fill_1 FILLER_104_1370 ();
 sg13g2_fill_1 FILLER_104_1380 ();
 sg13g2_fill_2 FILLER_104_1385 ();
 sg13g2_fill_1 FILLER_104_1387 ();
 sg13g2_fill_2 FILLER_104_1393 ();
 sg13g2_fill_1 FILLER_104_1395 ();
 sg13g2_decap_8 FILLER_104_1404 ();
 sg13g2_fill_2 FILLER_104_1420 ();
 sg13g2_decap_8 FILLER_104_1473 ();
 sg13g2_decap_8 FILLER_104_1480 ();
 sg13g2_decap_8 FILLER_104_1487 ();
 sg13g2_decap_8 FILLER_104_1494 ();
 sg13g2_decap_8 FILLER_104_1501 ();
 sg13g2_decap_8 FILLER_104_1508 ();
 sg13g2_decap_8 FILLER_104_1515 ();
 sg13g2_decap_8 FILLER_104_1522 ();
 sg13g2_decap_8 FILLER_104_1529 ();
 sg13g2_decap_8 FILLER_104_1536 ();
 sg13g2_decap_8 FILLER_104_1543 ();
 sg13g2_decap_8 FILLER_104_1550 ();
 sg13g2_decap_8 FILLER_104_1557 ();
 sg13g2_decap_8 FILLER_104_1564 ();
 sg13g2_decap_8 FILLER_104_1571 ();
 sg13g2_decap_8 FILLER_104_1578 ();
 sg13g2_decap_8 FILLER_104_1585 ();
 sg13g2_decap_8 FILLER_104_1592 ();
 sg13g2_decap_8 FILLER_104_1599 ();
 sg13g2_decap_8 FILLER_104_1606 ();
 sg13g2_decap_8 FILLER_104_1613 ();
 sg13g2_decap_4 FILLER_104_1620 ();
 sg13g2_fill_1 FILLER_104_1624 ();
 sg13g2_decap_8 FILLER_105_0 ();
 sg13g2_decap_8 FILLER_105_7 ();
 sg13g2_decap_8 FILLER_105_14 ();
 sg13g2_decap_8 FILLER_105_21 ();
 sg13g2_decap_8 FILLER_105_28 ();
 sg13g2_decap_8 FILLER_105_35 ();
 sg13g2_decap_4 FILLER_105_42 ();
 sg13g2_fill_1 FILLER_105_46 ();
 sg13g2_decap_4 FILLER_105_67 ();
 sg13g2_decap_4 FILLER_105_81 ();
 sg13g2_decap_4 FILLER_105_93 ();
 sg13g2_decap_4 FILLER_105_134 ();
 sg13g2_fill_2 FILLER_105_138 ();
 sg13g2_decap_4 FILLER_105_191 ();
 sg13g2_fill_2 FILLER_105_195 ();
 sg13g2_fill_2 FILLER_105_212 ();
 sg13g2_fill_1 FILLER_105_214 ();
 sg13g2_decap_4 FILLER_105_220 ();
 sg13g2_fill_2 FILLER_105_224 ();
 sg13g2_decap_8 FILLER_105_231 ();
 sg13g2_decap_8 FILLER_105_238 ();
 sg13g2_fill_1 FILLER_105_251 ();
 sg13g2_decap_4 FILLER_105_272 ();
 sg13g2_decap_8 FILLER_105_280 ();
 sg13g2_decap_8 FILLER_105_287 ();
 sg13g2_decap_8 FILLER_105_294 ();
 sg13g2_decap_8 FILLER_105_301 ();
 sg13g2_fill_1 FILLER_105_308 ();
 sg13g2_decap_8 FILLER_105_364 ();
 sg13g2_decap_8 FILLER_105_371 ();
 sg13g2_fill_2 FILLER_105_378 ();
 sg13g2_fill_1 FILLER_105_380 ();
 sg13g2_decap_8 FILLER_105_411 ();
 sg13g2_fill_2 FILLER_105_418 ();
 sg13g2_fill_1 FILLER_105_420 ();
 sg13g2_decap_8 FILLER_105_425 ();
 sg13g2_decap_4 FILLER_105_432 ();
 sg13g2_fill_1 FILLER_105_436 ();
 sg13g2_fill_2 FILLER_105_499 ();
 sg13g2_fill_2 FILLER_105_527 ();
 sg13g2_decap_4 FILLER_105_538 ();
 sg13g2_fill_2 FILLER_105_551 ();
 sg13g2_fill_2 FILLER_105_578 ();
 sg13g2_fill_1 FILLER_105_580 ();
 sg13g2_fill_2 FILLER_105_585 ();
 sg13g2_fill_1 FILLER_105_587 ();
 sg13g2_fill_1 FILLER_105_592 ();
 sg13g2_decap_8 FILLER_105_629 ();
 sg13g2_decap_8 FILLER_105_636 ();
 sg13g2_decap_8 FILLER_105_643 ();
 sg13g2_fill_2 FILLER_105_650 ();
 sg13g2_fill_1 FILLER_105_652 ();
 sg13g2_decap_8 FILLER_105_658 ();
 sg13g2_fill_2 FILLER_105_665 ();
 sg13g2_decap_4 FILLER_105_672 ();
 sg13g2_fill_1 FILLER_105_676 ();
 sg13g2_decap_8 FILLER_105_681 ();
 sg13g2_fill_2 FILLER_105_688 ();
 sg13g2_decap_8 FILLER_105_694 ();
 sg13g2_fill_2 FILLER_105_701 ();
 sg13g2_fill_1 FILLER_105_703 ();
 sg13g2_fill_2 FILLER_105_712 ();
 sg13g2_fill_1 FILLER_105_714 ();
 sg13g2_decap_8 FILLER_105_723 ();
 sg13g2_fill_2 FILLER_105_730 ();
 sg13g2_fill_1 FILLER_105_732 ();
 sg13g2_decap_8 FILLER_105_767 ();
 sg13g2_decap_4 FILLER_105_774 ();
 sg13g2_decap_8 FILLER_105_791 ();
 sg13g2_fill_1 FILLER_105_798 ();
 sg13g2_decap_8 FILLER_105_821 ();
 sg13g2_decap_8 FILLER_105_828 ();
 sg13g2_decap_4 FILLER_105_835 ();
 sg13g2_fill_2 FILLER_105_839 ();
 sg13g2_decap_8 FILLER_105_851 ();
 sg13g2_fill_2 FILLER_105_877 ();
 sg13g2_fill_1 FILLER_105_879 ();
 sg13g2_decap_4 FILLER_105_1014 ();
 sg13g2_decap_8 FILLER_105_1027 ();
 sg13g2_fill_2 FILLER_105_1034 ();
 sg13g2_fill_1 FILLER_105_1036 ();
 sg13g2_decap_8 FILLER_105_1055 ();
 sg13g2_decap_8 FILLER_105_1062 ();
 sg13g2_decap_8 FILLER_105_1069 ();
 sg13g2_decap_8 FILLER_105_1076 ();
 sg13g2_fill_1 FILLER_105_1083 ();
 sg13g2_fill_1 FILLER_105_1099 ();
 sg13g2_decap_4 FILLER_105_1105 ();
 sg13g2_decap_8 FILLER_105_1114 ();
 sg13g2_decap_8 FILLER_105_1121 ();
 sg13g2_decap_4 FILLER_105_1128 ();
 sg13g2_fill_2 FILLER_105_1132 ();
 sg13g2_decap_8 FILLER_105_1142 ();
 sg13g2_decap_4 FILLER_105_1154 ();
 sg13g2_decap_4 FILLER_105_1163 ();
 sg13g2_fill_2 FILLER_105_1189 ();
 sg13g2_decap_8 FILLER_105_1201 ();
 sg13g2_decap_4 FILLER_105_1208 ();
 sg13g2_decap_8 FILLER_105_1238 ();
 sg13g2_fill_2 FILLER_105_1245 ();
 sg13g2_fill_1 FILLER_105_1247 ();
 sg13g2_fill_2 FILLER_105_1284 ();
 sg13g2_decap_8 FILLER_105_1311 ();
 sg13g2_decap_4 FILLER_105_1326 ();
 sg13g2_fill_2 FILLER_105_1330 ();
 sg13g2_fill_2 FILLER_105_1414 ();
 sg13g2_fill_1 FILLER_105_1416 ();
 sg13g2_decap_8 FILLER_105_1468 ();
 sg13g2_decap_8 FILLER_105_1475 ();
 sg13g2_decap_8 FILLER_105_1482 ();
 sg13g2_decap_8 FILLER_105_1489 ();
 sg13g2_decap_8 FILLER_105_1496 ();
 sg13g2_decap_8 FILLER_105_1503 ();
 sg13g2_decap_8 FILLER_105_1510 ();
 sg13g2_decap_8 FILLER_105_1517 ();
 sg13g2_decap_8 FILLER_105_1524 ();
 sg13g2_decap_8 FILLER_105_1531 ();
 sg13g2_decap_8 FILLER_105_1538 ();
 sg13g2_decap_8 FILLER_105_1545 ();
 sg13g2_decap_8 FILLER_105_1552 ();
 sg13g2_decap_8 FILLER_105_1559 ();
 sg13g2_decap_8 FILLER_105_1566 ();
 sg13g2_decap_8 FILLER_105_1573 ();
 sg13g2_decap_8 FILLER_105_1580 ();
 sg13g2_decap_8 FILLER_105_1587 ();
 sg13g2_decap_8 FILLER_105_1594 ();
 sg13g2_decap_8 FILLER_105_1601 ();
 sg13g2_decap_8 FILLER_105_1608 ();
 sg13g2_decap_8 FILLER_105_1615 ();
 sg13g2_fill_2 FILLER_105_1622 ();
 sg13g2_fill_1 FILLER_105_1624 ();
 sg13g2_decap_8 FILLER_106_0 ();
 sg13g2_decap_8 FILLER_106_7 ();
 sg13g2_decap_8 FILLER_106_14 ();
 sg13g2_decap_8 FILLER_106_21 ();
 sg13g2_decap_8 FILLER_106_28 ();
 sg13g2_fill_1 FILLER_106_35 ();
 sg13g2_fill_2 FILLER_106_44 ();
 sg13g2_fill_1 FILLER_106_46 ();
 sg13g2_fill_2 FILLER_106_55 ();
 sg13g2_fill_1 FILLER_106_57 ();
 sg13g2_fill_1 FILLER_106_82 ();
 sg13g2_fill_1 FILLER_106_93 ();
 sg13g2_fill_2 FILLER_106_105 ();
 sg13g2_fill_1 FILLER_106_107 ();
 sg13g2_decap_8 FILLER_106_127 ();
 sg13g2_decap_8 FILLER_106_160 ();
 sg13g2_decap_8 FILLER_106_167 ();
 sg13g2_decap_8 FILLER_106_174 ();
 sg13g2_decap_8 FILLER_106_181 ();
 sg13g2_decap_8 FILLER_106_188 ();
 sg13g2_decap_8 FILLER_106_195 ();
 sg13g2_decap_4 FILLER_106_202 ();
 sg13g2_fill_1 FILLER_106_206 ();
 sg13g2_fill_2 FILLER_106_217 ();
 sg13g2_fill_1 FILLER_106_219 ();
 sg13g2_fill_1 FILLER_106_227 ();
 sg13g2_fill_2 FILLER_106_242 ();
 sg13g2_fill_1 FILLER_106_244 ();
 sg13g2_decap_8 FILLER_106_278 ();
 sg13g2_decap_4 FILLER_106_304 ();
 sg13g2_fill_1 FILLER_106_308 ();
 sg13g2_decap_4 FILLER_106_322 ();
 sg13g2_fill_2 FILLER_106_326 ();
 sg13g2_decap_8 FILLER_106_363 ();
 sg13g2_fill_2 FILLER_106_370 ();
 sg13g2_decap_8 FILLER_106_397 ();
 sg13g2_decap_4 FILLER_106_404 ();
 sg13g2_fill_2 FILLER_106_408 ();
 sg13g2_decap_8 FILLER_106_435 ();
 sg13g2_decap_4 FILLER_106_442 ();
 sg13g2_fill_2 FILLER_106_446 ();
 sg13g2_fill_2 FILLER_106_452 ();
 sg13g2_decap_8 FILLER_106_459 ();
 sg13g2_fill_2 FILLER_106_466 ();
 sg13g2_fill_1 FILLER_106_468 ();
 sg13g2_decap_8 FILLER_106_473 ();
 sg13g2_fill_1 FILLER_106_480 ();
 sg13g2_fill_2 FILLER_106_494 ();
 sg13g2_fill_1 FILLER_106_501 ();
 sg13g2_decap_8 FILLER_106_506 ();
 sg13g2_decap_4 FILLER_106_513 ();
 sg13g2_fill_1 FILLER_106_517 ();
 sg13g2_decap_4 FILLER_106_556 ();
 sg13g2_fill_2 FILLER_106_560 ();
 sg13g2_fill_2 FILLER_106_567 ();
 sg13g2_fill_1 FILLER_106_569 ();
 sg13g2_decap_4 FILLER_106_600 ();
 sg13g2_decap_8 FILLER_106_614 ();
 sg13g2_fill_2 FILLER_106_621 ();
 sg13g2_decap_8 FILLER_106_633 ();
 sg13g2_fill_1 FILLER_106_648 ();
 sg13g2_fill_2 FILLER_106_679 ();
 sg13g2_decap_8 FILLER_106_707 ();
 sg13g2_decap_8 FILLER_106_714 ();
 sg13g2_decap_4 FILLER_106_721 ();
 sg13g2_fill_1 FILLER_106_725 ();
 sg13g2_decap_8 FILLER_106_759 ();
 sg13g2_fill_1 FILLER_106_766 ();
 sg13g2_decap_8 FILLER_106_771 ();
 sg13g2_decap_8 FILLER_106_778 ();
 sg13g2_decap_4 FILLER_106_785 ();
 sg13g2_decap_8 FILLER_106_797 ();
 sg13g2_fill_2 FILLER_106_804 ();
 sg13g2_fill_1 FILLER_106_806 ();
 sg13g2_decap_8 FILLER_106_821 ();
 sg13g2_decap_4 FILLER_106_833 ();
 sg13g2_decap_8 FILLER_106_844 ();
 sg13g2_decap_8 FILLER_106_851 ();
 sg13g2_fill_1 FILLER_106_858 ();
 sg13g2_fill_2 FILLER_106_866 ();
 sg13g2_fill_1 FILLER_106_868 ();
 sg13g2_decap_8 FILLER_106_880 ();
 sg13g2_decap_4 FILLER_106_887 ();
 sg13g2_fill_1 FILLER_106_891 ();
 sg13g2_decap_8 FILLER_106_930 ();
 sg13g2_decap_4 FILLER_106_942 ();
 sg13g2_fill_2 FILLER_106_959 ();
 sg13g2_decap_8 FILLER_106_996 ();
 sg13g2_decap_8 FILLER_106_1003 ();
 sg13g2_decap_8 FILLER_106_1036 ();
 sg13g2_decap_8 FILLER_106_1043 ();
 sg13g2_decap_8 FILLER_106_1050 ();
 sg13g2_fill_1 FILLER_106_1057 ();
 sg13g2_decap_8 FILLER_106_1062 ();
 sg13g2_decap_8 FILLER_106_1069 ();
 sg13g2_decap_8 FILLER_106_1076 ();
 sg13g2_decap_4 FILLER_106_1083 ();
 sg13g2_decap_4 FILLER_106_1102 ();
 sg13g2_fill_1 FILLER_106_1106 ();
 sg13g2_fill_1 FILLER_106_1125 ();
 sg13g2_decap_8 FILLER_106_1136 ();
 sg13g2_fill_2 FILLER_106_1143 ();
 sg13g2_fill_1 FILLER_106_1150 ();
 sg13g2_fill_2 FILLER_106_1161 ();
 sg13g2_fill_1 FILLER_106_1163 ();
 sg13g2_decap_8 FILLER_106_1177 ();
 sg13g2_decap_8 FILLER_106_1184 ();
 sg13g2_fill_1 FILLER_106_1201 ();
 sg13g2_decap_4 FILLER_106_1209 ();
 sg13g2_fill_2 FILLER_106_1242 ();
 sg13g2_decap_4 FILLER_106_1269 ();
 sg13g2_fill_2 FILLER_106_1313 ();
 sg13g2_fill_1 FILLER_106_1327 ();
 sg13g2_decap_4 FILLER_106_1333 ();
 sg13g2_fill_2 FILLER_106_1337 ();
 sg13g2_decap_8 FILLER_106_1365 ();
 sg13g2_fill_2 FILLER_106_1372 ();
 sg13g2_fill_1 FILLER_106_1379 ();
 sg13g2_fill_1 FILLER_106_1405 ();
 sg13g2_fill_1 FILLER_106_1441 ();
 sg13g2_decap_8 FILLER_106_1446 ();
 sg13g2_decap_8 FILLER_106_1453 ();
 sg13g2_decap_8 FILLER_106_1460 ();
 sg13g2_decap_8 FILLER_106_1467 ();
 sg13g2_decap_8 FILLER_106_1474 ();
 sg13g2_decap_8 FILLER_106_1481 ();
 sg13g2_decap_8 FILLER_106_1488 ();
 sg13g2_decap_8 FILLER_106_1495 ();
 sg13g2_decap_8 FILLER_106_1502 ();
 sg13g2_decap_8 FILLER_106_1509 ();
 sg13g2_decap_8 FILLER_106_1516 ();
 sg13g2_decap_8 FILLER_106_1523 ();
 sg13g2_decap_8 FILLER_106_1530 ();
 sg13g2_decap_8 FILLER_106_1537 ();
 sg13g2_decap_8 FILLER_106_1544 ();
 sg13g2_decap_8 FILLER_106_1551 ();
 sg13g2_decap_8 FILLER_106_1558 ();
 sg13g2_decap_8 FILLER_106_1565 ();
 sg13g2_decap_8 FILLER_106_1572 ();
 sg13g2_decap_8 FILLER_106_1579 ();
 sg13g2_decap_8 FILLER_106_1586 ();
 sg13g2_decap_8 FILLER_106_1593 ();
 sg13g2_decap_8 FILLER_106_1600 ();
 sg13g2_decap_8 FILLER_106_1607 ();
 sg13g2_decap_8 FILLER_106_1614 ();
 sg13g2_decap_4 FILLER_106_1621 ();
 sg13g2_decap_8 FILLER_107_0 ();
 sg13g2_decap_8 FILLER_107_7 ();
 sg13g2_decap_8 FILLER_107_14 ();
 sg13g2_decap_8 FILLER_107_21 ();
 sg13g2_fill_2 FILLER_107_28 ();
 sg13g2_fill_1 FILLER_107_30 ();
 sg13g2_decap_8 FILLER_107_57 ();
 sg13g2_decap_8 FILLER_107_64 ();
 sg13g2_decap_4 FILLER_107_71 ();
 sg13g2_decap_4 FILLER_107_83 ();
 sg13g2_decap_4 FILLER_107_92 ();
 sg13g2_fill_2 FILLER_107_96 ();
 sg13g2_fill_2 FILLER_107_109 ();
 sg13g2_fill_1 FILLER_107_116 ();
 sg13g2_decap_8 FILLER_107_124 ();
 sg13g2_decap_8 FILLER_107_131 ();
 sg13g2_fill_2 FILLER_107_138 ();
 sg13g2_fill_1 FILLER_107_140 ();
 sg13g2_decap_8 FILLER_107_145 ();
 sg13g2_decap_4 FILLER_107_152 ();
 sg13g2_decap_8 FILLER_107_160 ();
 sg13g2_decap_4 FILLER_107_167 ();
 sg13g2_fill_1 FILLER_107_171 ();
 sg13g2_fill_2 FILLER_107_180 ();
 sg13g2_decap_8 FILLER_107_211 ();
 sg13g2_decap_8 FILLER_107_218 ();
 sg13g2_fill_2 FILLER_107_225 ();
 sg13g2_fill_2 FILLER_107_316 ();
 sg13g2_decap_8 FILLER_107_381 ();
 sg13g2_fill_2 FILLER_107_388 ();
 sg13g2_fill_1 FILLER_107_390 ();
 sg13g2_decap_4 FILLER_107_396 ();
 sg13g2_fill_2 FILLER_107_400 ();
 sg13g2_decap_8 FILLER_107_437 ();
 sg13g2_decap_8 FILLER_107_444 ();
 sg13g2_decap_8 FILLER_107_451 ();
 sg13g2_decap_4 FILLER_107_458 ();
 sg13g2_fill_1 FILLER_107_488 ();
 sg13g2_decap_8 FILLER_107_514 ();
 sg13g2_fill_2 FILLER_107_641 ();
 sg13g2_fill_1 FILLER_107_643 ();
 sg13g2_fill_1 FILLER_107_670 ();
 sg13g2_fill_2 FILLER_107_685 ();
 sg13g2_fill_1 FILLER_107_687 ();
 sg13g2_decap_8 FILLER_107_692 ();
 sg13g2_fill_2 FILLER_107_699 ();
 sg13g2_fill_1 FILLER_107_701 ();
 sg13g2_decap_4 FILLER_107_754 ();
 sg13g2_fill_2 FILLER_107_758 ();
 sg13g2_decap_8 FILLER_107_786 ();
 sg13g2_fill_1 FILLER_107_793 ();
 sg13g2_decap_4 FILLER_107_798 ();
 sg13g2_fill_1 FILLER_107_802 ();
 sg13g2_fill_2 FILLER_107_808 ();
 sg13g2_fill_1 FILLER_107_810 ();
 sg13g2_decap_8 FILLER_107_820 ();
 sg13g2_fill_2 FILLER_107_841 ();
 sg13g2_decap_4 FILLER_107_849 ();
 sg13g2_fill_1 FILLER_107_853 ();
 sg13g2_fill_1 FILLER_107_863 ();
 sg13g2_decap_8 FILLER_107_873 ();
 sg13g2_decap_8 FILLER_107_880 ();
 sg13g2_fill_1 FILLER_107_918 ();
 sg13g2_decap_8 FILLER_107_932 ();
 sg13g2_decap_4 FILLER_107_939 ();
 sg13g2_fill_2 FILLER_107_943 ();
 sg13g2_fill_2 FILLER_107_985 ();
 sg13g2_fill_1 FILLER_107_987 ();
 sg13g2_decap_4 FILLER_107_1046 ();
 sg13g2_decap_8 FILLER_107_1082 ();
 sg13g2_decap_8 FILLER_107_1089 ();
 sg13g2_decap_8 FILLER_107_1096 ();
 sg13g2_decap_8 FILLER_107_1103 ();
 sg13g2_decap_8 FILLER_107_1110 ();
 sg13g2_decap_8 FILLER_107_1117 ();
 sg13g2_fill_1 FILLER_107_1139 ();
 sg13g2_decap_4 FILLER_107_1156 ();
 sg13g2_fill_2 FILLER_107_1160 ();
 sg13g2_decap_4 FILLER_107_1184 ();
 sg13g2_fill_2 FILLER_107_1188 ();
 sg13g2_fill_1 FILLER_107_1200 ();
 sg13g2_decap_8 FILLER_107_1206 ();
 sg13g2_fill_1 FILLER_107_1213 ();
 sg13g2_fill_1 FILLER_107_1240 ();
 sg13g2_decap_8 FILLER_107_1267 ();
 sg13g2_decap_4 FILLER_107_1300 ();
 sg13g2_fill_2 FILLER_107_1304 ();
 sg13g2_fill_1 FILLER_107_1316 ();
 sg13g2_decap_8 FILLER_107_1329 ();
 sg13g2_decap_8 FILLER_107_1336 ();
 sg13g2_fill_2 FILLER_107_1343 ();
 sg13g2_fill_1 FILLER_107_1345 ();
 sg13g2_fill_1 FILLER_107_1350 ();
 sg13g2_decap_8 FILLER_107_1355 ();
 sg13g2_decap_8 FILLER_107_1362 ();
 sg13g2_decap_4 FILLER_107_1369 ();
 sg13g2_fill_1 FILLER_107_1373 ();
 sg13g2_decap_8 FILLER_107_1400 ();
 sg13g2_decap_4 FILLER_107_1407 ();
 sg13g2_fill_1 FILLER_107_1411 ();
 sg13g2_decap_8 FILLER_107_1416 ();
 sg13g2_decap_8 FILLER_107_1423 ();
 sg13g2_decap_8 FILLER_107_1430 ();
 sg13g2_decap_8 FILLER_107_1437 ();
 sg13g2_decap_8 FILLER_107_1444 ();
 sg13g2_decap_8 FILLER_107_1451 ();
 sg13g2_decap_8 FILLER_107_1458 ();
 sg13g2_decap_8 FILLER_107_1465 ();
 sg13g2_decap_8 FILLER_107_1472 ();
 sg13g2_decap_8 FILLER_107_1479 ();
 sg13g2_decap_8 FILLER_107_1486 ();
 sg13g2_decap_8 FILLER_107_1493 ();
 sg13g2_decap_8 FILLER_107_1500 ();
 sg13g2_decap_8 FILLER_107_1507 ();
 sg13g2_decap_8 FILLER_107_1514 ();
 sg13g2_decap_8 FILLER_107_1521 ();
 sg13g2_decap_8 FILLER_107_1528 ();
 sg13g2_decap_8 FILLER_107_1535 ();
 sg13g2_decap_8 FILLER_107_1542 ();
 sg13g2_decap_8 FILLER_107_1549 ();
 sg13g2_decap_8 FILLER_107_1556 ();
 sg13g2_decap_8 FILLER_107_1563 ();
 sg13g2_decap_8 FILLER_107_1570 ();
 sg13g2_decap_8 FILLER_107_1577 ();
 sg13g2_decap_8 FILLER_107_1584 ();
 sg13g2_decap_8 FILLER_107_1591 ();
 sg13g2_decap_8 FILLER_107_1598 ();
 sg13g2_decap_8 FILLER_107_1605 ();
 sg13g2_decap_8 FILLER_107_1612 ();
 sg13g2_decap_4 FILLER_107_1619 ();
 sg13g2_fill_2 FILLER_107_1623 ();
 sg13g2_decap_8 FILLER_108_0 ();
 sg13g2_decap_8 FILLER_108_7 ();
 sg13g2_decap_8 FILLER_108_14 ();
 sg13g2_decap_8 FILLER_108_21 ();
 sg13g2_decap_8 FILLER_108_28 ();
 sg13g2_decap_8 FILLER_108_35 ();
 sg13g2_decap_8 FILLER_108_42 ();
 sg13g2_decap_8 FILLER_108_49 ();
 sg13g2_decap_8 FILLER_108_56 ();
 sg13g2_decap_8 FILLER_108_63 ();
 sg13g2_decap_8 FILLER_108_70 ();
 sg13g2_decap_8 FILLER_108_77 ();
 sg13g2_fill_1 FILLER_108_84 ();
 sg13g2_decap_4 FILLER_108_90 ();
 sg13g2_fill_1 FILLER_108_94 ();
 sg13g2_decap_8 FILLER_108_101 ();
 sg13g2_fill_1 FILLER_108_108 ();
 sg13g2_decap_8 FILLER_108_120 ();
 sg13g2_fill_2 FILLER_108_127 ();
 sg13g2_decap_8 FILLER_108_133 ();
 sg13g2_decap_4 FILLER_108_140 ();
 sg13g2_fill_2 FILLER_108_144 ();
 sg13g2_decap_8 FILLER_108_205 ();
 sg13g2_decap_8 FILLER_108_212 ();
 sg13g2_decap_8 FILLER_108_219 ();
 sg13g2_decap_8 FILLER_108_226 ();
 sg13g2_decap_4 FILLER_108_233 ();
 sg13g2_fill_1 FILLER_108_279 ();
 sg13g2_fill_1 FILLER_108_284 ();
 sg13g2_fill_2 FILLER_108_311 ();
 sg13g2_fill_1 FILLER_108_313 ();
 sg13g2_fill_2 FILLER_108_332 ();
 sg13g2_fill_2 FILLER_108_350 ();
 sg13g2_fill_2 FILLER_108_360 ();
 sg13g2_fill_1 FILLER_108_362 ();
 sg13g2_fill_2 FILLER_108_394 ();
 sg13g2_decap_8 FILLER_108_402 ();
 sg13g2_fill_1 FILLER_108_409 ();
 sg13g2_decap_4 FILLER_108_414 ();
 sg13g2_fill_1 FILLER_108_418 ();
 sg13g2_decap_4 FILLER_108_422 ();
 sg13g2_decap_8 FILLER_108_452 ();
 sg13g2_decap_4 FILLER_108_459 ();
 sg13g2_fill_2 FILLER_108_531 ();
 sg13g2_fill_2 FILLER_108_593 ();
 sg13g2_fill_1 FILLER_108_595 ();
 sg13g2_decap_4 FILLER_108_631 ();
 sg13g2_fill_2 FILLER_108_635 ();
 sg13g2_fill_1 FILLER_108_651 ();
 sg13g2_decap_4 FILLER_108_657 ();
 sg13g2_fill_1 FILLER_108_661 ();
 sg13g2_decap_4 FILLER_108_672 ();
 sg13g2_decap_8 FILLER_108_680 ();
 sg13g2_decap_8 FILLER_108_687 ();
 sg13g2_decap_8 FILLER_108_694 ();
 sg13g2_decap_4 FILLER_108_701 ();
 sg13g2_fill_1 FILLER_108_705 ();
 sg13g2_decap_8 FILLER_108_714 ();
 sg13g2_fill_2 FILLER_108_721 ();
 sg13g2_fill_1 FILLER_108_723 ();
 sg13g2_decap_4 FILLER_108_728 ();
 sg13g2_fill_2 FILLER_108_732 ();
 sg13g2_decap_4 FILLER_108_748 ();
 sg13g2_decap_8 FILLER_108_766 ();
 sg13g2_decap_8 FILLER_108_773 ();
 sg13g2_decap_8 FILLER_108_780 ();
 sg13g2_decap_4 FILLER_108_787 ();
 sg13g2_decap_4 FILLER_108_801 ();
 sg13g2_fill_2 FILLER_108_805 ();
 sg13g2_decap_8 FILLER_108_820 ();
 sg13g2_decap_4 FILLER_108_827 ();
 sg13g2_fill_2 FILLER_108_831 ();
 sg13g2_fill_1 FILLER_108_841 ();
 sg13g2_decap_4 FILLER_108_848 ();
 sg13g2_decap_8 FILLER_108_869 ();
 sg13g2_decap_8 FILLER_108_876 ();
 sg13g2_fill_1 FILLER_108_883 ();
 sg13g2_fill_1 FILLER_108_922 ();
 sg13g2_decap_8 FILLER_108_935 ();
 sg13g2_decap_8 FILLER_108_942 ();
 sg13g2_fill_2 FILLER_108_949 ();
 sg13g2_fill_1 FILLER_108_951 ();
 sg13g2_fill_2 FILLER_108_957 ();
 sg13g2_fill_1 FILLER_108_959 ();
 sg13g2_fill_1 FILLER_108_964 ();
 sg13g2_decap_4 FILLER_108_980 ();
 sg13g2_fill_2 FILLER_108_984 ();
 sg13g2_decap_8 FILLER_108_1012 ();
 sg13g2_fill_2 FILLER_108_1019 ();
 sg13g2_fill_1 FILLER_108_1021 ();
 sg13g2_decap_8 FILLER_108_1048 ();
 sg13g2_decap_8 FILLER_108_1055 ();
 sg13g2_decap_4 FILLER_108_1062 ();
 sg13g2_decap_8 FILLER_108_1071 ();
 sg13g2_decap_8 FILLER_108_1084 ();
 sg13g2_decap_8 FILLER_108_1091 ();
 sg13g2_decap_8 FILLER_108_1098 ();
 sg13g2_decap_8 FILLER_108_1105 ();
 sg13g2_decap_4 FILLER_108_1112 ();
 sg13g2_fill_1 FILLER_108_1116 ();
 sg13g2_decap_8 FILLER_108_1121 ();
 sg13g2_decap_8 FILLER_108_1128 ();
 sg13g2_decap_8 FILLER_108_1135 ();
 sg13g2_decap_8 FILLER_108_1142 ();
 sg13g2_decap_4 FILLER_108_1149 ();
 sg13g2_fill_2 FILLER_108_1153 ();
 sg13g2_decap_8 FILLER_108_1159 ();
 sg13g2_decap_8 FILLER_108_1166 ();
 sg13g2_decap_8 FILLER_108_1173 ();
 sg13g2_decap_8 FILLER_108_1180 ();
 sg13g2_decap_8 FILLER_108_1187 ();
 sg13g2_fill_2 FILLER_108_1194 ();
 sg13g2_decap_8 FILLER_108_1203 ();
 sg13g2_fill_2 FILLER_108_1210 ();
 sg13g2_fill_1 FILLER_108_1212 ();
 sg13g2_decap_8 FILLER_108_1217 ();
 sg13g2_decap_8 FILLER_108_1224 ();
 sg13g2_decap_8 FILLER_108_1231 ();
 sg13g2_decap_4 FILLER_108_1238 ();
 sg13g2_fill_2 FILLER_108_1242 ();
 sg13g2_decap_4 FILLER_108_1258 ();
 sg13g2_fill_2 FILLER_108_1262 ();
 sg13g2_decap_8 FILLER_108_1274 ();
 sg13g2_fill_1 FILLER_108_1281 ();
 sg13g2_decap_8 FILLER_108_1310 ();
 sg13g2_decap_8 FILLER_108_1317 ();
 sg13g2_decap_8 FILLER_108_1324 ();
 sg13g2_decap_4 FILLER_108_1331 ();
 sg13g2_fill_2 FILLER_108_1335 ();
 sg13g2_decap_8 FILLER_108_1345 ();
 sg13g2_decap_8 FILLER_108_1352 ();
 sg13g2_decap_8 FILLER_108_1359 ();
 sg13g2_decap_8 FILLER_108_1366 ();
 sg13g2_decap_8 FILLER_108_1373 ();
 sg13g2_fill_1 FILLER_108_1380 ();
 sg13g2_decap_4 FILLER_108_1385 ();
 sg13g2_decap_8 FILLER_108_1393 ();
 sg13g2_decap_8 FILLER_108_1400 ();
 sg13g2_decap_8 FILLER_108_1407 ();
 sg13g2_decap_8 FILLER_108_1414 ();
 sg13g2_decap_8 FILLER_108_1421 ();
 sg13g2_decap_8 FILLER_108_1428 ();
 sg13g2_decap_8 FILLER_108_1435 ();
 sg13g2_decap_8 FILLER_108_1442 ();
 sg13g2_decap_8 FILLER_108_1449 ();
 sg13g2_decap_8 FILLER_108_1456 ();
 sg13g2_decap_8 FILLER_108_1463 ();
 sg13g2_decap_8 FILLER_108_1470 ();
 sg13g2_decap_8 FILLER_108_1477 ();
 sg13g2_decap_8 FILLER_108_1484 ();
 sg13g2_decap_8 FILLER_108_1491 ();
 sg13g2_decap_8 FILLER_108_1498 ();
 sg13g2_decap_8 FILLER_108_1505 ();
 sg13g2_decap_8 FILLER_108_1512 ();
 sg13g2_decap_8 FILLER_108_1519 ();
 sg13g2_decap_8 FILLER_108_1526 ();
 sg13g2_decap_8 FILLER_108_1533 ();
 sg13g2_decap_8 FILLER_108_1540 ();
 sg13g2_decap_8 FILLER_108_1547 ();
 sg13g2_decap_8 FILLER_108_1554 ();
 sg13g2_decap_8 FILLER_108_1561 ();
 sg13g2_decap_8 FILLER_108_1568 ();
 sg13g2_decap_8 FILLER_108_1575 ();
 sg13g2_decap_8 FILLER_108_1582 ();
 sg13g2_decap_8 FILLER_108_1589 ();
 sg13g2_decap_8 FILLER_108_1596 ();
 sg13g2_decap_8 FILLER_108_1603 ();
 sg13g2_decap_8 FILLER_108_1610 ();
 sg13g2_decap_8 FILLER_108_1617 ();
 sg13g2_fill_1 FILLER_108_1624 ();
 sg13g2_decap_8 FILLER_109_0 ();
 sg13g2_decap_8 FILLER_109_7 ();
 sg13g2_decap_8 FILLER_109_14 ();
 sg13g2_decap_8 FILLER_109_21 ();
 sg13g2_decap_8 FILLER_109_28 ();
 sg13g2_decap_8 FILLER_109_35 ();
 sg13g2_decap_8 FILLER_109_42 ();
 sg13g2_decap_8 FILLER_109_49 ();
 sg13g2_fill_1 FILLER_109_56 ();
 sg13g2_decap_8 FILLER_109_61 ();
 sg13g2_fill_1 FILLER_109_68 ();
 sg13g2_decap_8 FILLER_109_74 ();
 sg13g2_fill_2 FILLER_109_81 ();
 sg13g2_fill_1 FILLER_109_83 ();
 sg13g2_decap_4 FILLER_109_92 ();
 sg13g2_fill_2 FILLER_109_96 ();
 sg13g2_fill_2 FILLER_109_106 ();
 sg13g2_fill_1 FILLER_109_114 ();
 sg13g2_fill_2 FILLER_109_119 ();
 sg13g2_fill_1 FILLER_109_152 ();
 sg13g2_decap_8 FILLER_109_157 ();
 sg13g2_fill_2 FILLER_109_164 ();
 sg13g2_decap_8 FILLER_109_170 ();
 sg13g2_decap_4 FILLER_109_182 ();
 sg13g2_fill_1 FILLER_109_186 ();
 sg13g2_decap_8 FILLER_109_191 ();
 sg13g2_fill_1 FILLER_109_198 ();
 sg13g2_decap_8 FILLER_109_209 ();
 sg13g2_fill_1 FILLER_109_216 ();
 sg13g2_fill_1 FILLER_109_247 ();
 sg13g2_fill_2 FILLER_109_274 ();
 sg13g2_fill_1 FILLER_109_276 ();
 sg13g2_fill_1 FILLER_109_293 ();
 sg13g2_decap_8 FILLER_109_361 ();
 sg13g2_decap_4 FILLER_109_368 ();
 sg13g2_fill_2 FILLER_109_372 ();
 sg13g2_decap_4 FILLER_109_378 ();
 sg13g2_decap_4 FILLER_109_386 ();
 sg13g2_fill_2 FILLER_109_395 ();
 sg13g2_fill_1 FILLER_109_402 ();
 sg13g2_decap_8 FILLER_109_458 ();
 sg13g2_fill_2 FILLER_109_465 ();
 sg13g2_decap_4 FILLER_109_493 ();
 sg13g2_fill_2 FILLER_109_497 ();
 sg13g2_decap_8 FILLER_109_503 ();
 sg13g2_decap_4 FILLER_109_510 ();
 sg13g2_fill_2 FILLER_109_514 ();
 sg13g2_decap_8 FILLER_109_568 ();
 sg13g2_fill_2 FILLER_109_575 ();
 sg13g2_fill_1 FILLER_109_577 ();
 sg13g2_decap_4 FILLER_109_639 ();
 sg13g2_decap_8 FILLER_109_647 ();
 sg13g2_decap_8 FILLER_109_659 ();
 sg13g2_decap_8 FILLER_109_666 ();
 sg13g2_decap_8 FILLER_109_673 ();
 sg13g2_fill_1 FILLER_109_680 ();
 sg13g2_decap_8 FILLER_109_709 ();
 sg13g2_decap_8 FILLER_109_716 ();
 sg13g2_fill_1 FILLER_109_723 ();
 sg13g2_fill_2 FILLER_109_728 ();
 sg13g2_fill_1 FILLER_109_730 ();
 sg13g2_decap_4 FILLER_109_738 ();
 sg13g2_decap_8 FILLER_109_752 ();
 sg13g2_fill_1 FILLER_109_759 ();
 sg13g2_decap_4 FILLER_109_764 ();
 sg13g2_fill_2 FILLER_109_768 ();
 sg13g2_fill_2 FILLER_109_801 ();
 sg13g2_decap_4 FILLER_109_807 ();
 sg13g2_fill_1 FILLER_109_811 ();
 sg13g2_decap_4 FILLER_109_827 ();
 sg13g2_fill_2 FILLER_109_831 ();
 sg13g2_fill_1 FILLER_109_840 ();
 sg13g2_fill_1 FILLER_109_845 ();
 sg13g2_fill_1 FILLER_109_854 ();
 sg13g2_fill_2 FILLER_109_863 ();
 sg13g2_decap_8 FILLER_109_869 ();
 sg13g2_fill_2 FILLER_109_876 ();
 sg13g2_fill_1 FILLER_109_878 ();
 sg13g2_decap_4 FILLER_109_905 ();
 sg13g2_decap_8 FILLER_109_913 ();
 sg13g2_decap_8 FILLER_109_920 ();
 sg13g2_fill_2 FILLER_109_927 ();
 sg13g2_fill_1 FILLER_109_929 ();
 sg13g2_decap_8 FILLER_109_938 ();
 sg13g2_fill_1 FILLER_109_945 ();
 sg13g2_fill_2 FILLER_109_960 ();
 sg13g2_decap_8 FILLER_109_974 ();
 sg13g2_decap_8 FILLER_109_989 ();
 sg13g2_fill_2 FILLER_109_996 ();
 sg13g2_fill_1 FILLER_109_998 ();
 sg13g2_decap_4 FILLER_109_1003 ();
 sg13g2_fill_2 FILLER_109_1007 ();
 sg13g2_decap_4 FILLER_109_1018 ();
 sg13g2_decap_8 FILLER_109_1031 ();
 sg13g2_decap_8 FILLER_109_1038 ();
 sg13g2_decap_4 FILLER_109_1045 ();
 sg13g2_fill_2 FILLER_109_1049 ();
 sg13g2_decap_8 FILLER_109_1068 ();
 sg13g2_fill_2 FILLER_109_1075 ();
 sg13g2_fill_1 FILLER_109_1077 ();
 sg13g2_decap_4 FILLER_109_1083 ();
 sg13g2_decap_8 FILLER_109_1101 ();
 sg13g2_fill_2 FILLER_109_1108 ();
 sg13g2_decap_8 FILLER_109_1136 ();
 sg13g2_decap_4 FILLER_109_1143 ();
 sg13g2_decap_8 FILLER_109_1173 ();
 sg13g2_fill_2 FILLER_109_1180 ();
 sg13g2_decap_8 FILLER_109_1186 ();
 sg13g2_decap_8 FILLER_109_1193 ();
 sg13g2_decap_4 FILLER_109_1200 ();
 sg13g2_fill_1 FILLER_109_1204 ();
 sg13g2_decap_8 FILLER_109_1231 ();
 sg13g2_decap_8 FILLER_109_1238 ();
 sg13g2_fill_1 FILLER_109_1245 ();
 sg13g2_fill_2 FILLER_109_1271 ();
 sg13g2_decap_8 FILLER_109_1289 ();
 sg13g2_decap_4 FILLER_109_1296 ();
 sg13g2_decap_4 FILLER_109_1304 ();
 sg13g2_fill_2 FILLER_109_1308 ();
 sg13g2_decap_8 FILLER_109_1314 ();
 sg13g2_decap_4 FILLER_109_1321 ();
 sg13g2_decap_8 FILLER_109_1349 ();
 sg13g2_decap_8 FILLER_109_1356 ();
 sg13g2_decap_8 FILLER_109_1363 ();
 sg13g2_decap_8 FILLER_109_1370 ();
 sg13g2_decap_8 FILLER_109_1377 ();
 sg13g2_decap_8 FILLER_109_1384 ();
 sg13g2_decap_8 FILLER_109_1391 ();
 sg13g2_decap_8 FILLER_109_1398 ();
 sg13g2_decap_8 FILLER_109_1405 ();
 sg13g2_decap_8 FILLER_109_1412 ();
 sg13g2_decap_8 FILLER_109_1419 ();
 sg13g2_decap_8 FILLER_109_1426 ();
 sg13g2_decap_8 FILLER_109_1433 ();
 sg13g2_decap_8 FILLER_109_1440 ();
 sg13g2_decap_8 FILLER_109_1447 ();
 sg13g2_decap_8 FILLER_109_1454 ();
 sg13g2_decap_8 FILLER_109_1461 ();
 sg13g2_decap_8 FILLER_109_1468 ();
 sg13g2_decap_8 FILLER_109_1475 ();
 sg13g2_decap_8 FILLER_109_1482 ();
 sg13g2_decap_8 FILLER_109_1489 ();
 sg13g2_decap_8 FILLER_109_1496 ();
 sg13g2_decap_8 FILLER_109_1503 ();
 sg13g2_decap_8 FILLER_109_1510 ();
 sg13g2_decap_8 FILLER_109_1517 ();
 sg13g2_decap_8 FILLER_109_1524 ();
 sg13g2_decap_8 FILLER_109_1531 ();
 sg13g2_decap_8 FILLER_109_1538 ();
 sg13g2_decap_8 FILLER_109_1545 ();
 sg13g2_decap_8 FILLER_109_1552 ();
 sg13g2_decap_8 FILLER_109_1559 ();
 sg13g2_decap_8 FILLER_109_1566 ();
 sg13g2_decap_8 FILLER_109_1573 ();
 sg13g2_decap_8 FILLER_109_1580 ();
 sg13g2_decap_8 FILLER_109_1587 ();
 sg13g2_decap_8 FILLER_109_1594 ();
 sg13g2_decap_8 FILLER_109_1601 ();
 sg13g2_decap_8 FILLER_109_1608 ();
 sg13g2_decap_8 FILLER_109_1615 ();
 sg13g2_fill_2 FILLER_109_1622 ();
 sg13g2_fill_1 FILLER_109_1624 ();
 sg13g2_decap_8 FILLER_110_0 ();
 sg13g2_decap_8 FILLER_110_7 ();
 sg13g2_decap_8 FILLER_110_14 ();
 sg13g2_decap_8 FILLER_110_21 ();
 sg13g2_decap_8 FILLER_110_28 ();
 sg13g2_decap_8 FILLER_110_35 ();
 sg13g2_decap_8 FILLER_110_42 ();
 sg13g2_fill_1 FILLER_110_49 ();
 sg13g2_fill_2 FILLER_110_76 ();
 sg13g2_fill_1 FILLER_110_78 ();
 sg13g2_decap_8 FILLER_110_109 ();
 sg13g2_decap_8 FILLER_110_116 ();
 sg13g2_fill_2 FILLER_110_160 ();
 sg13g2_fill_1 FILLER_110_162 ();
 sg13g2_decap_8 FILLER_110_167 ();
 sg13g2_decap_4 FILLER_110_174 ();
 sg13g2_fill_2 FILLER_110_178 ();
 sg13g2_decap_8 FILLER_110_206 ();
 sg13g2_decap_8 FILLER_110_239 ();
 sg13g2_decap_4 FILLER_110_246 ();
 sg13g2_fill_2 FILLER_110_250 ();
 sg13g2_decap_4 FILLER_110_259 ();
 sg13g2_fill_2 FILLER_110_263 ();
 sg13g2_fill_2 FILLER_110_269 ();
 sg13g2_decap_4 FILLER_110_275 ();
 sg13g2_fill_1 FILLER_110_279 ();
 sg13g2_fill_2 FILLER_110_306 ();
 sg13g2_fill_2 FILLER_110_313 ();
 sg13g2_fill_2 FILLER_110_320 ();
 sg13g2_fill_2 FILLER_110_332 ();
 sg13g2_decap_8 FILLER_110_354 ();
 sg13g2_decap_4 FILLER_110_361 ();
 sg13g2_fill_2 FILLER_110_365 ();
 sg13g2_fill_1 FILLER_110_403 ();
 sg13g2_decap_4 FILLER_110_409 ();
 sg13g2_fill_1 FILLER_110_413 ();
 sg13g2_decap_8 FILLER_110_432 ();
 sg13g2_fill_1 FILLER_110_439 ();
 sg13g2_fill_1 FILLER_110_472 ();
 sg13g2_decap_4 FILLER_110_479 ();
 sg13g2_fill_1 FILLER_110_483 ();
 sg13g2_decap_4 FILLER_110_509 ();
 sg13g2_fill_1 FILLER_110_513 ();
 sg13g2_decap_8 FILLER_110_557 ();
 sg13g2_fill_2 FILLER_110_564 ();
 sg13g2_fill_2 FILLER_110_621 ();
 sg13g2_fill_1 FILLER_110_623 ();
 sg13g2_fill_2 FILLER_110_634 ();
 sg13g2_decap_8 FILLER_110_662 ();
 sg13g2_fill_1 FILLER_110_669 ();
 sg13g2_decap_4 FILLER_110_675 ();
 sg13g2_fill_1 FILLER_110_679 ();
 sg13g2_decap_8 FILLER_110_705 ();
 sg13g2_decap_4 FILLER_110_712 ();
 sg13g2_fill_2 FILLER_110_742 ();
 sg13g2_decap_8 FILLER_110_809 ();
 sg13g2_decap_8 FILLER_110_816 ();
 sg13g2_decap_4 FILLER_110_823 ();
 sg13g2_decap_8 FILLER_110_848 ();
 sg13g2_decap_8 FILLER_110_855 ();
 sg13g2_fill_2 FILLER_110_862 ();
 sg13g2_decap_4 FILLER_110_874 ();
 sg13g2_decap_8 FILLER_110_883 ();
 sg13g2_fill_2 FILLER_110_890 ();
 sg13g2_decap_4 FILLER_110_897 ();
 sg13g2_decap_4 FILLER_110_927 ();
 sg13g2_fill_1 FILLER_110_948 ();
 sg13g2_decap_8 FILLER_110_957 ();
 sg13g2_fill_1 FILLER_110_977 ();
 sg13g2_decap_8 FILLER_110_983 ();
 sg13g2_fill_2 FILLER_110_990 ();
 sg13g2_decap_8 FILLER_110_1022 ();
 sg13g2_fill_1 FILLER_110_1029 ();
 sg13g2_decap_8 FILLER_110_1038 ();
 sg13g2_decap_4 FILLER_110_1045 ();
 sg13g2_decap_8 FILLER_110_1075 ();
 sg13g2_fill_2 FILLER_110_1114 ();
 sg13g2_fill_1 FILLER_110_1116 ();
 sg13g2_decap_8 FILLER_110_1122 ();
 sg13g2_decap_8 FILLER_110_1129 ();
 sg13g2_decap_4 FILLER_110_1136 ();
 sg13g2_fill_1 FILLER_110_1140 ();
 sg13g2_decap_8 FILLER_110_1151 ();
 sg13g2_decap_8 FILLER_110_1158 ();
 sg13g2_fill_1 FILLER_110_1165 ();
 sg13g2_decap_4 FILLER_110_1169 ();
 sg13g2_fill_2 FILLER_110_1173 ();
 sg13g2_decap_8 FILLER_110_1201 ();
 sg13g2_fill_1 FILLER_110_1208 ();
 sg13g2_decap_8 FILLER_110_1213 ();
 sg13g2_decap_4 FILLER_110_1220 ();
 sg13g2_fill_2 FILLER_110_1224 ();
 sg13g2_decap_4 FILLER_110_1246 ();
 sg13g2_fill_2 FILLER_110_1250 ();
 sg13g2_decap_8 FILLER_110_1256 ();
 sg13g2_decap_8 FILLER_110_1263 ();
 sg13g2_decap_4 FILLER_110_1270 ();
 sg13g2_fill_2 FILLER_110_1274 ();
 sg13g2_decap_4 FILLER_110_1280 ();
 sg13g2_fill_1 FILLER_110_1284 ();
 sg13g2_fill_2 FILLER_110_1289 ();
 sg13g2_fill_2 FILLER_110_1317 ();
 sg13g2_decap_8 FILLER_110_1339 ();
 sg13g2_decap_8 FILLER_110_1346 ();
 sg13g2_decap_8 FILLER_110_1353 ();
 sg13g2_decap_8 FILLER_110_1360 ();
 sg13g2_decap_8 FILLER_110_1367 ();
 sg13g2_decap_8 FILLER_110_1374 ();
 sg13g2_decap_8 FILLER_110_1381 ();
 sg13g2_decap_8 FILLER_110_1388 ();
 sg13g2_decap_8 FILLER_110_1395 ();
 sg13g2_decap_8 FILLER_110_1402 ();
 sg13g2_decap_8 FILLER_110_1409 ();
 sg13g2_decap_8 FILLER_110_1416 ();
 sg13g2_decap_8 FILLER_110_1423 ();
 sg13g2_decap_8 FILLER_110_1430 ();
 sg13g2_decap_8 FILLER_110_1437 ();
 sg13g2_decap_8 FILLER_110_1444 ();
 sg13g2_decap_8 FILLER_110_1451 ();
 sg13g2_decap_8 FILLER_110_1458 ();
 sg13g2_decap_8 FILLER_110_1465 ();
 sg13g2_decap_8 FILLER_110_1472 ();
 sg13g2_decap_8 FILLER_110_1479 ();
 sg13g2_decap_8 FILLER_110_1486 ();
 sg13g2_decap_8 FILLER_110_1493 ();
 sg13g2_decap_8 FILLER_110_1500 ();
 sg13g2_decap_8 FILLER_110_1507 ();
 sg13g2_decap_8 FILLER_110_1514 ();
 sg13g2_decap_8 FILLER_110_1521 ();
 sg13g2_decap_8 FILLER_110_1528 ();
 sg13g2_decap_8 FILLER_110_1535 ();
 sg13g2_decap_8 FILLER_110_1542 ();
 sg13g2_decap_8 FILLER_110_1549 ();
 sg13g2_decap_8 FILLER_110_1556 ();
 sg13g2_decap_8 FILLER_110_1563 ();
 sg13g2_decap_8 FILLER_110_1570 ();
 sg13g2_decap_8 FILLER_110_1577 ();
 sg13g2_decap_8 FILLER_110_1584 ();
 sg13g2_decap_8 FILLER_110_1591 ();
 sg13g2_decap_8 FILLER_110_1598 ();
 sg13g2_decap_8 FILLER_110_1605 ();
 sg13g2_decap_8 FILLER_110_1612 ();
 sg13g2_decap_4 FILLER_110_1619 ();
 sg13g2_fill_2 FILLER_110_1623 ();
 sg13g2_decap_8 FILLER_111_0 ();
 sg13g2_decap_8 FILLER_111_7 ();
 sg13g2_decap_8 FILLER_111_14 ();
 sg13g2_decap_8 FILLER_111_21 ();
 sg13g2_decap_8 FILLER_111_28 ();
 sg13g2_decap_8 FILLER_111_35 ();
 sg13g2_decap_8 FILLER_111_42 ();
 sg13g2_decap_8 FILLER_111_49 ();
 sg13g2_decap_8 FILLER_111_56 ();
 sg13g2_decap_4 FILLER_111_63 ();
 sg13g2_fill_2 FILLER_111_67 ();
 sg13g2_fill_2 FILLER_111_88 ();
 sg13g2_decap_8 FILLER_111_94 ();
 sg13g2_decap_8 FILLER_111_101 ();
 sg13g2_decap_8 FILLER_111_108 ();
 sg13g2_decap_4 FILLER_111_150 ();
 sg13g2_fill_2 FILLER_111_154 ();
 sg13g2_decap_8 FILLER_111_182 ();
 sg13g2_decap_8 FILLER_111_189 ();
 sg13g2_fill_2 FILLER_111_196 ();
 sg13g2_fill_1 FILLER_111_198 ();
 sg13g2_decap_8 FILLER_111_209 ();
 sg13g2_fill_2 FILLER_111_281 ();
 sg13g2_fill_2 FILLER_111_324 ();
 sg13g2_fill_2 FILLER_111_337 ();
 sg13g2_decap_8 FILLER_111_365 ();
 sg13g2_decap_8 FILLER_111_372 ();
 sg13g2_fill_1 FILLER_111_379 ();
 sg13g2_fill_2 FILLER_111_394 ();
 sg13g2_fill_1 FILLER_111_396 ();
 sg13g2_fill_2 FILLER_111_422 ();
 sg13g2_fill_1 FILLER_111_424 ();
 sg13g2_decap_4 FILLER_111_435 ();
 sg13g2_decap_8 FILLER_111_453 ();
 sg13g2_fill_1 FILLER_111_460 ();
 sg13g2_fill_1 FILLER_111_467 ();
 sg13g2_fill_2 FILLER_111_477 ();
 sg13g2_decap_4 FILLER_111_487 ();
 sg13g2_decap_8 FILLER_111_517 ();
 sg13g2_decap_4 FILLER_111_550 ();
 sg13g2_fill_1 FILLER_111_554 ();
 sg13g2_decap_4 FILLER_111_624 ();
 sg13g2_decap_8 FILLER_111_638 ();
 sg13g2_decap_4 FILLER_111_645 ();
 sg13g2_decap_8 FILLER_111_658 ();
 sg13g2_decap_8 FILLER_111_665 ();
 sg13g2_decap_8 FILLER_111_672 ();
 sg13g2_fill_2 FILLER_111_679 ();
 sg13g2_fill_1 FILLER_111_681 ();
 sg13g2_fill_1 FILLER_111_686 ();
 sg13g2_fill_1 FILLER_111_692 ();
 sg13g2_fill_1 FILLER_111_706 ();
 sg13g2_decap_8 FILLER_111_720 ();
 sg13g2_decap_4 FILLER_111_727 ();
 sg13g2_fill_1 FILLER_111_731 ();
 sg13g2_fill_2 FILLER_111_737 ();
 sg13g2_fill_2 FILLER_111_744 ();
 sg13g2_fill_1 FILLER_111_746 ();
 sg13g2_decap_8 FILLER_111_752 ();
 sg13g2_decap_8 FILLER_111_759 ();
 sg13g2_decap_8 FILLER_111_766 ();
 sg13g2_fill_2 FILLER_111_773 ();
 sg13g2_decap_8 FILLER_111_815 ();
 sg13g2_decap_8 FILLER_111_827 ();
 sg13g2_fill_2 FILLER_111_834 ();
 sg13g2_decap_8 FILLER_111_840 ();
 sg13g2_decap_8 FILLER_111_847 ();
 sg13g2_decap_8 FILLER_111_854 ();
 sg13g2_decap_8 FILLER_111_861 ();
 sg13g2_decap_8 FILLER_111_868 ();
 sg13g2_fill_1 FILLER_111_875 ();
 sg13g2_decap_4 FILLER_111_890 ();
 sg13g2_fill_2 FILLER_111_903 ();
 sg13g2_fill_2 FILLER_111_934 ();
 sg13g2_fill_2 FILLER_111_941 ();
 sg13g2_decap_8 FILLER_111_952 ();
 sg13g2_decap_8 FILLER_111_959 ();
 sg13g2_fill_2 FILLER_111_966 ();
 sg13g2_decap_8 FILLER_111_988 ();
 sg13g2_decap_8 FILLER_111_995 ();
 sg13g2_decap_4 FILLER_111_1002 ();
 sg13g2_fill_2 FILLER_111_1006 ();
 sg13g2_decap_8 FILLER_111_1013 ();
 sg13g2_fill_1 FILLER_111_1020 ();
 sg13g2_decap_8 FILLER_111_1064 ();
 sg13g2_decap_8 FILLER_111_1071 ();
 sg13g2_decap_4 FILLER_111_1078 ();
 sg13g2_decap_8 FILLER_111_1092 ();
 sg13g2_decap_8 FILLER_111_1099 ();
 sg13g2_decap_4 FILLER_111_1106 ();
 sg13g2_fill_2 FILLER_111_1110 ();
 sg13g2_decap_4 FILLER_111_1116 ();
 sg13g2_fill_1 FILLER_111_1120 ();
 sg13g2_fill_1 FILLER_111_1134 ();
 sg13g2_decap_8 FILLER_111_1149 ();
 sg13g2_decap_4 FILLER_111_1156 ();
 sg13g2_fill_2 FILLER_111_1196 ();
 sg13g2_fill_1 FILLER_111_1198 ();
 sg13g2_decap_8 FILLER_111_1271 ();
 sg13g2_decap_8 FILLER_111_1278 ();
 sg13g2_decap_4 FILLER_111_1285 ();
 sg13g2_fill_1 FILLER_111_1294 ();
 sg13g2_decap_4 FILLER_111_1303 ();
 sg13g2_fill_2 FILLER_111_1317 ();
 sg13g2_decap_8 FILLER_111_1324 ();
 sg13g2_decap_8 FILLER_111_1331 ();
 sg13g2_decap_8 FILLER_111_1338 ();
 sg13g2_decap_8 FILLER_111_1345 ();
 sg13g2_decap_8 FILLER_111_1352 ();
 sg13g2_decap_8 FILLER_111_1359 ();
 sg13g2_decap_8 FILLER_111_1366 ();
 sg13g2_decap_8 FILLER_111_1373 ();
 sg13g2_decap_8 FILLER_111_1380 ();
 sg13g2_decap_8 FILLER_111_1387 ();
 sg13g2_decap_8 FILLER_111_1394 ();
 sg13g2_decap_8 FILLER_111_1401 ();
 sg13g2_decap_8 FILLER_111_1408 ();
 sg13g2_decap_8 FILLER_111_1415 ();
 sg13g2_decap_8 FILLER_111_1422 ();
 sg13g2_decap_8 FILLER_111_1429 ();
 sg13g2_decap_8 FILLER_111_1436 ();
 sg13g2_decap_8 FILLER_111_1443 ();
 sg13g2_decap_8 FILLER_111_1450 ();
 sg13g2_decap_8 FILLER_111_1457 ();
 sg13g2_decap_8 FILLER_111_1464 ();
 sg13g2_decap_8 FILLER_111_1471 ();
 sg13g2_decap_8 FILLER_111_1478 ();
 sg13g2_decap_8 FILLER_111_1485 ();
 sg13g2_decap_8 FILLER_111_1492 ();
 sg13g2_decap_8 FILLER_111_1499 ();
 sg13g2_decap_8 FILLER_111_1506 ();
 sg13g2_decap_8 FILLER_111_1513 ();
 sg13g2_decap_8 FILLER_111_1520 ();
 sg13g2_decap_8 FILLER_111_1527 ();
 sg13g2_decap_8 FILLER_111_1534 ();
 sg13g2_decap_8 FILLER_111_1541 ();
 sg13g2_decap_8 FILLER_111_1548 ();
 sg13g2_decap_8 FILLER_111_1555 ();
 sg13g2_decap_8 FILLER_111_1562 ();
 sg13g2_decap_8 FILLER_111_1569 ();
 sg13g2_decap_8 FILLER_111_1576 ();
 sg13g2_decap_8 FILLER_111_1583 ();
 sg13g2_decap_8 FILLER_111_1590 ();
 sg13g2_decap_8 FILLER_111_1597 ();
 sg13g2_decap_8 FILLER_111_1604 ();
 sg13g2_decap_8 FILLER_111_1611 ();
 sg13g2_decap_8 FILLER_111_1618 ();
 sg13g2_decap_8 FILLER_112_0 ();
 sg13g2_decap_8 FILLER_112_7 ();
 sg13g2_decap_8 FILLER_112_14 ();
 sg13g2_decap_8 FILLER_112_21 ();
 sg13g2_decap_8 FILLER_112_28 ();
 sg13g2_decap_8 FILLER_112_35 ();
 sg13g2_decap_8 FILLER_112_42 ();
 sg13g2_decap_4 FILLER_112_49 ();
 sg13g2_fill_2 FILLER_112_82 ();
 sg13g2_fill_2 FILLER_112_93 ();
 sg13g2_decap_8 FILLER_112_99 ();
 sg13g2_decap_8 FILLER_112_106 ();
 sg13g2_decap_4 FILLER_112_113 ();
 sg13g2_decap_4 FILLER_112_122 ();
 sg13g2_decap_8 FILLER_112_133 ();
 sg13g2_decap_8 FILLER_112_140 ();
 sg13g2_decap_4 FILLER_112_147 ();
 sg13g2_fill_2 FILLER_112_185 ();
 sg13g2_fill_1 FILLER_112_187 ();
 sg13g2_fill_1 FILLER_112_192 ();
 sg13g2_fill_2 FILLER_112_218 ();
 sg13g2_decap_4 FILLER_112_224 ();
 sg13g2_fill_2 FILLER_112_253 ();
 sg13g2_fill_1 FILLER_112_255 ();
 sg13g2_decap_4 FILLER_112_282 ();
 sg13g2_fill_1 FILLER_112_286 ();
 sg13g2_fill_1 FILLER_112_313 ();
 sg13g2_fill_1 FILLER_112_319 ();
 sg13g2_decap_4 FILLER_112_326 ();
 sg13g2_decap_8 FILLER_112_336 ();
 sg13g2_fill_2 FILLER_112_343 ();
 sg13g2_fill_1 FILLER_112_345 ();
 sg13g2_fill_1 FILLER_112_350 ();
 sg13g2_fill_2 FILLER_112_376 ();
 sg13g2_fill_1 FILLER_112_378 ();
 sg13g2_fill_1 FILLER_112_431 ();
 sg13g2_decap_8 FILLER_112_450 ();
 sg13g2_fill_2 FILLER_112_457 ();
 sg13g2_fill_1 FILLER_112_459 ();
 sg13g2_fill_1 FILLER_112_464 ();
 sg13g2_fill_2 FILLER_112_469 ();
 sg13g2_fill_2 FILLER_112_476 ();
 sg13g2_fill_2 FILLER_112_483 ();
 sg13g2_decap_8 FILLER_112_489 ();
 sg13g2_decap_8 FILLER_112_496 ();
 sg13g2_decap_8 FILLER_112_503 ();
 sg13g2_decap_8 FILLER_112_510 ();
 sg13g2_decap_8 FILLER_112_517 ();
 sg13g2_decap_8 FILLER_112_524 ();
 sg13g2_fill_1 FILLER_112_531 ();
 sg13g2_decap_4 FILLER_112_535 ();
 sg13g2_decap_8 FILLER_112_543 ();
 sg13g2_decap_8 FILLER_112_550 ();
 sg13g2_decap_4 FILLER_112_557 ();
 sg13g2_fill_1 FILLER_112_561 ();
 sg13g2_decap_4 FILLER_112_602 ();
 sg13g2_fill_2 FILLER_112_606 ();
 sg13g2_decap_8 FILLER_112_631 ();
 sg13g2_decap_8 FILLER_112_638 ();
 sg13g2_decap_8 FILLER_112_645 ();
 sg13g2_decap_8 FILLER_112_652 ();
 sg13g2_fill_2 FILLER_112_659 ();
 sg13g2_decap_8 FILLER_112_665 ();
 sg13g2_fill_1 FILLER_112_672 ();
 sg13g2_fill_1 FILLER_112_685 ();
 sg13g2_decap_8 FILLER_112_691 ();
 sg13g2_decap_8 FILLER_112_698 ();
 sg13g2_decap_8 FILLER_112_705 ();
 sg13g2_decap_8 FILLER_112_712 ();
 sg13g2_decap_8 FILLER_112_719 ();
 sg13g2_decap_8 FILLER_112_726 ();
 sg13g2_fill_2 FILLER_112_733 ();
 sg13g2_fill_1 FILLER_112_735 ();
 sg13g2_decap_8 FILLER_112_740 ();
 sg13g2_decap_4 FILLER_112_747 ();
 sg13g2_fill_1 FILLER_112_751 ();
 sg13g2_decap_8 FILLER_112_756 ();
 sg13g2_decap_8 FILLER_112_763 ();
 sg13g2_decap_8 FILLER_112_770 ();
 sg13g2_decap_8 FILLER_112_794 ();
 sg13g2_decap_8 FILLER_112_801 ();
 sg13g2_decap_8 FILLER_112_812 ();
 sg13g2_fill_1 FILLER_112_819 ();
 sg13g2_decap_8 FILLER_112_855 ();
 sg13g2_decap_8 FILLER_112_862 ();
 sg13g2_decap_8 FILLER_112_869 ();
 sg13g2_decap_8 FILLER_112_876 ();
 sg13g2_fill_2 FILLER_112_883 ();
 sg13g2_decap_8 FILLER_112_894 ();
 sg13g2_fill_2 FILLER_112_901 ();
 sg13g2_fill_1 FILLER_112_903 ();
 sg13g2_decap_4 FILLER_112_934 ();
 sg13g2_decap_8 FILLER_112_958 ();
 sg13g2_fill_1 FILLER_112_965 ();
 sg13g2_decap_4 FILLER_112_976 ();
 sg13g2_fill_1 FILLER_112_980 ();
 sg13g2_decap_8 FILLER_112_986 ();
 sg13g2_decap_8 FILLER_112_993 ();
 sg13g2_decap_8 FILLER_112_1000 ();
 sg13g2_decap_4 FILLER_112_1007 ();
 sg13g2_fill_2 FILLER_112_1050 ();
 sg13g2_fill_1 FILLER_112_1052 ();
 sg13g2_fill_2 FILLER_112_1078 ();
 sg13g2_fill_1 FILLER_112_1080 ();
 sg13g2_decap_8 FILLER_112_1091 ();
 sg13g2_decap_8 FILLER_112_1098 ();
 sg13g2_fill_2 FILLER_112_1105 ();
 sg13g2_fill_1 FILLER_112_1115 ();
 sg13g2_fill_1 FILLER_112_1125 ();
 sg13g2_fill_1 FILLER_112_1139 ();
 sg13g2_decap_4 FILLER_112_1145 ();
 sg13g2_fill_1 FILLER_112_1149 ();
 sg13g2_fill_2 FILLER_112_1171 ();
 sg13g2_decap_8 FILLER_112_1177 ();
 sg13g2_decap_4 FILLER_112_1184 ();
 sg13g2_fill_2 FILLER_112_1188 ();
 sg13g2_decap_8 FILLER_112_1226 ();
 sg13g2_decap_8 FILLER_112_1233 ();
 sg13g2_fill_2 FILLER_112_1240 ();
 sg13g2_fill_1 FILLER_112_1242 ();
 sg13g2_decap_4 FILLER_112_1276 ();
 sg13g2_fill_2 FILLER_112_1280 ();
 sg13g2_decap_8 FILLER_112_1291 ();
 sg13g2_fill_1 FILLER_112_1298 ();
 sg13g2_decap_8 FILLER_112_1328 ();
 sg13g2_decap_8 FILLER_112_1335 ();
 sg13g2_fill_1 FILLER_112_1342 ();
 sg13g2_decap_8 FILLER_112_1347 ();
 sg13g2_decap_8 FILLER_112_1354 ();
 sg13g2_decap_8 FILLER_112_1361 ();
 sg13g2_decap_8 FILLER_112_1368 ();
 sg13g2_decap_8 FILLER_112_1375 ();
 sg13g2_decap_8 FILLER_112_1382 ();
 sg13g2_decap_8 FILLER_112_1389 ();
 sg13g2_decap_8 FILLER_112_1396 ();
 sg13g2_decap_8 FILLER_112_1403 ();
 sg13g2_decap_8 FILLER_112_1410 ();
 sg13g2_decap_8 FILLER_112_1417 ();
 sg13g2_decap_8 FILLER_112_1424 ();
 sg13g2_decap_8 FILLER_112_1431 ();
 sg13g2_decap_8 FILLER_112_1438 ();
 sg13g2_decap_8 FILLER_112_1445 ();
 sg13g2_decap_8 FILLER_112_1452 ();
 sg13g2_decap_8 FILLER_112_1459 ();
 sg13g2_decap_8 FILLER_112_1466 ();
 sg13g2_decap_8 FILLER_112_1473 ();
 sg13g2_decap_8 FILLER_112_1480 ();
 sg13g2_decap_8 FILLER_112_1487 ();
 sg13g2_decap_8 FILLER_112_1494 ();
 sg13g2_decap_8 FILLER_112_1501 ();
 sg13g2_decap_8 FILLER_112_1508 ();
 sg13g2_decap_8 FILLER_112_1515 ();
 sg13g2_decap_8 FILLER_112_1522 ();
 sg13g2_decap_8 FILLER_112_1529 ();
 sg13g2_decap_8 FILLER_112_1536 ();
 sg13g2_decap_8 FILLER_112_1543 ();
 sg13g2_decap_8 FILLER_112_1550 ();
 sg13g2_decap_8 FILLER_112_1557 ();
 sg13g2_decap_8 FILLER_112_1564 ();
 sg13g2_decap_8 FILLER_112_1571 ();
 sg13g2_decap_8 FILLER_112_1578 ();
 sg13g2_decap_8 FILLER_112_1585 ();
 sg13g2_decap_8 FILLER_112_1592 ();
 sg13g2_decap_8 FILLER_112_1599 ();
 sg13g2_decap_8 FILLER_112_1606 ();
 sg13g2_decap_8 FILLER_112_1613 ();
 sg13g2_decap_4 FILLER_112_1620 ();
 sg13g2_fill_1 FILLER_112_1624 ();
 sg13g2_decap_8 FILLER_113_0 ();
 sg13g2_decap_8 FILLER_113_7 ();
 sg13g2_decap_8 FILLER_113_14 ();
 sg13g2_decap_8 FILLER_113_21 ();
 sg13g2_decap_8 FILLER_113_28 ();
 sg13g2_decap_8 FILLER_113_35 ();
 sg13g2_decap_8 FILLER_113_42 ();
 sg13g2_decap_4 FILLER_113_49 ();
 sg13g2_fill_1 FILLER_113_53 ();
 sg13g2_fill_2 FILLER_113_80 ();
 sg13g2_decap_4 FILLER_113_113 ();
 sg13g2_fill_1 FILLER_113_117 ();
 sg13g2_decap_8 FILLER_113_122 ();
 sg13g2_decap_8 FILLER_113_129 ();
 sg13g2_decap_8 FILLER_113_136 ();
 sg13g2_decap_8 FILLER_113_143 ();
 sg13g2_decap_4 FILLER_113_150 ();
 sg13g2_fill_1 FILLER_113_154 ();
 sg13g2_fill_2 FILLER_113_212 ();
 sg13g2_fill_1 FILLER_113_214 ();
 sg13g2_decap_4 FILLER_113_275 ();
 sg13g2_fill_1 FILLER_113_279 ();
 sg13g2_decap_4 FILLER_113_284 ();
 sg13g2_fill_1 FILLER_113_288 ();
 sg13g2_fill_2 FILLER_113_310 ();
 sg13g2_fill_1 FILLER_113_312 ();
 sg13g2_fill_1 FILLER_113_323 ();
 sg13g2_decap_8 FILLER_113_330 ();
 sg13g2_decap_8 FILLER_113_337 ();
 sg13g2_decap_8 FILLER_113_344 ();
 sg13g2_decap_8 FILLER_113_384 ();
 sg13g2_fill_2 FILLER_113_391 ();
 sg13g2_fill_1 FILLER_113_393 ();
 sg13g2_decap_8 FILLER_113_404 ();
 sg13g2_decap_4 FILLER_113_411 ();
 sg13g2_fill_1 FILLER_113_415 ();
 sg13g2_decap_8 FILLER_113_420 ();
 sg13g2_fill_1 FILLER_113_427 ();
 sg13g2_fill_1 FILLER_113_444 ();
 sg13g2_decap_8 FILLER_113_455 ();
 sg13g2_decap_4 FILLER_113_462 ();
 sg13g2_fill_2 FILLER_113_466 ();
 sg13g2_decap_4 FILLER_113_472 ();
 sg13g2_fill_2 FILLER_113_486 ();
 sg13g2_decap_8 FILLER_113_493 ();
 sg13g2_decap_8 FILLER_113_500 ();
 sg13g2_decap_4 FILLER_113_507 ();
 sg13g2_fill_1 FILLER_113_511 ();
 sg13g2_decap_8 FILLER_113_516 ();
 sg13g2_decap_4 FILLER_113_523 ();
 sg13g2_fill_1 FILLER_113_527 ();
 sg13g2_decap_8 FILLER_113_557 ();
 sg13g2_fill_2 FILLER_113_564 ();
 sg13g2_decap_8 FILLER_113_571 ();
 sg13g2_decap_8 FILLER_113_578 ();
 sg13g2_decap_8 FILLER_113_585 ();
 sg13g2_decap_8 FILLER_113_592 ();
 sg13g2_decap_8 FILLER_113_599 ();
 sg13g2_fill_2 FILLER_113_606 ();
 sg13g2_fill_2 FILLER_113_613 ();
 sg13g2_decap_8 FILLER_113_619 ();
 sg13g2_fill_2 FILLER_113_626 ();
 sg13g2_fill_1 FILLER_113_628 ();
 sg13g2_fill_2 FILLER_113_647 ();
 sg13g2_fill_1 FILLER_113_649 ();
 sg13g2_decap_8 FILLER_113_655 ();
 sg13g2_decap_4 FILLER_113_662 ();
 sg13g2_fill_1 FILLER_113_666 ();
 sg13g2_decap_8 FILLER_113_675 ();
 sg13g2_fill_2 FILLER_113_708 ();
 sg13g2_decap_8 FILLER_113_714 ();
 sg13g2_fill_1 FILLER_113_721 ();
 sg13g2_decap_8 FILLER_113_726 ();
 sg13g2_fill_2 FILLER_113_733 ();
 sg13g2_decap_8 FILLER_113_774 ();
 sg13g2_decap_8 FILLER_113_781 ();
 sg13g2_decap_4 FILLER_113_788 ();
 sg13g2_fill_2 FILLER_113_792 ();
 sg13g2_decap_8 FILLER_113_819 ();
 sg13g2_decap_8 FILLER_113_826 ();
 sg13g2_decap_8 FILLER_113_833 ();
 sg13g2_fill_2 FILLER_113_840 ();
 sg13g2_fill_1 FILLER_113_842 ();
 sg13g2_fill_2 FILLER_113_876 ();
 sg13g2_fill_1 FILLER_113_878 ();
 sg13g2_decap_8 FILLER_113_888 ();
 sg13g2_decap_8 FILLER_113_895 ();
 sg13g2_fill_2 FILLER_113_902 ();
 sg13g2_fill_1 FILLER_113_904 ();
 sg13g2_decap_8 FILLER_113_910 ();
 sg13g2_decap_8 FILLER_113_917 ();
 sg13g2_decap_8 FILLER_113_924 ();
 sg13g2_decap_8 FILLER_113_931 ();
 sg13g2_decap_8 FILLER_113_943 ();
 sg13g2_decap_8 FILLER_113_950 ();
 sg13g2_decap_8 FILLER_113_957 ();
 sg13g2_decap_4 FILLER_113_964 ();
 sg13g2_fill_2 FILLER_113_968 ();
 sg13g2_fill_2 FILLER_113_975 ();
 sg13g2_fill_1 FILLER_113_1073 ();
 sg13g2_fill_2 FILLER_113_1094 ();
 sg13g2_fill_1 FILLER_113_1096 ();
 sg13g2_decap_8 FILLER_113_1105 ();
 sg13g2_decap_8 FILLER_113_1120 ();
 sg13g2_decap_8 FILLER_113_1127 ();
 sg13g2_decap_8 FILLER_113_1134 ();
 sg13g2_decap_8 FILLER_113_1141 ();
 sg13g2_decap_8 FILLER_113_1148 ();
 sg13g2_decap_4 FILLER_113_1160 ();
 sg13g2_fill_2 FILLER_113_1164 ();
 sg13g2_decap_4 FILLER_113_1180 ();
 sg13g2_fill_2 FILLER_113_1184 ();
 sg13g2_fill_2 FILLER_113_1202 ();
 sg13g2_decap_8 FILLER_113_1209 ();
 sg13g2_decap_4 FILLER_113_1216 ();
 sg13g2_fill_2 FILLER_113_1220 ();
 sg13g2_fill_1 FILLER_113_1232 ();
 sg13g2_decap_4 FILLER_113_1300 ();
 sg13g2_fill_1 FILLER_113_1304 ();
 sg13g2_decap_8 FILLER_113_1365 ();
 sg13g2_decap_8 FILLER_113_1372 ();
 sg13g2_decap_8 FILLER_113_1379 ();
 sg13g2_decap_8 FILLER_113_1386 ();
 sg13g2_decap_8 FILLER_113_1393 ();
 sg13g2_decap_8 FILLER_113_1400 ();
 sg13g2_decap_8 FILLER_113_1407 ();
 sg13g2_decap_8 FILLER_113_1414 ();
 sg13g2_decap_8 FILLER_113_1421 ();
 sg13g2_decap_8 FILLER_113_1428 ();
 sg13g2_decap_8 FILLER_113_1435 ();
 sg13g2_decap_8 FILLER_113_1442 ();
 sg13g2_decap_8 FILLER_113_1449 ();
 sg13g2_decap_8 FILLER_113_1456 ();
 sg13g2_decap_8 FILLER_113_1463 ();
 sg13g2_decap_8 FILLER_113_1470 ();
 sg13g2_decap_8 FILLER_113_1477 ();
 sg13g2_decap_8 FILLER_113_1484 ();
 sg13g2_decap_8 FILLER_113_1491 ();
 sg13g2_decap_8 FILLER_113_1498 ();
 sg13g2_decap_8 FILLER_113_1505 ();
 sg13g2_decap_8 FILLER_113_1512 ();
 sg13g2_decap_8 FILLER_113_1519 ();
 sg13g2_decap_8 FILLER_113_1526 ();
 sg13g2_decap_8 FILLER_113_1533 ();
 sg13g2_decap_8 FILLER_113_1540 ();
 sg13g2_decap_8 FILLER_113_1547 ();
 sg13g2_decap_8 FILLER_113_1554 ();
 sg13g2_decap_8 FILLER_113_1561 ();
 sg13g2_decap_8 FILLER_113_1568 ();
 sg13g2_decap_8 FILLER_113_1575 ();
 sg13g2_decap_8 FILLER_113_1582 ();
 sg13g2_decap_8 FILLER_113_1589 ();
 sg13g2_decap_8 FILLER_113_1596 ();
 sg13g2_decap_8 FILLER_113_1603 ();
 sg13g2_decap_8 FILLER_113_1610 ();
 sg13g2_decap_8 FILLER_113_1617 ();
 sg13g2_fill_1 FILLER_113_1624 ();
 sg13g2_decap_8 FILLER_114_0 ();
 sg13g2_decap_8 FILLER_114_7 ();
 sg13g2_decap_8 FILLER_114_14 ();
 sg13g2_decap_8 FILLER_114_21 ();
 sg13g2_decap_8 FILLER_114_28 ();
 sg13g2_decap_8 FILLER_114_35 ();
 sg13g2_decap_8 FILLER_114_42 ();
 sg13g2_decap_8 FILLER_114_49 ();
 sg13g2_decap_8 FILLER_114_56 ();
 sg13g2_decap_8 FILLER_114_63 ();
 sg13g2_decap_4 FILLER_114_70 ();
 sg13g2_fill_1 FILLER_114_74 ();
 sg13g2_fill_1 FILLER_114_79 ();
 sg13g2_fill_2 FILLER_114_84 ();
 sg13g2_fill_1 FILLER_114_90 ();
 sg13g2_decap_4 FILLER_114_95 ();
 sg13g2_decap_8 FILLER_114_104 ();
 sg13g2_fill_1 FILLER_114_111 ();
 sg13g2_decap_4 FILLER_114_138 ();
 sg13g2_fill_1 FILLER_114_142 ();
 sg13g2_decap_4 FILLER_114_148 ();
 sg13g2_decap_8 FILLER_114_162 ();
 sg13g2_decap_8 FILLER_114_169 ();
 sg13g2_decap_8 FILLER_114_176 ();
 sg13g2_decap_8 FILLER_114_183 ();
 sg13g2_decap_8 FILLER_114_190 ();
 sg13g2_decap_8 FILLER_114_197 ();
 sg13g2_decap_4 FILLER_114_204 ();
 sg13g2_fill_2 FILLER_114_208 ();
 sg13g2_fill_2 FILLER_114_236 ();
 sg13g2_fill_1 FILLER_114_253 ();
 sg13g2_decap_8 FILLER_114_329 ();
 sg13g2_decap_8 FILLER_114_336 ();
 sg13g2_fill_2 FILLER_114_343 ();
 sg13g2_fill_1 FILLER_114_345 ();
 sg13g2_fill_2 FILLER_114_372 ();
 sg13g2_fill_1 FILLER_114_374 ();
 sg13g2_decap_4 FILLER_114_405 ();
 sg13g2_fill_2 FILLER_114_409 ();
 sg13g2_decap_8 FILLER_114_420 ();
 sg13g2_decap_8 FILLER_114_427 ();
 sg13g2_decap_8 FILLER_114_443 ();
 sg13g2_decap_8 FILLER_114_450 ();
 sg13g2_decap_8 FILLER_114_457 ();
 sg13g2_fill_2 FILLER_114_464 ();
 sg13g2_fill_1 FILLER_114_466 ();
 sg13g2_decap_8 FILLER_114_477 ();
 sg13g2_decap_8 FILLER_114_484 ();
 sg13g2_decap_8 FILLER_114_491 ();
 sg13g2_decap_4 FILLER_114_498 ();
 sg13g2_fill_2 FILLER_114_502 ();
 sg13g2_decap_8 FILLER_114_555 ();
 sg13g2_decap_4 FILLER_114_562 ();
 sg13g2_decap_8 FILLER_114_570 ();
 sg13g2_decap_8 FILLER_114_577 ();
 sg13g2_decap_8 FILLER_114_584 ();
 sg13g2_fill_1 FILLER_114_595 ();
 sg13g2_decap_4 FILLER_114_600 ();
 sg13g2_fill_1 FILLER_114_604 ();
 sg13g2_fill_2 FILLER_114_620 ();
 sg13g2_decap_4 FILLER_114_632 ();
 sg13g2_fill_2 FILLER_114_636 ();
 sg13g2_fill_1 FILLER_114_643 ();
 sg13g2_fill_2 FILLER_114_661 ();
 sg13g2_fill_2 FILLER_114_676 ();
 sg13g2_fill_1 FILLER_114_678 ();
 sg13g2_decap_4 FILLER_114_692 ();
 sg13g2_fill_1 FILLER_114_696 ();
 sg13g2_fill_1 FILLER_114_702 ();
 sg13g2_fill_2 FILLER_114_712 ();
 sg13g2_fill_1 FILLER_114_714 ();
 sg13g2_fill_2 FILLER_114_741 ();
 sg13g2_decap_8 FILLER_114_748 ();
 sg13g2_decap_8 FILLER_114_755 ();
 sg13g2_fill_1 FILLER_114_762 ();
 sg13g2_decap_4 FILLER_114_794 ();
 sg13g2_fill_1 FILLER_114_798 ();
 sg13g2_decap_8 FILLER_114_825 ();
 sg13g2_fill_2 FILLER_114_832 ();
 sg13g2_fill_1 FILLER_114_838 ();
 sg13g2_fill_2 FILLER_114_869 ();
 sg13g2_fill_1 FILLER_114_871 ();
 sg13g2_decap_8 FILLER_114_903 ();
 sg13g2_decap_8 FILLER_114_910 ();
 sg13g2_fill_1 FILLER_114_917 ();
 sg13g2_decap_8 FILLER_114_943 ();
 sg13g2_fill_2 FILLER_114_950 ();
 sg13g2_fill_1 FILLER_114_952 ();
 sg13g2_decap_8 FILLER_114_1008 ();
 sg13g2_fill_1 FILLER_114_1015 ();
 sg13g2_decap_8 FILLER_114_1021 ();
 sg13g2_decap_8 FILLER_114_1028 ();
 sg13g2_decap_4 FILLER_114_1035 ();
 sg13g2_decap_8 FILLER_114_1044 ();
 sg13g2_decap_8 FILLER_114_1055 ();
 sg13g2_decap_8 FILLER_114_1062 ();
 sg13g2_decap_4 FILLER_114_1069 ();
 sg13g2_fill_1 FILLER_114_1073 ();
 sg13g2_fill_1 FILLER_114_1087 ();
 sg13g2_fill_1 FILLER_114_1096 ();
 sg13g2_decap_4 FILLER_114_1105 ();
 sg13g2_decap_8 FILLER_114_1118 ();
 sg13g2_decap_8 FILLER_114_1125 ();
 sg13g2_decap_4 FILLER_114_1132 ();
 sg13g2_fill_2 FILLER_114_1136 ();
 sg13g2_fill_2 FILLER_114_1143 ();
 sg13g2_decap_8 FILLER_114_1157 ();
 sg13g2_decap_8 FILLER_114_1164 ();
 sg13g2_decap_8 FILLER_114_1171 ();
 sg13g2_fill_1 FILLER_114_1192 ();
 sg13g2_decap_8 FILLER_114_1197 ();
 sg13g2_decap_8 FILLER_114_1204 ();
 sg13g2_fill_2 FILLER_114_1211 ();
 sg13g2_fill_1 FILLER_114_1213 ();
 sg13g2_decap_8 FILLER_114_1227 ();
 sg13g2_decap_8 FILLER_114_1234 ();
 sg13g2_fill_1 FILLER_114_1241 ();
 sg13g2_decap_8 FILLER_114_1256 ();
 sg13g2_decap_8 FILLER_114_1263 ();
 sg13g2_decap_4 FILLER_114_1270 ();
 sg13g2_decap_8 FILLER_114_1278 ();
 sg13g2_decap_8 FILLER_114_1285 ();
 sg13g2_decap_8 FILLER_114_1292 ();
 sg13g2_decap_8 FILLER_114_1299 ();
 sg13g2_fill_2 FILLER_114_1310 ();
 sg13g2_decap_8 FILLER_114_1316 ();
 sg13g2_decap_8 FILLER_114_1323 ();
 sg13g2_fill_2 FILLER_114_1330 ();
 sg13g2_decap_8 FILLER_114_1336 ();
 sg13g2_decap_4 FILLER_114_1343 ();
 sg13g2_fill_1 FILLER_114_1347 ();
 sg13g2_decap_8 FILLER_114_1378 ();
 sg13g2_decap_8 FILLER_114_1385 ();
 sg13g2_decap_8 FILLER_114_1392 ();
 sg13g2_decap_8 FILLER_114_1399 ();
 sg13g2_decap_8 FILLER_114_1406 ();
 sg13g2_decap_8 FILLER_114_1413 ();
 sg13g2_decap_8 FILLER_114_1420 ();
 sg13g2_decap_8 FILLER_114_1427 ();
 sg13g2_decap_8 FILLER_114_1434 ();
 sg13g2_decap_8 FILLER_114_1441 ();
 sg13g2_decap_8 FILLER_114_1448 ();
 sg13g2_decap_8 FILLER_114_1455 ();
 sg13g2_decap_8 FILLER_114_1462 ();
 sg13g2_decap_8 FILLER_114_1469 ();
 sg13g2_decap_8 FILLER_114_1476 ();
 sg13g2_decap_8 FILLER_114_1483 ();
 sg13g2_decap_8 FILLER_114_1490 ();
 sg13g2_decap_8 FILLER_114_1497 ();
 sg13g2_decap_8 FILLER_114_1504 ();
 sg13g2_decap_8 FILLER_114_1511 ();
 sg13g2_decap_8 FILLER_114_1518 ();
 sg13g2_decap_8 FILLER_114_1525 ();
 sg13g2_decap_8 FILLER_114_1532 ();
 sg13g2_decap_8 FILLER_114_1539 ();
 sg13g2_decap_8 FILLER_114_1546 ();
 sg13g2_decap_8 FILLER_114_1553 ();
 sg13g2_decap_8 FILLER_114_1560 ();
 sg13g2_decap_8 FILLER_114_1567 ();
 sg13g2_decap_8 FILLER_114_1574 ();
 sg13g2_decap_8 FILLER_114_1581 ();
 sg13g2_decap_8 FILLER_114_1588 ();
 sg13g2_decap_8 FILLER_114_1595 ();
 sg13g2_decap_8 FILLER_114_1602 ();
 sg13g2_decap_8 FILLER_114_1609 ();
 sg13g2_decap_8 FILLER_114_1616 ();
 sg13g2_fill_2 FILLER_114_1623 ();
 sg13g2_decap_8 FILLER_115_0 ();
 sg13g2_decap_8 FILLER_115_7 ();
 sg13g2_decap_8 FILLER_115_14 ();
 sg13g2_decap_8 FILLER_115_21 ();
 sg13g2_decap_8 FILLER_115_28 ();
 sg13g2_decap_8 FILLER_115_35 ();
 sg13g2_decap_8 FILLER_115_42 ();
 sg13g2_decap_8 FILLER_115_49 ();
 sg13g2_decap_8 FILLER_115_56 ();
 sg13g2_decap_8 FILLER_115_63 ();
 sg13g2_fill_2 FILLER_115_70 ();
 sg13g2_fill_1 FILLER_115_72 ();
 sg13g2_fill_1 FILLER_115_104 ();
 sg13g2_fill_2 FILLER_115_110 ();
 sg13g2_decap_8 FILLER_115_119 ();
 sg13g2_fill_2 FILLER_115_126 ();
 sg13g2_fill_2 FILLER_115_143 ();
 sg13g2_fill_2 FILLER_115_157 ();
 sg13g2_decap_4 FILLER_115_164 ();
 sg13g2_fill_2 FILLER_115_168 ();
 sg13g2_decap_8 FILLER_115_175 ();
 sg13g2_decap_8 FILLER_115_182 ();
 sg13g2_fill_2 FILLER_115_189 ();
 sg13g2_decap_4 FILLER_115_195 ();
 sg13g2_fill_2 FILLER_115_226 ();
 sg13g2_fill_2 FILLER_115_271 ();
 sg13g2_fill_1 FILLER_115_309 ();
 sg13g2_fill_2 FILLER_115_320 ();
 sg13g2_decap_8 FILLER_115_339 ();
 sg13g2_decap_8 FILLER_115_346 ();
 sg13g2_decap_8 FILLER_115_353 ();
 sg13g2_decap_8 FILLER_115_360 ();
 sg13g2_fill_2 FILLER_115_367 ();
 sg13g2_fill_1 FILLER_115_369 ();
 sg13g2_fill_2 FILLER_115_385 ();
 sg13g2_fill_1 FILLER_115_387 ();
 sg13g2_fill_2 FILLER_115_419 ();
 sg13g2_fill_1 FILLER_115_421 ();
 sg13g2_fill_2 FILLER_115_427 ();
 sg13g2_decap_8 FILLER_115_455 ();
 sg13g2_decap_4 FILLER_115_462 ();
 sg13g2_fill_2 FILLER_115_466 ();
 sg13g2_fill_1 FILLER_115_489 ();
 sg13g2_decap_8 FILLER_115_505 ();
 sg13g2_decap_8 FILLER_115_512 ();
 sg13g2_fill_1 FILLER_115_528 ();
 sg13g2_fill_2 FILLER_115_538 ();
 sg13g2_decap_4 FILLER_115_545 ();
 sg13g2_fill_2 FILLER_115_553 ();
 sg13g2_decap_8 FILLER_115_616 ();
 sg13g2_fill_2 FILLER_115_623 ();
 sg13g2_decap_4 FILLER_115_629 ();
 sg13g2_decap_8 FILLER_115_637 ();
 sg13g2_decap_8 FILLER_115_644 ();
 sg13g2_decap_8 FILLER_115_651 ();
 sg13g2_decap_4 FILLER_115_658 ();
 sg13g2_fill_1 FILLER_115_662 ();
 sg13g2_decap_4 FILLER_115_670 ();
 sg13g2_fill_1 FILLER_115_674 ();
 sg13g2_decap_8 FILLER_115_679 ();
 sg13g2_fill_2 FILLER_115_686 ();
 sg13g2_decap_8 FILLER_115_711 ();
 sg13g2_fill_2 FILLER_115_718 ();
 sg13g2_fill_1 FILLER_115_720 ();
 sg13g2_decap_8 FILLER_115_767 ();
 sg13g2_decap_8 FILLER_115_774 ();
 sg13g2_decap_8 FILLER_115_781 ();
 sg13g2_decap_8 FILLER_115_788 ();
 sg13g2_decap_8 FILLER_115_807 ();
 sg13g2_decap_4 FILLER_115_814 ();
 sg13g2_fill_1 FILLER_115_853 ();
 sg13g2_fill_2 FILLER_115_862 ();
 sg13g2_fill_1 FILLER_115_864 ();
 sg13g2_fill_2 FILLER_115_894 ();
 sg13g2_decap_4 FILLER_115_904 ();
 sg13g2_fill_2 FILLER_115_908 ();
 sg13g2_decap_8 FILLER_115_946 ();
 sg13g2_decap_8 FILLER_115_953 ();
 sg13g2_fill_2 FILLER_115_960 ();
 sg13g2_fill_1 FILLER_115_962 ();
 sg13g2_decap_4 FILLER_115_967 ();
 sg13g2_decap_4 FILLER_115_979 ();
 sg13g2_fill_2 FILLER_115_992 ();
 sg13g2_decap_8 FILLER_115_998 ();
 sg13g2_decap_8 FILLER_115_1005 ();
 sg13g2_decap_8 FILLER_115_1012 ();
 sg13g2_decap_8 FILLER_115_1019 ();
 sg13g2_decap_8 FILLER_115_1026 ();
 sg13g2_decap_8 FILLER_115_1033 ();
 sg13g2_fill_2 FILLER_115_1040 ();
 sg13g2_fill_1 FILLER_115_1042 ();
 sg13g2_decap_8 FILLER_115_1047 ();
 sg13g2_decap_8 FILLER_115_1054 ();
 sg13g2_decap_8 FILLER_115_1065 ();
 sg13g2_decap_8 FILLER_115_1072 ();
 sg13g2_fill_2 FILLER_115_1079 ();
 sg13g2_fill_1 FILLER_115_1081 ();
 sg13g2_decap_8 FILLER_115_1090 ();
 sg13g2_decap_4 FILLER_115_1097 ();
 sg13g2_fill_1 FILLER_115_1101 ();
 sg13g2_fill_1 FILLER_115_1118 ();
 sg13g2_fill_2 FILLER_115_1123 ();
 sg13g2_fill_2 FILLER_115_1137 ();
 sg13g2_fill_2 FILLER_115_1142 ();
 sg13g2_fill_1 FILLER_115_1152 ();
 sg13g2_decap_4 FILLER_115_1158 ();
 sg13g2_fill_1 FILLER_115_1162 ();
 sg13g2_decap_8 FILLER_115_1178 ();
 sg13g2_decap_8 FILLER_115_1185 ();
 sg13g2_fill_2 FILLER_115_1192 ();
 sg13g2_fill_1 FILLER_115_1194 ();
 sg13g2_decap_8 FILLER_115_1200 ();
 sg13g2_decap_8 FILLER_115_1207 ();
 sg13g2_fill_2 FILLER_115_1240 ();
 sg13g2_fill_1 FILLER_115_1242 ();
 sg13g2_decap_8 FILLER_115_1248 ();
 sg13g2_decap_8 FILLER_115_1259 ();
 sg13g2_decap_4 FILLER_115_1266 ();
 sg13g2_decap_8 FILLER_115_1285 ();
 sg13g2_fill_2 FILLER_115_1292 ();
 sg13g2_fill_2 FILLER_115_1339 ();
 sg13g2_fill_1 FILLER_115_1341 ();
 sg13g2_fill_1 FILLER_115_1352 ();
 sg13g2_decap_8 FILLER_115_1383 ();
 sg13g2_decap_8 FILLER_115_1390 ();
 sg13g2_decap_8 FILLER_115_1397 ();
 sg13g2_decap_8 FILLER_115_1404 ();
 sg13g2_decap_8 FILLER_115_1411 ();
 sg13g2_decap_8 FILLER_115_1418 ();
 sg13g2_decap_8 FILLER_115_1425 ();
 sg13g2_decap_8 FILLER_115_1432 ();
 sg13g2_decap_8 FILLER_115_1439 ();
 sg13g2_decap_8 FILLER_115_1446 ();
 sg13g2_decap_8 FILLER_115_1453 ();
 sg13g2_decap_8 FILLER_115_1460 ();
 sg13g2_decap_8 FILLER_115_1467 ();
 sg13g2_decap_8 FILLER_115_1474 ();
 sg13g2_decap_8 FILLER_115_1481 ();
 sg13g2_decap_8 FILLER_115_1488 ();
 sg13g2_decap_8 FILLER_115_1495 ();
 sg13g2_decap_8 FILLER_115_1502 ();
 sg13g2_decap_8 FILLER_115_1509 ();
 sg13g2_decap_8 FILLER_115_1516 ();
 sg13g2_decap_8 FILLER_115_1523 ();
 sg13g2_decap_8 FILLER_115_1530 ();
 sg13g2_decap_8 FILLER_115_1537 ();
 sg13g2_decap_8 FILLER_115_1544 ();
 sg13g2_decap_8 FILLER_115_1551 ();
 sg13g2_decap_8 FILLER_115_1558 ();
 sg13g2_decap_8 FILLER_115_1565 ();
 sg13g2_decap_8 FILLER_115_1572 ();
 sg13g2_decap_8 FILLER_115_1579 ();
 sg13g2_decap_8 FILLER_115_1586 ();
 sg13g2_decap_8 FILLER_115_1593 ();
 sg13g2_decap_8 FILLER_115_1600 ();
 sg13g2_decap_8 FILLER_115_1607 ();
 sg13g2_decap_8 FILLER_115_1614 ();
 sg13g2_decap_4 FILLER_115_1621 ();
 sg13g2_decap_8 FILLER_116_0 ();
 sg13g2_decap_8 FILLER_116_7 ();
 sg13g2_decap_8 FILLER_116_14 ();
 sg13g2_decap_8 FILLER_116_21 ();
 sg13g2_decap_8 FILLER_116_28 ();
 sg13g2_decap_8 FILLER_116_35 ();
 sg13g2_decap_8 FILLER_116_42 ();
 sg13g2_decap_8 FILLER_116_49 ();
 sg13g2_decap_8 FILLER_116_56 ();
 sg13g2_decap_8 FILLER_116_63 ();
 sg13g2_decap_4 FILLER_116_103 ();
 sg13g2_decap_4 FILLER_116_117 ();
 sg13g2_fill_1 FILLER_116_121 ();
 sg13g2_fill_2 FILLER_116_144 ();
 sg13g2_fill_1 FILLER_116_146 ();
 sg13g2_decap_4 FILLER_116_152 ();
 sg13g2_fill_2 FILLER_116_181 ();
 sg13g2_fill_1 FILLER_116_183 ();
 sg13g2_fill_2 FILLER_116_215 ();
 sg13g2_fill_2 FILLER_116_222 ();
 sg13g2_fill_1 FILLER_116_229 ();
 sg13g2_fill_1 FILLER_116_247 ();
 sg13g2_decap_8 FILLER_116_274 ();
 sg13g2_decap_8 FILLER_116_281 ();
 sg13g2_decap_8 FILLER_116_288 ();
 sg13g2_fill_2 FILLER_116_295 ();
 sg13g2_fill_1 FILLER_116_297 ();
 sg13g2_fill_2 FILLER_116_311 ();
 sg13g2_decap_8 FILLER_116_339 ();
 sg13g2_decap_4 FILLER_116_355 ();
 sg13g2_fill_2 FILLER_116_359 ();
 sg13g2_decap_8 FILLER_116_365 ();
 sg13g2_decap_8 FILLER_116_389 ();
 sg13g2_decap_8 FILLER_116_396 ();
 sg13g2_decap_8 FILLER_116_403 ();
 sg13g2_decap_4 FILLER_116_410 ();
 sg13g2_decap_8 FILLER_116_419 ();
 sg13g2_fill_2 FILLER_116_426 ();
 sg13g2_fill_1 FILLER_116_428 ();
 sg13g2_decap_4 FILLER_116_439 ();
 sg13g2_fill_2 FILLER_116_446 ();
 sg13g2_fill_1 FILLER_116_448 ();
 sg13g2_decap_4 FILLER_116_470 ();
 sg13g2_fill_1 FILLER_116_474 ();
 sg13g2_fill_2 FILLER_116_479 ();
 sg13g2_fill_1 FILLER_116_489 ();
 sg13g2_decap_4 FILLER_116_501 ();
 sg13g2_fill_2 FILLER_116_505 ();
 sg13g2_decap_8 FILLER_116_511 ();
 sg13g2_decap_8 FILLER_116_518 ();
 sg13g2_fill_1 FILLER_116_525 ();
 sg13g2_decap_4 FILLER_116_531 ();
 sg13g2_fill_1 FILLER_116_535 ();
 sg13g2_decap_8 FILLER_116_566 ();
 sg13g2_decap_8 FILLER_116_573 ();
 sg13g2_decap_8 FILLER_116_580 ();
 sg13g2_decap_4 FILLER_116_587 ();
 sg13g2_fill_1 FILLER_116_591 ();
 sg13g2_decap_8 FILLER_116_600 ();
 sg13g2_decap_8 FILLER_116_607 ();
 sg13g2_decap_8 FILLER_116_618 ();
 sg13g2_fill_1 FILLER_116_625 ();
 sg13g2_decap_8 FILLER_116_652 ();
 sg13g2_decap_8 FILLER_116_659 ();
 sg13g2_decap_4 FILLER_116_666 ();
 sg13g2_fill_2 FILLER_116_670 ();
 sg13g2_fill_1 FILLER_116_680 ();
 sg13g2_decap_4 FILLER_116_686 ();
 sg13g2_fill_2 FILLER_116_690 ();
 sg13g2_decap_8 FILLER_116_699 ();
 sg13g2_fill_2 FILLER_116_706 ();
 sg13g2_decap_8 FILLER_116_714 ();
 sg13g2_decap_8 FILLER_116_721 ();
 sg13g2_decap_8 FILLER_116_728 ();
 sg13g2_decap_8 FILLER_116_735 ();
 sg13g2_fill_1 FILLER_116_742 ();
 sg13g2_fill_1 FILLER_116_748 ();
 sg13g2_decap_4 FILLER_116_753 ();
 sg13g2_decap_8 FILLER_116_766 ();
 sg13g2_decap_8 FILLER_116_773 ();
 sg13g2_fill_1 FILLER_116_780 ();
 sg13g2_fill_1 FILLER_116_786 ();
 sg13g2_fill_1 FILLER_116_793 ();
 sg13g2_fill_1 FILLER_116_804 ();
 sg13g2_fill_2 FILLER_116_809 ();
 sg13g2_decap_8 FILLER_116_824 ();
 sg13g2_decap_8 FILLER_116_831 ();
 sg13g2_decap_4 FILLER_116_838 ();
 sg13g2_fill_1 FILLER_116_842 ();
 sg13g2_decap_4 FILLER_116_847 ();
 sg13g2_fill_1 FILLER_116_851 ();
 sg13g2_decap_8 FILLER_116_888 ();
 sg13g2_decap_4 FILLER_116_895 ();
 sg13g2_decap_8 FILLER_116_907 ();
 sg13g2_fill_1 FILLER_116_914 ();
 sg13g2_decap_8 FILLER_116_929 ();
 sg13g2_decap_4 FILLER_116_936 ();
 sg13g2_fill_2 FILLER_116_940 ();
 sg13g2_fill_2 FILLER_116_959 ();
 sg13g2_fill_1 FILLER_116_961 ();
 sg13g2_decap_8 FILLER_116_972 ();
 sg13g2_fill_1 FILLER_116_979 ();
 sg13g2_fill_1 FILLER_116_1006 ();
 sg13g2_decap_4 FILLER_116_1011 ();
 sg13g2_fill_1 FILLER_116_1015 ();
 sg13g2_fill_2 FILLER_116_1026 ();
 sg13g2_fill_1 FILLER_116_1033 ();
 sg13g2_fill_1 FILLER_116_1039 ();
 sg13g2_decap_8 FILLER_116_1045 ();
 sg13g2_decap_8 FILLER_116_1086 ();
 sg13g2_fill_2 FILLER_116_1093 ();
 sg13g2_decap_8 FILLER_116_1100 ();
 sg13g2_fill_1 FILLER_116_1107 ();
 sg13g2_decap_4 FILLER_116_1116 ();
 sg13g2_decap_8 FILLER_116_1124 ();
 sg13g2_decap_8 FILLER_116_1131 ();
 sg13g2_decap_8 FILLER_116_1138 ();
 sg13g2_decap_4 FILLER_116_1145 ();
 sg13g2_fill_1 FILLER_116_1149 ();
 sg13g2_decap_4 FILLER_116_1158 ();
 sg13g2_fill_2 FILLER_116_1162 ();
 sg13g2_decap_4 FILLER_116_1180 ();
 sg13g2_fill_2 FILLER_116_1184 ();
 sg13g2_decap_8 FILLER_116_1206 ();
 sg13g2_decap_8 FILLER_116_1213 ();
 sg13g2_fill_1 FILLER_116_1220 ();
 sg13g2_fill_1 FILLER_116_1230 ();
 sg13g2_fill_2 FILLER_116_1239 ();
 sg13g2_fill_1 FILLER_116_1245 ();
 sg13g2_fill_1 FILLER_116_1272 ();
 sg13g2_decap_4 FILLER_116_1277 ();
 sg13g2_fill_2 FILLER_116_1281 ();
 sg13g2_decap_8 FILLER_116_1287 ();
 sg13g2_fill_2 FILLER_116_1294 ();
 sg13g2_fill_1 FILLER_116_1310 ();
 sg13g2_fill_1 FILLER_116_1317 ();
 sg13g2_decap_8 FILLER_116_1322 ();
 sg13g2_decap_8 FILLER_116_1329 ();
 sg13g2_decap_8 FILLER_116_1336 ();
 sg13g2_decap_8 FILLER_116_1377 ();
 sg13g2_decap_8 FILLER_116_1384 ();
 sg13g2_decap_8 FILLER_116_1391 ();
 sg13g2_decap_8 FILLER_116_1398 ();
 sg13g2_decap_8 FILLER_116_1405 ();
 sg13g2_decap_8 FILLER_116_1412 ();
 sg13g2_decap_8 FILLER_116_1419 ();
 sg13g2_decap_8 FILLER_116_1426 ();
 sg13g2_decap_8 FILLER_116_1433 ();
 sg13g2_decap_8 FILLER_116_1440 ();
 sg13g2_decap_8 FILLER_116_1447 ();
 sg13g2_decap_8 FILLER_116_1454 ();
 sg13g2_decap_8 FILLER_116_1461 ();
 sg13g2_decap_8 FILLER_116_1468 ();
 sg13g2_decap_8 FILLER_116_1475 ();
 sg13g2_decap_8 FILLER_116_1482 ();
 sg13g2_decap_8 FILLER_116_1489 ();
 sg13g2_decap_8 FILLER_116_1496 ();
 sg13g2_decap_8 FILLER_116_1503 ();
 sg13g2_decap_8 FILLER_116_1510 ();
 sg13g2_decap_8 FILLER_116_1517 ();
 sg13g2_decap_8 FILLER_116_1524 ();
 sg13g2_decap_8 FILLER_116_1531 ();
 sg13g2_decap_8 FILLER_116_1538 ();
 sg13g2_decap_8 FILLER_116_1545 ();
 sg13g2_decap_8 FILLER_116_1552 ();
 sg13g2_decap_8 FILLER_116_1559 ();
 sg13g2_decap_8 FILLER_116_1566 ();
 sg13g2_decap_8 FILLER_116_1573 ();
 sg13g2_decap_8 FILLER_116_1580 ();
 sg13g2_decap_8 FILLER_116_1587 ();
 sg13g2_decap_8 FILLER_116_1594 ();
 sg13g2_decap_8 FILLER_116_1601 ();
 sg13g2_decap_8 FILLER_116_1608 ();
 sg13g2_decap_8 FILLER_116_1615 ();
 sg13g2_fill_2 FILLER_116_1622 ();
 sg13g2_fill_1 FILLER_116_1624 ();
 sg13g2_decap_8 FILLER_117_0 ();
 sg13g2_decap_8 FILLER_117_7 ();
 sg13g2_decap_8 FILLER_117_14 ();
 sg13g2_decap_8 FILLER_117_21 ();
 sg13g2_decap_8 FILLER_117_28 ();
 sg13g2_decap_8 FILLER_117_35 ();
 sg13g2_decap_8 FILLER_117_42 ();
 sg13g2_decap_8 FILLER_117_49 ();
 sg13g2_decap_8 FILLER_117_56 ();
 sg13g2_decap_8 FILLER_117_63 ();
 sg13g2_decap_4 FILLER_117_70 ();
 sg13g2_decap_4 FILLER_117_100 ();
 sg13g2_decap_4 FILLER_117_114 ();
 sg13g2_decap_8 FILLER_117_123 ();
 sg13g2_decap_4 FILLER_117_130 ();
 sg13g2_fill_2 FILLER_117_134 ();
 sg13g2_decap_8 FILLER_117_151 ();
 sg13g2_fill_1 FILLER_117_158 ();
 sg13g2_fill_1 FILLER_117_169 ();
 sg13g2_decap_8 FILLER_117_177 ();
 sg13g2_fill_2 FILLER_117_184 ();
 sg13g2_fill_2 FILLER_117_214 ();
 sg13g2_decap_8 FILLER_117_221 ();
 sg13g2_decap_8 FILLER_117_228 ();
 sg13g2_fill_2 FILLER_117_235 ();
 sg13g2_decap_8 FILLER_117_247 ();
 sg13g2_decap_4 FILLER_117_254 ();
 sg13g2_fill_1 FILLER_117_258 ();
 sg13g2_decap_8 FILLER_117_263 ();
 sg13g2_decap_8 FILLER_117_270 ();
 sg13g2_fill_2 FILLER_117_277 ();
 sg13g2_fill_1 FILLER_117_279 ();
 sg13g2_fill_2 FILLER_117_309 ();
 sg13g2_fill_2 FILLER_117_315 ();
 sg13g2_fill_1 FILLER_117_317 ();
 sg13g2_fill_2 FILLER_117_349 ();
 sg13g2_decap_4 FILLER_117_377 ();
 sg13g2_fill_2 FILLER_117_381 ();
 sg13g2_decap_8 FILLER_117_388 ();
 sg13g2_decap_8 FILLER_117_395 ();
 sg13g2_fill_2 FILLER_117_402 ();
 sg13g2_fill_1 FILLER_117_410 ();
 sg13g2_decap_8 FILLER_117_416 ();
 sg13g2_decap_4 FILLER_117_423 ();
 sg13g2_fill_1 FILLER_117_427 ();
 sg13g2_decap_8 FILLER_117_435 ();
 sg13g2_decap_8 FILLER_117_442 ();
 sg13g2_fill_1 FILLER_117_449 ();
 sg13g2_decap_4 FILLER_117_476 ();
 sg13g2_fill_1 FILLER_117_485 ();
 sg13g2_decap_8 FILLER_117_491 ();
 sg13g2_fill_2 FILLER_117_498 ();
 sg13g2_fill_1 FILLER_117_526 ();
 sg13g2_fill_1 FILLER_117_532 ();
 sg13g2_fill_1 FILLER_117_565 ();
 sg13g2_decap_8 FILLER_117_571 ();
 sg13g2_decap_8 FILLER_117_578 ();
 sg13g2_fill_1 FILLER_117_585 ();
 sg13g2_decap_8 FILLER_117_620 ();
 sg13g2_decap_8 FILLER_117_627 ();
 sg13g2_decap_8 FILLER_117_634 ();
 sg13g2_decap_8 FILLER_117_641 ();
 sg13g2_decap_4 FILLER_117_648 ();
 sg13g2_fill_1 FILLER_117_652 ();
 sg13g2_fill_1 FILLER_117_666 ();
 sg13g2_fill_1 FILLER_117_671 ();
 sg13g2_fill_1 FILLER_117_682 ();
 sg13g2_fill_1 FILLER_117_698 ();
 sg13g2_decap_8 FILLER_117_703 ();
 sg13g2_fill_2 FILLER_117_710 ();
 sg13g2_decap_8 FILLER_117_722 ();
 sg13g2_fill_2 FILLER_117_729 ();
 sg13g2_fill_1 FILLER_117_731 ();
 sg13g2_fill_2 FILLER_117_737 ();
 sg13g2_fill_1 FILLER_117_739 ();
 sg13g2_fill_2 FILLER_117_746 ();
 sg13g2_fill_1 FILLER_117_748 ();
 sg13g2_fill_1 FILLER_117_792 ();
 sg13g2_decap_8 FILLER_117_799 ();
 sg13g2_fill_1 FILLER_117_806 ();
 sg13g2_decap_8 FILLER_117_858 ();
 sg13g2_decap_4 FILLER_117_865 ();
 sg13g2_fill_2 FILLER_117_869 ();
 sg13g2_decap_8 FILLER_117_915 ();
 sg13g2_fill_2 FILLER_117_922 ();
 sg13g2_decap_4 FILLER_117_928 ();
 sg13g2_fill_1 FILLER_117_932 ();
 sg13g2_fill_1 FILLER_117_942 ();
 sg13g2_decap_4 FILLER_117_948 ();
 sg13g2_fill_1 FILLER_117_952 ();
 sg13g2_decap_8 FILLER_117_966 ();
 sg13g2_fill_1 FILLER_117_973 ();
 sg13g2_decap_8 FILLER_117_984 ();
 sg13g2_decap_8 FILLER_117_991 ();
 sg13g2_fill_1 FILLER_117_998 ();
 sg13g2_fill_1 FILLER_117_1025 ();
 sg13g2_decap_8 FILLER_117_1095 ();
 sg13g2_decap_4 FILLER_117_1102 ();
 sg13g2_fill_2 FILLER_117_1110 ();
 sg13g2_decap_8 FILLER_117_1138 ();
 sg13g2_fill_1 FILLER_117_1145 ();
 sg13g2_decap_8 FILLER_117_1152 ();
 sg13g2_fill_2 FILLER_117_1176 ();
 sg13g2_decap_4 FILLER_117_1182 ();
 sg13g2_fill_2 FILLER_117_1186 ();
 sg13g2_decap_8 FILLER_117_1208 ();
 sg13g2_fill_2 FILLER_117_1215 ();
 sg13g2_fill_1 FILLER_117_1217 ();
 sg13g2_decap_8 FILLER_117_1223 ();
 sg13g2_decap_4 FILLER_117_1270 ();
 sg13g2_decap_4 FILLER_117_1280 ();
 sg13g2_fill_1 FILLER_117_1284 ();
 sg13g2_decap_8 FILLER_117_1290 ();
 sg13g2_decap_8 FILLER_117_1297 ();
 sg13g2_decap_8 FILLER_117_1304 ();
 sg13g2_decap_4 FILLER_117_1311 ();
 sg13g2_fill_1 FILLER_117_1315 ();
 sg13g2_decap_4 FILLER_117_1320 ();
 sg13g2_fill_2 FILLER_117_1324 ();
 sg13g2_decap_8 FILLER_117_1331 ();
 sg13g2_decap_4 FILLER_117_1343 ();
 sg13g2_fill_1 FILLER_117_1347 ();
 sg13g2_fill_1 FILLER_117_1353 ();
 sg13g2_fill_1 FILLER_117_1359 ();
 sg13g2_decap_8 FILLER_117_1389 ();
 sg13g2_decap_8 FILLER_117_1396 ();
 sg13g2_decap_8 FILLER_117_1403 ();
 sg13g2_decap_8 FILLER_117_1410 ();
 sg13g2_decap_8 FILLER_117_1417 ();
 sg13g2_decap_8 FILLER_117_1424 ();
 sg13g2_decap_8 FILLER_117_1431 ();
 sg13g2_decap_8 FILLER_117_1438 ();
 sg13g2_decap_8 FILLER_117_1445 ();
 sg13g2_decap_8 FILLER_117_1452 ();
 sg13g2_decap_8 FILLER_117_1459 ();
 sg13g2_decap_8 FILLER_117_1466 ();
 sg13g2_decap_8 FILLER_117_1473 ();
 sg13g2_decap_8 FILLER_117_1480 ();
 sg13g2_decap_8 FILLER_117_1487 ();
 sg13g2_decap_8 FILLER_117_1494 ();
 sg13g2_decap_8 FILLER_117_1501 ();
 sg13g2_decap_8 FILLER_117_1508 ();
 sg13g2_decap_8 FILLER_117_1515 ();
 sg13g2_decap_8 FILLER_117_1522 ();
 sg13g2_decap_8 FILLER_117_1529 ();
 sg13g2_decap_8 FILLER_117_1536 ();
 sg13g2_decap_8 FILLER_117_1543 ();
 sg13g2_decap_8 FILLER_117_1550 ();
 sg13g2_decap_8 FILLER_117_1557 ();
 sg13g2_decap_8 FILLER_117_1564 ();
 sg13g2_decap_8 FILLER_117_1571 ();
 sg13g2_decap_8 FILLER_117_1578 ();
 sg13g2_decap_8 FILLER_117_1585 ();
 sg13g2_decap_8 FILLER_117_1592 ();
 sg13g2_decap_8 FILLER_117_1599 ();
 sg13g2_decap_8 FILLER_117_1606 ();
 sg13g2_decap_8 FILLER_117_1613 ();
 sg13g2_decap_4 FILLER_117_1620 ();
 sg13g2_fill_1 FILLER_117_1624 ();
 sg13g2_decap_8 FILLER_118_0 ();
 sg13g2_decap_8 FILLER_118_7 ();
 sg13g2_decap_8 FILLER_118_14 ();
 sg13g2_decap_8 FILLER_118_21 ();
 sg13g2_decap_8 FILLER_118_28 ();
 sg13g2_decap_8 FILLER_118_35 ();
 sg13g2_decap_8 FILLER_118_42 ();
 sg13g2_decap_8 FILLER_118_49 ();
 sg13g2_decap_8 FILLER_118_56 ();
 sg13g2_decap_4 FILLER_118_63 ();
 sg13g2_decap_8 FILLER_118_71 ();
 sg13g2_decap_8 FILLER_118_78 ();
 sg13g2_decap_8 FILLER_118_85 ();
 sg13g2_decap_8 FILLER_118_92 ();
 sg13g2_fill_2 FILLER_118_99 ();
 sg13g2_fill_1 FILLER_118_101 ();
 sg13g2_decap_8 FILLER_118_119 ();
 sg13g2_fill_1 FILLER_118_126 ();
 sg13g2_fill_1 FILLER_118_131 ();
 sg13g2_fill_1 FILLER_118_139 ();
 sg13g2_decap_8 FILLER_118_150 ();
 sg13g2_decap_8 FILLER_118_157 ();
 sg13g2_decap_4 FILLER_118_164 ();
 sg13g2_decap_8 FILLER_118_194 ();
 sg13g2_decap_4 FILLER_118_201 ();
 sg13g2_fill_2 FILLER_118_217 ();
 sg13g2_fill_1 FILLER_118_219 ();
 sg13g2_fill_2 FILLER_118_225 ();
 sg13g2_decap_4 FILLER_118_232 ();
 sg13g2_fill_1 FILLER_118_236 ();
 sg13g2_fill_1 FILLER_118_278 ();
 sg13g2_decap_8 FILLER_118_305 ();
 sg13g2_fill_2 FILLER_118_312 ();
 sg13g2_fill_1 FILLER_118_314 ();
 sg13g2_fill_2 FILLER_118_328 ();
 sg13g2_fill_1 FILLER_118_330 ();
 sg13g2_decap_8 FILLER_118_337 ();
 sg13g2_decap_8 FILLER_118_344 ();
 sg13g2_fill_1 FILLER_118_351 ();
 sg13g2_fill_2 FILLER_118_357 ();
 sg13g2_fill_1 FILLER_118_359 ();
 sg13g2_fill_2 FILLER_118_365 ();
 sg13g2_fill_1 FILLER_118_367 ();
 sg13g2_fill_2 FILLER_118_373 ();
 sg13g2_fill_2 FILLER_118_398 ();
 sg13g2_fill_1 FILLER_118_400 ();
 sg13g2_decap_4 FILLER_118_411 ();
 sg13g2_fill_2 FILLER_118_415 ();
 sg13g2_decap_8 FILLER_118_495 ();
 sg13g2_fill_2 FILLER_118_502 ();
 sg13g2_fill_2 FILLER_118_513 ();
 sg13g2_fill_1 FILLER_118_515 ();
 sg13g2_fill_1 FILLER_118_525 ();
 sg13g2_fill_1 FILLER_118_530 ();
 sg13g2_fill_1 FILLER_118_557 ();
 sg13g2_fill_1 FILLER_118_584 ();
 sg13g2_fill_1 FILLER_118_611 ();
 sg13g2_fill_1 FILLER_118_616 ();
 sg13g2_decap_8 FILLER_118_621 ();
 sg13g2_decap_4 FILLER_118_628 ();
 sg13g2_decap_4 FILLER_118_636 ();
 sg13g2_fill_2 FILLER_118_640 ();
 sg13g2_decap_8 FILLER_118_652 ();
 sg13g2_decap_8 FILLER_118_659 ();
 sg13g2_fill_1 FILLER_118_666 ();
 sg13g2_fill_2 FILLER_118_671 ();
 sg13g2_decap_4 FILLER_118_677 ();
 sg13g2_decap_8 FILLER_118_690 ();
 sg13g2_fill_1 FILLER_118_697 ();
 sg13g2_fill_1 FILLER_118_724 ();
 sg13g2_fill_1 FILLER_118_730 ();
 sg13g2_fill_1 FILLER_118_745 ();
 sg13g2_decap_8 FILLER_118_752 ();
 sg13g2_decap_4 FILLER_118_759 ();
 sg13g2_fill_2 FILLER_118_763 ();
 sg13g2_decap_8 FILLER_118_769 ();
 sg13g2_decap_8 FILLER_118_776 ();
 sg13g2_fill_2 FILLER_118_783 ();
 sg13g2_fill_1 FILLER_118_785 ();
 sg13g2_decap_8 FILLER_118_799 ();
 sg13g2_decap_4 FILLER_118_806 ();
 sg13g2_decap_8 FILLER_118_823 ();
 sg13g2_decap_8 FILLER_118_830 ();
 sg13g2_fill_1 FILLER_118_847 ();
 sg13g2_decap_8 FILLER_118_862 ();
 sg13g2_fill_2 FILLER_118_869 ();
 sg13g2_decap_8 FILLER_118_876 ();
 sg13g2_decap_4 FILLER_118_883 ();
 sg13g2_decap_8 FILLER_118_900 ();
 sg13g2_fill_1 FILLER_118_916 ();
 sg13g2_fill_1 FILLER_118_922 ();
 sg13g2_decap_8 FILLER_118_929 ();
 sg13g2_decap_4 FILLER_118_936 ();
 sg13g2_decap_8 FILLER_118_967 ();
 sg13g2_decap_8 FILLER_118_984 ();
 sg13g2_fill_2 FILLER_118_991 ();
 sg13g2_fill_1 FILLER_118_993 ();
 sg13g2_fill_1 FILLER_118_1023 ();
 sg13g2_fill_2 FILLER_118_1039 ();
 sg13g2_fill_1 FILLER_118_1041 ();
 sg13g2_decap_8 FILLER_118_1051 ();
 sg13g2_fill_2 FILLER_118_1093 ();
 sg13g2_fill_1 FILLER_118_1095 ();
 sg13g2_decap_8 FILLER_118_1110 ();
 sg13g2_fill_2 FILLER_118_1117 ();
 sg13g2_fill_1 FILLER_118_1119 ();
 sg13g2_decap_4 FILLER_118_1125 ();
 sg13g2_fill_1 FILLER_118_1129 ();
 sg13g2_fill_1 FILLER_118_1166 ();
 sg13g2_fill_2 FILLER_118_1182 ();
 sg13g2_decap_8 FILLER_118_1201 ();
 sg13g2_decap_8 FILLER_118_1208 ();
 sg13g2_decap_8 FILLER_118_1215 ();
 sg13g2_fill_2 FILLER_118_1222 ();
 sg13g2_fill_1 FILLER_118_1224 ();
 sg13g2_decap_8 FILLER_118_1230 ();
 sg13g2_decap_8 FILLER_118_1237 ();
 sg13g2_decap_4 FILLER_118_1244 ();
 sg13g2_decap_8 FILLER_118_1259 ();
 sg13g2_decap_8 FILLER_118_1266 ();
 sg13g2_fill_2 FILLER_118_1273 ();
 sg13g2_fill_1 FILLER_118_1275 ();
 sg13g2_decap_8 FILLER_118_1281 ();
 sg13g2_decap_8 FILLER_118_1294 ();
 sg13g2_decap_4 FILLER_118_1301 ();
 sg13g2_fill_2 FILLER_118_1305 ();
 sg13g2_fill_1 FILLER_118_1321 ();
 sg13g2_decap_8 FILLER_118_1331 ();
 sg13g2_decap_8 FILLER_118_1338 ();
 sg13g2_decap_4 FILLER_118_1345 ();
 sg13g2_fill_2 FILLER_118_1349 ();
 sg13g2_fill_1 FILLER_118_1360 ();
 sg13g2_decap_8 FILLER_118_1387 ();
 sg13g2_decap_8 FILLER_118_1394 ();
 sg13g2_decap_8 FILLER_118_1401 ();
 sg13g2_decap_8 FILLER_118_1408 ();
 sg13g2_decap_8 FILLER_118_1415 ();
 sg13g2_decap_8 FILLER_118_1422 ();
 sg13g2_decap_8 FILLER_118_1429 ();
 sg13g2_decap_8 FILLER_118_1436 ();
 sg13g2_decap_8 FILLER_118_1443 ();
 sg13g2_decap_8 FILLER_118_1450 ();
 sg13g2_decap_8 FILLER_118_1457 ();
 sg13g2_decap_8 FILLER_118_1464 ();
 sg13g2_decap_8 FILLER_118_1471 ();
 sg13g2_decap_8 FILLER_118_1478 ();
 sg13g2_decap_8 FILLER_118_1485 ();
 sg13g2_decap_8 FILLER_118_1492 ();
 sg13g2_decap_8 FILLER_118_1499 ();
 sg13g2_decap_8 FILLER_118_1506 ();
 sg13g2_decap_8 FILLER_118_1513 ();
 sg13g2_decap_8 FILLER_118_1520 ();
 sg13g2_decap_8 FILLER_118_1527 ();
 sg13g2_decap_8 FILLER_118_1534 ();
 sg13g2_decap_8 FILLER_118_1541 ();
 sg13g2_decap_8 FILLER_118_1548 ();
 sg13g2_decap_8 FILLER_118_1555 ();
 sg13g2_decap_8 FILLER_118_1562 ();
 sg13g2_decap_8 FILLER_118_1569 ();
 sg13g2_decap_8 FILLER_118_1576 ();
 sg13g2_decap_8 FILLER_118_1583 ();
 sg13g2_decap_8 FILLER_118_1590 ();
 sg13g2_decap_8 FILLER_118_1597 ();
 sg13g2_decap_8 FILLER_118_1604 ();
 sg13g2_decap_8 FILLER_118_1611 ();
 sg13g2_decap_8 FILLER_118_1618 ();
 sg13g2_decap_8 FILLER_119_0 ();
 sg13g2_decap_8 FILLER_119_7 ();
 sg13g2_decap_8 FILLER_119_14 ();
 sg13g2_decap_8 FILLER_119_21 ();
 sg13g2_decap_8 FILLER_119_28 ();
 sg13g2_decap_8 FILLER_119_35 ();
 sg13g2_decap_8 FILLER_119_42 ();
 sg13g2_decap_8 FILLER_119_49 ();
 sg13g2_decap_4 FILLER_119_56 ();
 sg13g2_fill_1 FILLER_119_60 ();
 sg13g2_decap_4 FILLER_119_87 ();
 sg13g2_decap_4 FILLER_119_118 ();
 sg13g2_decap_8 FILLER_119_153 ();
 sg13g2_decap_8 FILLER_119_160 ();
 sg13g2_decap_4 FILLER_119_167 ();
 sg13g2_decap_8 FILLER_119_180 ();
 sg13g2_decap_4 FILLER_119_187 ();
 sg13g2_fill_2 FILLER_119_191 ();
 sg13g2_decap_8 FILLER_119_197 ();
 sg13g2_fill_1 FILLER_119_204 ();
 sg13g2_decap_8 FILLER_119_225 ();
 sg13g2_decap_8 FILLER_119_232 ();
 sg13g2_fill_2 FILLER_119_251 ();
 sg13g2_fill_1 FILLER_119_253 ();
 sg13g2_decap_8 FILLER_119_279 ();
 sg13g2_decap_8 FILLER_119_286 ();
 sg13g2_decap_4 FILLER_119_293 ();
 sg13g2_fill_1 FILLER_119_297 ();
 sg13g2_fill_2 FILLER_119_313 ();
 sg13g2_decap_8 FILLER_119_337 ();
 sg13g2_decap_8 FILLER_119_344 ();
 sg13g2_decap_8 FILLER_119_351 ();
 sg13g2_decap_4 FILLER_119_358 ();
 sg13g2_fill_2 FILLER_119_362 ();
 sg13g2_fill_1 FILLER_119_372 ();
 sg13g2_decap_8 FILLER_119_388 ();
 sg13g2_decap_8 FILLER_119_395 ();
 sg13g2_decap_8 FILLER_119_402 ();
 sg13g2_decap_8 FILLER_119_409 ();
 sg13g2_fill_2 FILLER_119_416 ();
 sg13g2_fill_1 FILLER_119_418 ();
 sg13g2_fill_2 FILLER_119_424 ();
 sg13g2_decap_8 FILLER_119_431 ();
 sg13g2_decap_8 FILLER_119_438 ();
 sg13g2_fill_2 FILLER_119_445 ();
 sg13g2_decap_4 FILLER_119_453 ();
 sg13g2_decap_8 FILLER_119_471 ();
 sg13g2_decap_8 FILLER_119_478 ();
 sg13g2_decap_8 FILLER_119_485 ();
 sg13g2_fill_2 FILLER_119_492 ();
 sg13g2_fill_1 FILLER_119_494 ();
 sg13g2_fill_2 FILLER_119_500 ();
 sg13g2_fill_1 FILLER_119_502 ();
 sg13g2_decap_8 FILLER_119_528 ();
 sg13g2_decap_8 FILLER_119_535 ();
 sg13g2_decap_8 FILLER_119_542 ();
 sg13g2_decap_8 FILLER_119_549 ();
 sg13g2_decap_8 FILLER_119_556 ();
 sg13g2_fill_1 FILLER_119_563 ();
 sg13g2_decap_8 FILLER_119_572 ();
 sg13g2_decap_8 FILLER_119_579 ();
 sg13g2_decap_8 FILLER_119_586 ();
 sg13g2_decap_4 FILLER_119_593 ();
 sg13g2_fill_2 FILLER_119_597 ();
 sg13g2_fill_1 FILLER_119_611 ();
 sg13g2_decap_8 FILLER_119_634 ();
 sg13g2_fill_1 FILLER_119_641 ();
 sg13g2_fill_1 FILLER_119_672 ();
 sg13g2_fill_2 FILLER_119_681 ();
 sg13g2_fill_1 FILLER_119_687 ();
 sg13g2_fill_2 FILLER_119_693 ();
 sg13g2_fill_2 FILLER_119_699 ();
 sg13g2_decap_8 FILLER_119_705 ();
 sg13g2_decap_4 FILLER_119_712 ();
 sg13g2_fill_1 FILLER_119_726 ();
 sg13g2_fill_1 FILLER_119_731 ();
 sg13g2_fill_1 FILLER_119_737 ();
 sg13g2_fill_1 FILLER_119_743 ();
 sg13g2_decap_4 FILLER_119_751 ();
 sg13g2_decap_8 FILLER_119_761 ();
 sg13g2_decap_4 FILLER_119_773 ();
 sg13g2_fill_1 FILLER_119_777 ();
 sg13g2_fill_1 FILLER_119_784 ();
 sg13g2_decap_8 FILLER_119_791 ();
 sg13g2_decap_8 FILLER_119_798 ();
 sg13g2_fill_1 FILLER_119_805 ();
 sg13g2_fill_2 FILLER_119_813 ();
 sg13g2_decap_8 FILLER_119_825 ();
 sg13g2_decap_8 FILLER_119_832 ();
 sg13g2_decap_8 FILLER_119_839 ();
 sg13g2_decap_8 FILLER_119_855 ();
 sg13g2_decap_8 FILLER_119_870 ();
 sg13g2_decap_4 FILLER_119_881 ();
 sg13g2_fill_1 FILLER_119_885 ();
 sg13g2_fill_2 FILLER_119_894 ();
 sg13g2_fill_1 FILLER_119_896 ();
 sg13g2_decap_8 FILLER_119_902 ();
 sg13g2_decap_8 FILLER_119_909 ();
 sg13g2_decap_8 FILLER_119_916 ();
 sg13g2_fill_1 FILLER_119_928 ();
 sg13g2_decap_8 FILLER_119_935 ();
 sg13g2_fill_2 FILLER_119_942 ();
 sg13g2_decap_8 FILLER_119_958 ();
 sg13g2_decap_4 FILLER_119_965 ();
 sg13g2_fill_2 FILLER_119_969 ();
 sg13g2_fill_1 FILLER_119_981 ();
 sg13g2_fill_2 FILLER_119_990 ();
 sg13g2_fill_2 FILLER_119_1023 ();
 sg13g2_decap_8 FILLER_119_1055 ();
 sg13g2_fill_2 FILLER_119_1062 ();
 sg13g2_fill_1 FILLER_119_1064 ();
 sg13g2_decap_4 FILLER_119_1070 ();
 sg13g2_fill_1 FILLER_119_1074 ();
 sg13g2_fill_2 FILLER_119_1079 ();
 sg13g2_decap_4 FILLER_119_1095 ();
 sg13g2_fill_1 FILLER_119_1099 ();
 sg13g2_fill_2 FILLER_119_1126 ();
 sg13g2_fill_1 FILLER_119_1128 ();
 sg13g2_fill_2 FILLER_119_1133 ();
 sg13g2_fill_2 FILLER_119_1143 ();
 sg13g2_fill_1 FILLER_119_1145 ();
 sg13g2_decap_8 FILLER_119_1171 ();
 sg13g2_fill_1 FILLER_119_1196 ();
 sg13g2_fill_2 FILLER_119_1205 ();
 sg13g2_decap_8 FILLER_119_1215 ();
 sg13g2_fill_2 FILLER_119_1226 ();
 sg13g2_fill_1 FILLER_119_1228 ();
 sg13g2_fill_2 FILLER_119_1247 ();
 sg13g2_decap_8 FILLER_119_1255 ();
 sg13g2_decap_8 FILLER_119_1262 ();
 sg13g2_decap_4 FILLER_119_1269 ();
 sg13g2_fill_1 FILLER_119_1273 ();
 sg13g2_fill_1 FILLER_119_1278 ();
 sg13g2_fill_1 FILLER_119_1284 ();
 sg13g2_decap_8 FILLER_119_1291 ();
 sg13g2_decap_8 FILLER_119_1298 ();
 sg13g2_decap_8 FILLER_119_1318 ();
 sg13g2_fill_1 FILLER_119_1325 ();
 sg13g2_decap_4 FILLER_119_1341 ();
 sg13g2_decap_8 FILLER_119_1385 ();
 sg13g2_decap_8 FILLER_119_1392 ();
 sg13g2_decap_8 FILLER_119_1399 ();
 sg13g2_decap_8 FILLER_119_1406 ();
 sg13g2_decap_8 FILLER_119_1413 ();
 sg13g2_decap_8 FILLER_119_1420 ();
 sg13g2_decap_8 FILLER_119_1427 ();
 sg13g2_decap_8 FILLER_119_1434 ();
 sg13g2_decap_8 FILLER_119_1441 ();
 sg13g2_decap_8 FILLER_119_1448 ();
 sg13g2_decap_8 FILLER_119_1455 ();
 sg13g2_decap_8 FILLER_119_1462 ();
 sg13g2_decap_8 FILLER_119_1469 ();
 sg13g2_decap_8 FILLER_119_1476 ();
 sg13g2_decap_8 FILLER_119_1483 ();
 sg13g2_decap_8 FILLER_119_1490 ();
 sg13g2_decap_8 FILLER_119_1497 ();
 sg13g2_decap_8 FILLER_119_1504 ();
 sg13g2_decap_8 FILLER_119_1511 ();
 sg13g2_decap_8 FILLER_119_1518 ();
 sg13g2_decap_8 FILLER_119_1525 ();
 sg13g2_decap_8 FILLER_119_1532 ();
 sg13g2_decap_8 FILLER_119_1539 ();
 sg13g2_decap_8 FILLER_119_1546 ();
 sg13g2_decap_8 FILLER_119_1553 ();
 sg13g2_decap_8 FILLER_119_1560 ();
 sg13g2_decap_8 FILLER_119_1567 ();
 sg13g2_decap_8 FILLER_119_1574 ();
 sg13g2_decap_8 FILLER_119_1581 ();
 sg13g2_decap_8 FILLER_119_1588 ();
 sg13g2_decap_8 FILLER_119_1595 ();
 sg13g2_decap_8 FILLER_119_1602 ();
 sg13g2_decap_8 FILLER_119_1609 ();
 sg13g2_decap_8 FILLER_119_1616 ();
 sg13g2_fill_2 FILLER_119_1623 ();
 sg13g2_decap_8 FILLER_120_0 ();
 sg13g2_decap_8 FILLER_120_7 ();
 sg13g2_decap_8 FILLER_120_14 ();
 sg13g2_decap_8 FILLER_120_21 ();
 sg13g2_decap_8 FILLER_120_28 ();
 sg13g2_decap_8 FILLER_120_35 ();
 sg13g2_decap_8 FILLER_120_42 ();
 sg13g2_decap_8 FILLER_120_49 ();
 sg13g2_decap_4 FILLER_120_56 ();
 sg13g2_decap_8 FILLER_120_64 ();
 sg13g2_decap_8 FILLER_120_71 ();
 sg13g2_decap_8 FILLER_120_78 ();
 sg13g2_decap_8 FILLER_120_85 ();
 sg13g2_decap_4 FILLER_120_92 ();
 sg13g2_fill_2 FILLER_120_96 ();
 sg13g2_decap_8 FILLER_120_108 ();
 sg13g2_decap_8 FILLER_120_115 ();
 sg13g2_decap_8 FILLER_120_122 ();
 sg13g2_decap_8 FILLER_120_129 ();
 sg13g2_decap_8 FILLER_120_136 ();
 sg13g2_decap_8 FILLER_120_143 ();
 sg13g2_decap_8 FILLER_120_150 ();
 sg13g2_decap_8 FILLER_120_157 ();
 sg13g2_decap_8 FILLER_120_164 ();
 sg13g2_fill_2 FILLER_120_171 ();
 sg13g2_fill_1 FILLER_120_173 ();
 sg13g2_decap_8 FILLER_120_179 ();
 sg13g2_decap_8 FILLER_120_224 ();
 sg13g2_decap_8 FILLER_120_231 ();
 sg13g2_decap_4 FILLER_120_238 ();
 sg13g2_decap_8 FILLER_120_247 ();
 sg13g2_fill_2 FILLER_120_254 ();
 sg13g2_decap_8 FILLER_120_260 ();
 sg13g2_decap_8 FILLER_120_267 ();
 sg13g2_decap_8 FILLER_120_274 ();
 sg13g2_fill_1 FILLER_120_281 ();
 sg13g2_decap_8 FILLER_120_286 ();
 sg13g2_decap_8 FILLER_120_293 ();
 sg13g2_decap_8 FILLER_120_300 ();
 sg13g2_decap_8 FILLER_120_307 ();
 sg13g2_decap_8 FILLER_120_314 ();
 sg13g2_decap_8 FILLER_120_321 ();
 sg13g2_decap_8 FILLER_120_328 ();
 sg13g2_fill_2 FILLER_120_335 ();
 sg13g2_fill_1 FILLER_120_337 ();
 sg13g2_fill_2 FILLER_120_342 ();
 sg13g2_decap_8 FILLER_120_389 ();
 sg13g2_decap_8 FILLER_120_396 ();
 sg13g2_fill_2 FILLER_120_415 ();
 sg13g2_decap_8 FILLER_120_425 ();
 sg13g2_decap_4 FILLER_120_432 ();
 sg13g2_fill_2 FILLER_120_454 ();
 sg13g2_decap_8 FILLER_120_468 ();
 sg13g2_fill_2 FILLER_120_484 ();
 sg13g2_fill_1 FILLER_120_486 ();
 sg13g2_fill_1 FILLER_120_496 ();
 sg13g2_decap_8 FILLER_120_523 ();
 sg13g2_decap_8 FILLER_120_535 ();
 sg13g2_fill_2 FILLER_120_542 ();
 sg13g2_fill_2 FILLER_120_553 ();
 sg13g2_fill_1 FILLER_120_555 ();
 sg13g2_decap_4 FILLER_120_561 ();
 sg13g2_fill_1 FILLER_120_565 ();
 sg13g2_decap_8 FILLER_120_571 ();
 sg13g2_decap_8 FILLER_120_578 ();
 sg13g2_fill_1 FILLER_120_585 ();
 sg13g2_fill_2 FILLER_120_606 ();
 sg13g2_decap_8 FILLER_120_622 ();
 sg13g2_fill_2 FILLER_120_629 ();
 sg13g2_fill_1 FILLER_120_644 ();
 sg13g2_decap_8 FILLER_120_649 ();
 sg13g2_decap_8 FILLER_120_656 ();
 sg13g2_decap_8 FILLER_120_663 ();
 sg13g2_decap_8 FILLER_120_675 ();
 sg13g2_decap_8 FILLER_120_682 ();
 sg13g2_decap_8 FILLER_120_689 ();
 sg13g2_decap_4 FILLER_120_696 ();
 sg13g2_fill_2 FILLER_120_700 ();
 sg13g2_fill_2 FILLER_120_707 ();
 sg13g2_fill_1 FILLER_120_709 ();
 sg13g2_fill_2 FILLER_120_732 ();
 sg13g2_decap_8 FILLER_120_744 ();
 sg13g2_decap_8 FILLER_120_751 ();
 sg13g2_fill_2 FILLER_120_758 ();
 sg13g2_fill_1 FILLER_120_760 ();
 sg13g2_decap_8 FILLER_120_769 ();
 sg13g2_fill_2 FILLER_120_776 ();
 sg13g2_decap_4 FILLER_120_788 ();
 sg13g2_fill_2 FILLER_120_800 ();
 sg13g2_fill_2 FILLER_120_815 ();
 sg13g2_fill_1 FILLER_120_817 ();
 sg13g2_decap_4 FILLER_120_825 ();
 sg13g2_decap_8 FILLER_120_835 ();
 sg13g2_decap_8 FILLER_120_847 ();
 sg13g2_decap_8 FILLER_120_854 ();
 sg13g2_fill_2 FILLER_120_861 ();
 sg13g2_fill_2 FILLER_120_896 ();
 sg13g2_fill_1 FILLER_120_898 ();
 sg13g2_decap_8 FILLER_120_904 ();
 sg13g2_decap_8 FILLER_120_911 ();
 sg13g2_decap_8 FILLER_120_918 ();
 sg13g2_decap_8 FILLER_120_925 ();
 sg13g2_decap_8 FILLER_120_932 ();
 sg13g2_decap_8 FILLER_120_939 ();
 sg13g2_decap_8 FILLER_120_946 ();
 sg13g2_fill_2 FILLER_120_953 ();
 sg13g2_decap_8 FILLER_120_973 ();
 sg13g2_decap_8 FILLER_120_980 ();
 sg13g2_decap_8 FILLER_120_987 ();
 sg13g2_fill_1 FILLER_120_994 ();
 sg13g2_decap_8 FILLER_120_1002 ();
 sg13g2_decap_8 FILLER_120_1009 ();
 sg13g2_decap_8 FILLER_120_1016 ();
 sg13g2_decap_8 FILLER_120_1023 ();
 sg13g2_decap_4 FILLER_120_1033 ();
 sg13g2_fill_1 FILLER_120_1037 ();
 sg13g2_decap_8 FILLER_120_1064 ();
 sg13g2_fill_2 FILLER_120_1071 ();
 sg13g2_fill_1 FILLER_120_1073 ();
 sg13g2_decap_8 FILLER_120_1084 ();
 sg13g2_decap_8 FILLER_120_1091 ();
 sg13g2_decap_8 FILLER_120_1098 ();
 sg13g2_fill_2 FILLER_120_1105 ();
 sg13g2_fill_2 FILLER_120_1141 ();
 sg13g2_fill_1 FILLER_120_1143 ();
 sg13g2_decap_8 FILLER_120_1213 ();
 sg13g2_decap_8 FILLER_120_1220 ();
 sg13g2_fill_2 FILLER_120_1227 ();
 sg13g2_decap_8 FILLER_120_1255 ();
 sg13g2_fill_2 FILLER_120_1262 ();
 sg13g2_fill_1 FILLER_120_1264 ();
 sg13g2_decap_4 FILLER_120_1299 ();
 sg13g2_fill_2 FILLER_120_1303 ();
 sg13g2_decap_8 FILLER_120_1316 ();
 sg13g2_decap_8 FILLER_120_1333 ();
 sg13g2_fill_2 FILLER_120_1340 ();
 sg13g2_decap_8 FILLER_120_1347 ();
 sg13g2_decap_8 FILLER_120_1354 ();
 sg13g2_fill_2 FILLER_120_1361 ();
 sg13g2_decap_8 FILLER_120_1367 ();
 sg13g2_decap_8 FILLER_120_1374 ();
 sg13g2_decap_8 FILLER_120_1381 ();
 sg13g2_decap_8 FILLER_120_1388 ();
 sg13g2_decap_8 FILLER_120_1395 ();
 sg13g2_decap_8 FILLER_120_1402 ();
 sg13g2_decap_8 FILLER_120_1409 ();
 sg13g2_decap_8 FILLER_120_1416 ();
 sg13g2_decap_8 FILLER_120_1423 ();
 sg13g2_decap_8 FILLER_120_1430 ();
 sg13g2_decap_8 FILLER_120_1437 ();
 sg13g2_decap_8 FILLER_120_1444 ();
 sg13g2_decap_8 FILLER_120_1451 ();
 sg13g2_decap_8 FILLER_120_1458 ();
 sg13g2_decap_8 FILLER_120_1465 ();
 sg13g2_decap_8 FILLER_120_1472 ();
 sg13g2_decap_8 FILLER_120_1479 ();
 sg13g2_decap_8 FILLER_120_1486 ();
 sg13g2_decap_8 FILLER_120_1493 ();
 sg13g2_decap_8 FILLER_120_1500 ();
 sg13g2_decap_8 FILLER_120_1507 ();
 sg13g2_decap_8 FILLER_120_1514 ();
 sg13g2_decap_8 FILLER_120_1521 ();
 sg13g2_decap_8 FILLER_120_1528 ();
 sg13g2_decap_8 FILLER_120_1535 ();
 sg13g2_decap_8 FILLER_120_1542 ();
 sg13g2_decap_8 FILLER_120_1549 ();
 sg13g2_decap_8 FILLER_120_1556 ();
 sg13g2_decap_8 FILLER_120_1563 ();
 sg13g2_decap_8 FILLER_120_1570 ();
 sg13g2_decap_8 FILLER_120_1577 ();
 sg13g2_decap_8 FILLER_120_1584 ();
 sg13g2_decap_8 FILLER_120_1591 ();
 sg13g2_decap_8 FILLER_120_1598 ();
 sg13g2_decap_8 FILLER_120_1605 ();
 sg13g2_decap_8 FILLER_120_1612 ();
 sg13g2_decap_4 FILLER_120_1619 ();
 sg13g2_fill_2 FILLER_120_1623 ();
 sg13g2_decap_8 FILLER_121_0 ();
 sg13g2_decap_8 FILLER_121_7 ();
 sg13g2_decap_8 FILLER_121_14 ();
 sg13g2_decap_8 FILLER_121_21 ();
 sg13g2_decap_8 FILLER_121_28 ();
 sg13g2_decap_8 FILLER_121_35 ();
 sg13g2_decap_8 FILLER_121_42 ();
 sg13g2_decap_4 FILLER_121_49 ();
 sg13g2_fill_1 FILLER_121_53 ();
 sg13g2_fill_2 FILLER_121_92 ();
 sg13g2_fill_1 FILLER_121_94 ();
 sg13g2_decap_8 FILLER_121_100 ();
 sg13g2_decap_8 FILLER_121_107 ();
 sg13g2_decap_8 FILLER_121_114 ();
 sg13g2_decap_8 FILLER_121_121 ();
 sg13g2_decap_8 FILLER_121_128 ();
 sg13g2_fill_2 FILLER_121_135 ();
 sg13g2_decap_8 FILLER_121_141 ();
 sg13g2_decap_8 FILLER_121_148 ();
 sg13g2_decap_4 FILLER_121_155 ();
 sg13g2_fill_2 FILLER_121_159 ();
 sg13g2_decap_4 FILLER_121_183 ();
 sg13g2_fill_2 FILLER_121_187 ();
 sg13g2_decap_8 FILLER_121_193 ();
 sg13g2_decap_8 FILLER_121_200 ();
 sg13g2_decap_4 FILLER_121_207 ();
 sg13g2_fill_2 FILLER_121_211 ();
 sg13g2_fill_2 FILLER_121_218 ();
 sg13g2_fill_1 FILLER_121_220 ();
 sg13g2_fill_2 FILLER_121_226 ();
 sg13g2_fill_1 FILLER_121_274 ();
 sg13g2_decap_4 FILLER_121_301 ();
 sg13g2_fill_1 FILLER_121_305 ();
 sg13g2_fill_2 FILLER_121_321 ();
 sg13g2_fill_1 FILLER_121_323 ();
 sg13g2_decap_4 FILLER_121_332 ();
 sg13g2_fill_2 FILLER_121_336 ();
 sg13g2_decap_8 FILLER_121_342 ();
 sg13g2_decap_8 FILLER_121_349 ();
 sg13g2_decap_8 FILLER_121_356 ();
 sg13g2_decap_4 FILLER_121_363 ();
 sg13g2_fill_1 FILLER_121_379 ();
 sg13g2_fill_2 FILLER_121_385 ();
 sg13g2_decap_8 FILLER_121_399 ();
 sg13g2_decap_4 FILLER_121_423 ();
 sg13g2_fill_1 FILLER_121_427 ();
 sg13g2_decap_4 FILLER_121_443 ();
 sg13g2_decap_8 FILLER_121_453 ();
 sg13g2_decap_8 FILLER_121_460 ();
 sg13g2_fill_1 FILLER_121_467 ();
 sg13g2_decap_8 FILLER_121_533 ();
 sg13g2_decap_4 FILLER_121_566 ();
 sg13g2_fill_2 FILLER_121_570 ();
 sg13g2_decap_4 FILLER_121_581 ();
 sg13g2_decap_4 FILLER_121_590 ();
 sg13g2_fill_2 FILLER_121_602 ();
 sg13g2_fill_1 FILLER_121_604 ();
 sg13g2_decap_8 FILLER_121_613 ();
 sg13g2_decap_8 FILLER_121_620 ();
 sg13g2_fill_2 FILLER_121_627 ();
 sg13g2_decap_8 FILLER_121_633 ();
 sg13g2_decap_4 FILLER_121_640 ();
 sg13g2_fill_2 FILLER_121_644 ();
 sg13g2_decap_8 FILLER_121_655 ();
 sg13g2_fill_2 FILLER_121_662 ();
 sg13g2_decap_4 FILLER_121_669 ();
 sg13g2_fill_1 FILLER_121_673 ();
 sg13g2_fill_1 FILLER_121_679 ();
 sg13g2_decap_8 FILLER_121_684 ();
 sg13g2_decap_8 FILLER_121_691 ();
 sg13g2_fill_1 FILLER_121_698 ();
 sg13g2_decap_8 FILLER_121_716 ();
 sg13g2_decap_8 FILLER_121_723 ();
 sg13g2_decap_8 FILLER_121_730 ();
 sg13g2_decap_8 FILLER_121_737 ();
 sg13g2_decap_8 FILLER_121_744 ();
 sg13g2_fill_2 FILLER_121_751 ();
 sg13g2_fill_1 FILLER_121_753 ();
 sg13g2_decap_8 FILLER_121_771 ();
 sg13g2_fill_2 FILLER_121_778 ();
 sg13g2_fill_1 FILLER_121_780 ();
 sg13g2_decap_8 FILLER_121_796 ();
 sg13g2_decap_8 FILLER_121_803 ();
 sg13g2_decap_4 FILLER_121_810 ();
 sg13g2_fill_1 FILLER_121_814 ();
 sg13g2_fill_1 FILLER_121_832 ();
 sg13g2_fill_2 FILLER_121_845 ();
 sg13g2_fill_1 FILLER_121_847 ();
 sg13g2_fill_2 FILLER_121_853 ();
 sg13g2_fill_1 FILLER_121_870 ();
 sg13g2_decap_8 FILLER_121_880 ();
 sg13g2_fill_1 FILLER_121_887 ();
 sg13g2_decap_8 FILLER_121_892 ();
 sg13g2_decap_8 FILLER_121_899 ();
 sg13g2_decap_4 FILLER_121_906 ();
 sg13g2_fill_1 FILLER_121_910 ();
 sg13g2_decap_8 FILLER_121_921 ();
 sg13g2_decap_4 FILLER_121_928 ();
 sg13g2_fill_2 FILLER_121_962 ();
 sg13g2_decap_8 FILLER_121_968 ();
 sg13g2_decap_4 FILLER_121_975 ();
 sg13g2_fill_2 FILLER_121_979 ();
 sg13g2_fill_2 FILLER_121_985 ();
 sg13g2_fill_2 FILLER_121_1014 ();
 sg13g2_fill_1 FILLER_121_1016 ();
 sg13g2_decap_8 FILLER_121_1030 ();
 sg13g2_decap_8 FILLER_121_1037 ();
 sg13g2_fill_2 FILLER_121_1044 ();
 sg13g2_decap_8 FILLER_121_1050 ();
 sg13g2_decap_8 FILLER_121_1057 ();
 sg13g2_decap_8 FILLER_121_1064 ();
 sg13g2_decap_8 FILLER_121_1071 ();
 sg13g2_fill_2 FILLER_121_1078 ();
 sg13g2_fill_1 FILLER_121_1080 ();
 sg13g2_fill_2 FILLER_121_1090 ();
 sg13g2_fill_1 FILLER_121_1092 ();
 sg13g2_decap_8 FILLER_121_1097 ();
 sg13g2_decap_8 FILLER_121_1104 ();
 sg13g2_decap_8 FILLER_121_1111 ();
 sg13g2_fill_2 FILLER_121_1118 ();
 sg13g2_fill_1 FILLER_121_1120 ();
 sg13g2_decap_4 FILLER_121_1153 ();
 sg13g2_decap_8 FILLER_121_1161 ();
 sg13g2_decap_8 FILLER_121_1168 ();
 sg13g2_decap_4 FILLER_121_1175 ();
 sg13g2_decap_8 FILLER_121_1184 ();
 sg13g2_decap_4 FILLER_121_1191 ();
 sg13g2_fill_1 FILLER_121_1195 ();
 sg13g2_decap_8 FILLER_121_1204 ();
 sg13g2_decap_8 FILLER_121_1211 ();
 sg13g2_decap_4 FILLER_121_1218 ();
 sg13g2_decap_8 FILLER_121_1233 ();
 sg13g2_decap_8 FILLER_121_1240 ();
 sg13g2_fill_1 FILLER_121_1247 ();
 sg13g2_decap_4 FILLER_121_1259 ();
 sg13g2_fill_1 FILLER_121_1263 ();
 sg13g2_fill_1 FILLER_121_1278 ();
 sg13g2_decap_8 FILLER_121_1284 ();
 sg13g2_decap_8 FILLER_121_1291 ();
 sg13g2_decap_4 FILLER_121_1298 ();
 sg13g2_decap_4 FILLER_121_1313 ();
 sg13g2_fill_2 FILLER_121_1317 ();
 sg13g2_fill_1 FILLER_121_1323 ();
 sg13g2_fill_1 FILLER_121_1329 ();
 sg13g2_fill_1 FILLER_121_1336 ();
 sg13g2_fill_1 FILLER_121_1342 ();
 sg13g2_fill_2 FILLER_121_1351 ();
 sg13g2_decap_8 FILLER_121_1357 ();
 sg13g2_decap_8 FILLER_121_1364 ();
 sg13g2_decap_8 FILLER_121_1371 ();
 sg13g2_decap_8 FILLER_121_1378 ();
 sg13g2_decap_8 FILLER_121_1385 ();
 sg13g2_decap_8 FILLER_121_1392 ();
 sg13g2_decap_8 FILLER_121_1399 ();
 sg13g2_decap_8 FILLER_121_1406 ();
 sg13g2_decap_8 FILLER_121_1413 ();
 sg13g2_decap_8 FILLER_121_1420 ();
 sg13g2_decap_8 FILLER_121_1427 ();
 sg13g2_decap_8 FILLER_121_1434 ();
 sg13g2_decap_8 FILLER_121_1441 ();
 sg13g2_decap_8 FILLER_121_1448 ();
 sg13g2_decap_8 FILLER_121_1455 ();
 sg13g2_decap_8 FILLER_121_1462 ();
 sg13g2_decap_8 FILLER_121_1469 ();
 sg13g2_decap_8 FILLER_121_1476 ();
 sg13g2_decap_8 FILLER_121_1483 ();
 sg13g2_decap_8 FILLER_121_1490 ();
 sg13g2_decap_8 FILLER_121_1497 ();
 sg13g2_decap_8 FILLER_121_1504 ();
 sg13g2_decap_8 FILLER_121_1511 ();
 sg13g2_decap_8 FILLER_121_1518 ();
 sg13g2_decap_8 FILLER_121_1525 ();
 sg13g2_decap_8 FILLER_121_1532 ();
 sg13g2_decap_8 FILLER_121_1539 ();
 sg13g2_decap_8 FILLER_121_1546 ();
 sg13g2_decap_8 FILLER_121_1553 ();
 sg13g2_decap_8 FILLER_121_1560 ();
 sg13g2_decap_8 FILLER_121_1567 ();
 sg13g2_decap_8 FILLER_121_1574 ();
 sg13g2_decap_8 FILLER_121_1581 ();
 sg13g2_decap_8 FILLER_121_1588 ();
 sg13g2_decap_8 FILLER_121_1595 ();
 sg13g2_decap_8 FILLER_121_1602 ();
 sg13g2_decap_8 FILLER_121_1609 ();
 sg13g2_decap_8 FILLER_121_1616 ();
 sg13g2_fill_2 FILLER_121_1623 ();
 sg13g2_decap_8 FILLER_122_0 ();
 sg13g2_decap_8 FILLER_122_7 ();
 sg13g2_fill_2 FILLER_122_14 ();
 sg13g2_decap_8 FILLER_122_20 ();
 sg13g2_decap_8 FILLER_122_27 ();
 sg13g2_decap_8 FILLER_122_34 ();
 sg13g2_decap_8 FILLER_122_41 ();
 sg13g2_decap_8 FILLER_122_48 ();
 sg13g2_decap_8 FILLER_122_55 ();
 sg13g2_decap_8 FILLER_122_62 ();
 sg13g2_fill_1 FILLER_122_69 ();
 sg13g2_fill_1 FILLER_122_95 ();
 sg13g2_decap_8 FILLER_122_108 ();
 sg13g2_decap_4 FILLER_122_120 ();
 sg13g2_fill_1 FILLER_122_124 ();
 sg13g2_fill_1 FILLER_122_156 ();
 sg13g2_fill_1 FILLER_122_162 ();
 sg13g2_decap_8 FILLER_122_168 ();
 sg13g2_decap_4 FILLER_122_175 ();
 sg13g2_fill_2 FILLER_122_179 ();
 sg13g2_decap_8 FILLER_122_207 ();
 sg13g2_decap_8 FILLER_122_214 ();
 sg13g2_decap_8 FILLER_122_221 ();
 sg13g2_fill_2 FILLER_122_228 ();
 sg13g2_decap_8 FILLER_122_242 ();
 sg13g2_decap_8 FILLER_122_249 ();
 sg13g2_decap_8 FILLER_122_256 ();
 sg13g2_fill_1 FILLER_122_263 ();
 sg13g2_decap_8 FILLER_122_268 ();
 sg13g2_decap_8 FILLER_122_275 ();
 sg13g2_fill_1 FILLER_122_282 ();
 sg13g2_fill_2 FILLER_122_329 ();
 sg13g2_decap_4 FILLER_122_357 ();
 sg13g2_fill_1 FILLER_122_361 ();
 sg13g2_decap_8 FILLER_122_367 ();
 sg13g2_decap_8 FILLER_122_374 ();
 sg13g2_decap_4 FILLER_122_387 ();
 sg13g2_fill_1 FILLER_122_391 ();
 sg13g2_decap_8 FILLER_122_397 ();
 sg13g2_decap_8 FILLER_122_404 ();
 sg13g2_fill_1 FILLER_122_411 ();
 sg13g2_decap_8 FILLER_122_424 ();
 sg13g2_decap_8 FILLER_122_431 ();
 sg13g2_decap_4 FILLER_122_438 ();
 sg13g2_fill_2 FILLER_122_442 ();
 sg13g2_decap_8 FILLER_122_499 ();
 sg13g2_fill_1 FILLER_122_506 ();
 sg13g2_decap_8 FILLER_122_511 ();
 sg13g2_fill_2 FILLER_122_518 ();
 sg13g2_fill_1 FILLER_122_528 ();
 sg13g2_decap_4 FILLER_122_564 ();
 sg13g2_decap_8 FILLER_122_594 ();
 sg13g2_fill_2 FILLER_122_601 ();
 sg13g2_decap_8 FILLER_122_607 ();
 sg13g2_decap_4 FILLER_122_614 ();
 sg13g2_fill_2 FILLER_122_648 ();
 sg13g2_fill_1 FILLER_122_650 ();
 sg13g2_decap_4 FILLER_122_690 ();
 sg13g2_fill_1 FILLER_122_694 ();
 sg13g2_decap_4 FILLER_122_704 ();
 sg13g2_fill_2 FILLER_122_708 ();
 sg13g2_decap_8 FILLER_122_719 ();
 sg13g2_fill_1 FILLER_122_726 ();
 sg13g2_fill_1 FILLER_122_734 ();
 sg13g2_fill_2 FILLER_122_739 ();
 sg13g2_decap_4 FILLER_122_756 ();
 sg13g2_fill_1 FILLER_122_760 ();
 sg13g2_decap_4 FILLER_122_773 ();
 sg13g2_decap_4 FILLER_122_785 ();
 sg13g2_decap_8 FILLER_122_799 ();
 sg13g2_decap_4 FILLER_122_806 ();
 sg13g2_fill_1 FILLER_122_810 ();
 sg13g2_decap_8 FILLER_122_826 ();
 sg13g2_decap_8 FILLER_122_833 ();
 sg13g2_fill_2 FILLER_122_840 ();
 sg13g2_fill_1 FILLER_122_842 ();
 sg13g2_fill_1 FILLER_122_848 ();
 sg13g2_fill_2 FILLER_122_853 ();
 sg13g2_fill_1 FILLER_122_855 ();
 sg13g2_decap_8 FILLER_122_864 ();
 sg13g2_decap_8 FILLER_122_871 ();
 sg13g2_decap_4 FILLER_122_878 ();
 sg13g2_decap_8 FILLER_122_891 ();
 sg13g2_decap_4 FILLER_122_903 ();
 sg13g2_fill_2 FILLER_122_907 ();
 sg13g2_fill_1 FILLER_122_918 ();
 sg13g2_decap_4 FILLER_122_922 ();
 sg13g2_fill_2 FILLER_122_926 ();
 sg13g2_fill_2 FILLER_122_933 ();
 sg13g2_fill_1 FILLER_122_935 ();
 sg13g2_fill_1 FILLER_122_944 ();
 sg13g2_fill_2 FILLER_122_983 ();
 sg13g2_decap_8 FILLER_122_992 ();
 sg13g2_decap_8 FILLER_122_999 ();
 sg13g2_decap_8 FILLER_122_1006 ();
 sg13g2_fill_1 FILLER_122_1013 ();
 sg13g2_fill_1 FILLER_122_1024 ();
 sg13g2_decap_4 FILLER_122_1039 ();
 sg13g2_fill_2 FILLER_122_1064 ();
 sg13g2_fill_1 FILLER_122_1066 ();
 sg13g2_decap_4 FILLER_122_1079 ();
 sg13g2_fill_2 FILLER_122_1083 ();
 sg13g2_decap_8 FILLER_122_1111 ();
 sg13g2_decap_8 FILLER_122_1118 ();
 sg13g2_decap_8 FILLER_122_1125 ();
 sg13g2_decap_8 FILLER_122_1132 ();
 sg13g2_decap_8 FILLER_122_1139 ();
 sg13g2_fill_2 FILLER_122_1146 ();
 sg13g2_decap_8 FILLER_122_1153 ();
 sg13g2_decap_8 FILLER_122_1160 ();
 sg13g2_decap_8 FILLER_122_1167 ();
 sg13g2_decap_8 FILLER_122_1174 ();
 sg13g2_decap_8 FILLER_122_1181 ();
 sg13g2_decap_4 FILLER_122_1188 ();
 sg13g2_fill_1 FILLER_122_1192 ();
 sg13g2_decap_8 FILLER_122_1204 ();
 sg13g2_decap_8 FILLER_122_1211 ();
 sg13g2_fill_2 FILLER_122_1218 ();
 sg13g2_fill_1 FILLER_122_1220 ();
 sg13g2_decap_8 FILLER_122_1232 ();
 sg13g2_fill_1 FILLER_122_1239 ();
 sg13g2_fill_1 FILLER_122_1261 ();
 sg13g2_decap_8 FILLER_122_1267 ();
 sg13g2_fill_1 FILLER_122_1274 ();
 sg13g2_decap_8 FILLER_122_1279 ();
 sg13g2_fill_2 FILLER_122_1286 ();
 sg13g2_fill_1 FILLER_122_1288 ();
 sg13g2_fill_2 FILLER_122_1299 ();
 sg13g2_fill_1 FILLER_122_1306 ();
 sg13g2_fill_2 FILLER_122_1316 ();
 sg13g2_fill_1 FILLER_122_1318 ();
 sg13g2_fill_2 FILLER_122_1328 ();
 sg13g2_fill_1 FILLER_122_1346 ();
 sg13g2_decap_8 FILLER_122_1352 ();
 sg13g2_decap_8 FILLER_122_1359 ();
 sg13g2_decap_4 FILLER_122_1366 ();
 sg13g2_decap_4 FILLER_122_1375 ();
 sg13g2_fill_2 FILLER_122_1379 ();
 sg13g2_decap_8 FILLER_122_1385 ();
 sg13g2_decap_8 FILLER_122_1392 ();
 sg13g2_decap_8 FILLER_122_1399 ();
 sg13g2_decap_8 FILLER_122_1406 ();
 sg13g2_decap_8 FILLER_122_1413 ();
 sg13g2_decap_8 FILLER_122_1420 ();
 sg13g2_decap_8 FILLER_122_1427 ();
 sg13g2_decap_8 FILLER_122_1434 ();
 sg13g2_decap_8 FILLER_122_1441 ();
 sg13g2_decap_8 FILLER_122_1448 ();
 sg13g2_decap_8 FILLER_122_1455 ();
 sg13g2_decap_8 FILLER_122_1462 ();
 sg13g2_decap_8 FILLER_122_1469 ();
 sg13g2_decap_8 FILLER_122_1476 ();
 sg13g2_decap_8 FILLER_122_1483 ();
 sg13g2_decap_8 FILLER_122_1490 ();
 sg13g2_decap_8 FILLER_122_1497 ();
 sg13g2_decap_8 FILLER_122_1504 ();
 sg13g2_decap_8 FILLER_122_1511 ();
 sg13g2_decap_8 FILLER_122_1518 ();
 sg13g2_decap_8 FILLER_122_1525 ();
 sg13g2_decap_8 FILLER_122_1532 ();
 sg13g2_decap_8 FILLER_122_1539 ();
 sg13g2_decap_8 FILLER_122_1546 ();
 sg13g2_decap_8 FILLER_122_1553 ();
 sg13g2_decap_8 FILLER_122_1560 ();
 sg13g2_decap_8 FILLER_122_1567 ();
 sg13g2_decap_8 FILLER_122_1574 ();
 sg13g2_decap_8 FILLER_122_1581 ();
 sg13g2_decap_8 FILLER_122_1588 ();
 sg13g2_decap_8 FILLER_122_1595 ();
 sg13g2_decap_8 FILLER_122_1602 ();
 sg13g2_decap_8 FILLER_122_1609 ();
 sg13g2_decap_8 FILLER_122_1616 ();
 sg13g2_fill_2 FILLER_122_1623 ();
 sg13g2_decap_8 FILLER_123_0 ();
 sg13g2_fill_2 FILLER_123_7 ();
 sg13g2_fill_1 FILLER_123_9 ();
 sg13g2_decap_8 FILLER_123_36 ();
 sg13g2_decap_8 FILLER_123_43 ();
 sg13g2_fill_1 FILLER_123_50 ();
 sg13g2_decap_4 FILLER_123_55 ();
 sg13g2_fill_2 FILLER_123_97 ();
 sg13g2_fill_1 FILLER_123_99 ();
 sg13g2_fill_1 FILLER_123_105 ();
 sg13g2_decap_4 FILLER_123_116 ();
 sg13g2_fill_1 FILLER_123_120 ();
 sg13g2_decap_8 FILLER_123_131 ();
 sg13g2_decap_8 FILLER_123_138 ();
 sg13g2_decap_4 FILLER_123_150 ();
 sg13g2_fill_1 FILLER_123_154 ();
 sg13g2_decap_8 FILLER_123_167 ();
 sg13g2_decap_8 FILLER_123_174 ();
 sg13g2_decap_8 FILLER_123_181 ();
 sg13g2_fill_2 FILLER_123_188 ();
 sg13g2_decap_8 FILLER_123_215 ();
 sg13g2_decap_4 FILLER_123_222 ();
 sg13g2_fill_1 FILLER_123_226 ();
 sg13g2_fill_1 FILLER_123_254 ();
 sg13g2_decap_4 FILLER_123_281 ();
 sg13g2_fill_2 FILLER_123_304 ();
 sg13g2_fill_1 FILLER_123_306 ();
 sg13g2_fill_2 FILLER_123_312 ();
 sg13g2_fill_1 FILLER_123_314 ();
 sg13g2_fill_2 FILLER_123_320 ();
 sg13g2_decap_8 FILLER_123_331 ();
 sg13g2_decap_8 FILLER_123_338 ();
 sg13g2_decap_4 FILLER_123_345 ();
 sg13g2_fill_1 FILLER_123_349 ();
 sg13g2_decap_8 FILLER_123_359 ();
 sg13g2_fill_1 FILLER_123_366 ();
 sg13g2_decap_8 FILLER_123_372 ();
 sg13g2_decap_8 FILLER_123_379 ();
 sg13g2_decap_8 FILLER_123_386 ();
 sg13g2_decap_8 FILLER_123_393 ();
 sg13g2_decap_8 FILLER_123_400 ();
 sg13g2_fill_2 FILLER_123_407 ();
 sg13g2_fill_2 FILLER_123_413 ();
 sg13g2_decap_8 FILLER_123_433 ();
 sg13g2_decap_8 FILLER_123_440 ();
 sg13g2_fill_2 FILLER_123_447 ();
 sg13g2_fill_1 FILLER_123_454 ();
 sg13g2_fill_1 FILLER_123_467 ();
 sg13g2_fill_2 FILLER_123_474 ();
 sg13g2_fill_1 FILLER_123_476 ();
 sg13g2_decap_8 FILLER_123_488 ();
 sg13g2_decap_4 FILLER_123_495 ();
 sg13g2_fill_1 FILLER_123_499 ();
 sg13g2_decap_8 FILLER_123_504 ();
 sg13g2_decap_8 FILLER_123_511 ();
 sg13g2_decap_8 FILLER_123_518 ();
 sg13g2_decap_8 FILLER_123_525 ();
 sg13g2_decap_8 FILLER_123_532 ();
 sg13g2_fill_1 FILLER_123_539 ();
 sg13g2_decap_8 FILLER_123_558 ();
 sg13g2_decap_8 FILLER_123_565 ();
 sg13g2_fill_2 FILLER_123_572 ();
 sg13g2_fill_2 FILLER_123_583 ();
 sg13g2_fill_1 FILLER_123_585 ();
 sg13g2_fill_2 FILLER_123_590 ();
 sg13g2_fill_2 FILLER_123_646 ();
 sg13g2_fill_2 FILLER_123_681 ();
 sg13g2_fill_1 FILLER_123_683 ();
 sg13g2_fill_2 FILLER_123_689 ();
 sg13g2_decap_8 FILLER_123_699 ();
 sg13g2_fill_1 FILLER_123_706 ();
 sg13g2_decap_4 FILLER_123_711 ();
 sg13g2_decap_4 FILLER_123_723 ();
 sg13g2_fill_2 FILLER_123_731 ();
 sg13g2_fill_1 FILLER_123_733 ();
 sg13g2_fill_1 FILLER_123_742 ();
 sg13g2_fill_1 FILLER_123_748 ();
 sg13g2_decap_4 FILLER_123_761 ();
 sg13g2_fill_2 FILLER_123_768 ();
 sg13g2_fill_1 FILLER_123_770 ();
 sg13g2_decap_8 FILLER_123_776 ();
 sg13g2_fill_2 FILLER_123_783 ();
 sg13g2_fill_1 FILLER_123_785 ();
 sg13g2_fill_2 FILLER_123_799 ();
 sg13g2_fill_2 FILLER_123_809 ();
 sg13g2_decap_8 FILLER_123_826 ();
 sg13g2_decap_8 FILLER_123_833 ();
 sg13g2_fill_1 FILLER_123_844 ();
 sg13g2_decap_8 FILLER_123_849 ();
 sg13g2_decap_8 FILLER_123_856 ();
 sg13g2_decap_4 FILLER_123_870 ();
 sg13g2_fill_1 FILLER_123_874 ();
 sg13g2_decap_8 FILLER_123_888 ();
 sg13g2_decap_8 FILLER_123_895 ();
 sg13g2_fill_1 FILLER_123_902 ();
 sg13g2_fill_2 FILLER_123_908 ();
 sg13g2_fill_1 FILLER_123_910 ();
 sg13g2_decap_4 FILLER_123_921 ();
 sg13g2_fill_2 FILLER_123_972 ();
 sg13g2_decap_4 FILLER_123_991 ();
 sg13g2_fill_2 FILLER_123_995 ();
 sg13g2_decap_8 FILLER_123_1001 ();
 sg13g2_decap_8 FILLER_123_1008 ();
 sg13g2_decap_4 FILLER_123_1015 ();
 sg13g2_fill_2 FILLER_123_1027 ();
 sg13g2_fill_1 FILLER_123_1029 ();
 sg13g2_fill_1 FILLER_123_1045 ();
 sg13g2_fill_1 FILLER_123_1051 ();
 sg13g2_fill_1 FILLER_123_1060 ();
 sg13g2_fill_2 FILLER_123_1066 ();
 sg13g2_decap_4 FILLER_123_1074 ();
 sg13g2_fill_2 FILLER_123_1078 ();
 sg13g2_decap_8 FILLER_123_1088 ();
 sg13g2_decap_4 FILLER_123_1095 ();
 sg13g2_fill_2 FILLER_123_1099 ();
 sg13g2_decap_8 FILLER_123_1118 ();
 sg13g2_fill_1 FILLER_123_1125 ();
 sg13g2_decap_8 FILLER_123_1134 ();
 sg13g2_fill_1 FILLER_123_1141 ();
 sg13g2_decap_8 FILLER_123_1153 ();
 sg13g2_decap_8 FILLER_123_1160 ();
 sg13g2_fill_2 FILLER_123_1167 ();
 sg13g2_fill_1 FILLER_123_1173 ();
 sg13g2_decap_8 FILLER_123_1180 ();
 sg13g2_fill_1 FILLER_123_1187 ();
 sg13g2_fill_2 FILLER_123_1204 ();
 sg13g2_decap_8 FILLER_123_1216 ();
 sg13g2_fill_2 FILLER_123_1223 ();
 sg13g2_fill_1 FILLER_123_1237 ();
 sg13g2_decap_4 FILLER_123_1257 ();
 sg13g2_decap_8 FILLER_123_1265 ();
 sg13g2_fill_1 FILLER_123_1272 ();
 sg13g2_decap_4 FILLER_123_1277 ();
 sg13g2_decap_8 FILLER_123_1313 ();
 sg13g2_decap_4 FILLER_123_1320 ();
 sg13g2_decap_8 FILLER_123_1329 ();
 sg13g2_fill_2 FILLER_123_1344 ();
 sg13g2_fill_1 FILLER_123_1346 ();
 sg13g2_fill_1 FILLER_123_1365 ();
 sg13g2_decap_4 FILLER_123_1369 ();
 sg13g2_decap_8 FILLER_123_1399 ();
 sg13g2_decap_8 FILLER_123_1406 ();
 sg13g2_decap_8 FILLER_123_1413 ();
 sg13g2_decap_8 FILLER_123_1420 ();
 sg13g2_decap_8 FILLER_123_1427 ();
 sg13g2_decap_8 FILLER_123_1434 ();
 sg13g2_decap_8 FILLER_123_1441 ();
 sg13g2_decap_8 FILLER_123_1448 ();
 sg13g2_decap_8 FILLER_123_1455 ();
 sg13g2_decap_8 FILLER_123_1462 ();
 sg13g2_decap_8 FILLER_123_1469 ();
 sg13g2_decap_8 FILLER_123_1476 ();
 sg13g2_decap_8 FILLER_123_1483 ();
 sg13g2_decap_8 FILLER_123_1490 ();
 sg13g2_decap_8 FILLER_123_1497 ();
 sg13g2_decap_8 FILLER_123_1504 ();
 sg13g2_decap_8 FILLER_123_1511 ();
 sg13g2_decap_8 FILLER_123_1518 ();
 sg13g2_decap_8 FILLER_123_1525 ();
 sg13g2_decap_8 FILLER_123_1532 ();
 sg13g2_decap_8 FILLER_123_1539 ();
 sg13g2_decap_8 FILLER_123_1546 ();
 sg13g2_decap_8 FILLER_123_1553 ();
 sg13g2_decap_8 FILLER_123_1560 ();
 sg13g2_decap_8 FILLER_123_1567 ();
 sg13g2_decap_8 FILLER_123_1574 ();
 sg13g2_decap_8 FILLER_123_1581 ();
 sg13g2_decap_8 FILLER_123_1588 ();
 sg13g2_decap_8 FILLER_123_1595 ();
 sg13g2_decap_8 FILLER_123_1602 ();
 sg13g2_decap_8 FILLER_123_1609 ();
 sg13g2_decap_8 FILLER_123_1616 ();
 sg13g2_fill_2 FILLER_123_1623 ();
 sg13g2_decap_8 FILLER_124_0 ();
 sg13g2_fill_2 FILLER_124_11 ();
 sg13g2_fill_1 FILLER_124_13 ();
 sg13g2_fill_2 FILLER_124_40 ();
 sg13g2_decap_8 FILLER_124_46 ();
 sg13g2_decap_4 FILLER_124_53 ();
 sg13g2_fill_1 FILLER_124_57 ();
 sg13g2_decap_4 FILLER_124_97 ();
 sg13g2_fill_1 FILLER_124_106 ();
 sg13g2_decap_8 FILLER_124_112 ();
 sg13g2_decap_8 FILLER_124_119 ();
 sg13g2_fill_1 FILLER_124_126 ();
 sg13g2_decap_4 FILLER_124_137 ();
 sg13g2_fill_1 FILLER_124_141 ();
 sg13g2_fill_2 FILLER_124_152 ();
 sg13g2_fill_1 FILLER_124_154 ();
 sg13g2_decap_4 FILLER_124_160 ();
 sg13g2_fill_2 FILLER_124_189 ();
 sg13g2_fill_1 FILLER_124_191 ();
 sg13g2_fill_2 FILLER_124_201 ();
 sg13g2_decap_8 FILLER_124_208 ();
 sg13g2_fill_2 FILLER_124_215 ();
 sg13g2_fill_1 FILLER_124_217 ();
 sg13g2_decap_4 FILLER_124_227 ();
 sg13g2_fill_1 FILLER_124_231 ();
 sg13g2_decap_8 FILLER_124_237 ();
 sg13g2_fill_1 FILLER_124_244 ();
 sg13g2_decap_8 FILLER_124_250 ();
 sg13g2_decap_8 FILLER_124_257 ();
 sg13g2_decap_8 FILLER_124_264 ();
 sg13g2_decap_8 FILLER_124_271 ();
 sg13g2_decap_4 FILLER_124_278 ();
 sg13g2_fill_2 FILLER_124_310 ();
 sg13g2_fill_2 FILLER_124_337 ();
 sg13g2_decap_4 FILLER_124_343 ();
 sg13g2_fill_2 FILLER_124_347 ();
 sg13g2_decap_8 FILLER_124_358 ();
 sg13g2_fill_2 FILLER_124_365 ();
 sg13g2_fill_2 FILLER_124_372 ();
 sg13g2_fill_1 FILLER_124_374 ();
 sg13g2_decap_8 FILLER_124_384 ();
 sg13g2_fill_1 FILLER_124_397 ();
 sg13g2_decap_8 FILLER_124_402 ();
 sg13g2_decap_8 FILLER_124_414 ();
 sg13g2_decap_4 FILLER_124_421 ();
 sg13g2_fill_2 FILLER_124_425 ();
 sg13g2_decap_4 FILLER_124_440 ();
 sg13g2_fill_2 FILLER_124_444 ();
 sg13g2_fill_1 FILLER_124_466 ();
 sg13g2_decap_8 FILLER_124_472 ();
 sg13g2_decap_8 FILLER_124_479 ();
 sg13g2_fill_2 FILLER_124_486 ();
 sg13g2_fill_2 FILLER_124_519 ();
 sg13g2_fill_2 FILLER_124_565 ();
 sg13g2_decap_4 FILLER_124_626 ();
 sg13g2_decap_8 FILLER_124_691 ();
 sg13g2_decap_4 FILLER_124_698 ();
 sg13g2_fill_2 FILLER_124_702 ();
 sg13g2_decap_8 FILLER_124_716 ();
 sg13g2_decap_8 FILLER_124_723 ();
 sg13g2_decap_8 FILLER_124_730 ();
 sg13g2_decap_8 FILLER_124_737 ();
 sg13g2_decap_8 FILLER_124_744 ();
 sg13g2_decap_4 FILLER_124_761 ();
 sg13g2_fill_2 FILLER_124_770 ();
 sg13g2_decap_8 FILLER_124_776 ();
 sg13g2_fill_2 FILLER_124_783 ();
 sg13g2_fill_1 FILLER_124_790 ();
 sg13g2_fill_1 FILLER_124_795 ();
 sg13g2_decap_8 FILLER_124_802 ();
 sg13g2_decap_4 FILLER_124_809 ();
 sg13g2_fill_2 FILLER_124_813 ();
 sg13g2_decap_8 FILLER_124_826 ();
 sg13g2_decap_4 FILLER_124_833 ();
 sg13g2_decap_8 FILLER_124_862 ();
 sg13g2_decap_8 FILLER_124_869 ();
 sg13g2_decap_4 FILLER_124_876 ();
 sg13g2_decap_8 FILLER_124_885 ();
 sg13g2_fill_1 FILLER_124_892 ();
 sg13g2_decap_8 FILLER_124_898 ();
 sg13g2_decap_8 FILLER_124_905 ();
 sg13g2_decap_8 FILLER_124_912 ();
 sg13g2_decap_4 FILLER_124_919 ();
 sg13g2_fill_2 FILLER_124_923 ();
 sg13g2_fill_2 FILLER_124_931 ();
 sg13g2_decap_4 FILLER_124_939 ();
 sg13g2_fill_1 FILLER_124_943 ();
 sg13g2_decap_8 FILLER_124_951 ();
 sg13g2_decap_8 FILLER_124_958 ();
 sg13g2_decap_4 FILLER_124_965 ();
 sg13g2_decap_4 FILLER_124_974 ();
 sg13g2_decap_4 FILLER_124_986 ();
 sg13g2_decap_8 FILLER_124_1016 ();
 sg13g2_decap_8 FILLER_124_1029 ();
 sg13g2_decap_8 FILLER_124_1036 ();
 sg13g2_decap_4 FILLER_124_1043 ();
 sg13g2_fill_2 FILLER_124_1065 ();
 sg13g2_fill_1 FILLER_124_1067 ();
 sg13g2_fill_1 FILLER_124_1079 ();
 sg13g2_decap_8 FILLER_124_1085 ();
 sg13g2_decap_8 FILLER_124_1092 ();
 sg13g2_fill_2 FILLER_124_1099 ();
 sg13g2_decap_4 FILLER_124_1104 ();
 sg13g2_decap_8 FILLER_124_1112 ();
 sg13g2_decap_4 FILLER_124_1119 ();
 sg13g2_fill_1 FILLER_124_1123 ();
 sg13g2_decap_8 FILLER_124_1146 ();
 sg13g2_fill_2 FILLER_124_1153 ();
 sg13g2_fill_1 FILLER_124_1155 ();
 sg13g2_fill_2 FILLER_124_1160 ();
 sg13g2_fill_1 FILLER_124_1193 ();
 sg13g2_decap_4 FILLER_124_1200 ();
 sg13g2_fill_2 FILLER_124_1204 ();
 sg13g2_fill_2 FILLER_124_1214 ();
 sg13g2_fill_1 FILLER_124_1221 ();
 sg13g2_fill_2 FILLER_124_1226 ();
 sg13g2_decap_4 FILLER_124_1233 ();
 sg13g2_fill_1 FILLER_124_1237 ();
 sg13g2_decap_8 FILLER_124_1243 ();
 sg13g2_decap_8 FILLER_124_1250 ();
 sg13g2_fill_2 FILLER_124_1262 ();
 sg13g2_fill_2 FILLER_124_1271 ();
 sg13g2_fill_1 FILLER_124_1273 ();
 sg13g2_fill_2 FILLER_124_1294 ();
 sg13g2_fill_1 FILLER_124_1296 ();
 sg13g2_fill_1 FILLER_124_1301 ();
 sg13g2_decap_8 FILLER_124_1310 ();
 sg13g2_decap_4 FILLER_124_1317 ();
 sg13g2_decap_4 FILLER_124_1335 ();
 sg13g2_fill_1 FILLER_124_1350 ();
 sg13g2_decap_8 FILLER_124_1363 ();
 sg13g2_decap_4 FILLER_124_1370 ();
 sg13g2_fill_1 FILLER_124_1374 ();
 sg13g2_decap_8 FILLER_124_1380 ();
 sg13g2_decap_8 FILLER_124_1387 ();
 sg13g2_decap_8 FILLER_124_1394 ();
 sg13g2_decap_8 FILLER_124_1401 ();
 sg13g2_decap_8 FILLER_124_1408 ();
 sg13g2_decap_8 FILLER_124_1415 ();
 sg13g2_decap_8 FILLER_124_1422 ();
 sg13g2_decap_8 FILLER_124_1429 ();
 sg13g2_decap_8 FILLER_124_1436 ();
 sg13g2_decap_8 FILLER_124_1443 ();
 sg13g2_decap_8 FILLER_124_1450 ();
 sg13g2_decap_8 FILLER_124_1457 ();
 sg13g2_decap_8 FILLER_124_1464 ();
 sg13g2_decap_8 FILLER_124_1471 ();
 sg13g2_decap_8 FILLER_124_1478 ();
 sg13g2_decap_8 FILLER_124_1485 ();
 sg13g2_decap_8 FILLER_124_1492 ();
 sg13g2_decap_8 FILLER_124_1499 ();
 sg13g2_decap_8 FILLER_124_1506 ();
 sg13g2_decap_8 FILLER_124_1513 ();
 sg13g2_decap_8 FILLER_124_1520 ();
 sg13g2_decap_8 FILLER_124_1527 ();
 sg13g2_decap_8 FILLER_124_1534 ();
 sg13g2_decap_8 FILLER_124_1541 ();
 sg13g2_decap_8 FILLER_124_1548 ();
 sg13g2_decap_8 FILLER_124_1555 ();
 sg13g2_decap_8 FILLER_124_1562 ();
 sg13g2_decap_8 FILLER_124_1569 ();
 sg13g2_decap_8 FILLER_124_1576 ();
 sg13g2_decap_8 FILLER_124_1583 ();
 sg13g2_decap_8 FILLER_124_1590 ();
 sg13g2_decap_8 FILLER_124_1597 ();
 sg13g2_decap_8 FILLER_124_1604 ();
 sg13g2_decap_8 FILLER_124_1611 ();
 sg13g2_decap_8 FILLER_124_1618 ();
 sg13g2_decap_8 FILLER_125_0 ();
 sg13g2_decap_4 FILLER_125_7 ();
 sg13g2_fill_2 FILLER_125_11 ();
 sg13g2_fill_1 FILLER_125_17 ();
 sg13g2_decap_4 FILLER_125_22 ();
 sg13g2_fill_2 FILLER_125_30 ();
 sg13g2_fill_1 FILLER_125_32 ();
 sg13g2_fill_1 FILLER_125_59 ();
 sg13g2_fill_2 FILLER_125_86 ();
 sg13g2_fill_1 FILLER_125_93 ();
 sg13g2_fill_1 FILLER_125_99 ();
 sg13g2_fill_1 FILLER_125_105 ();
 sg13g2_fill_1 FILLER_125_113 ();
 sg13g2_fill_2 FILLER_125_119 ();
 sg13g2_fill_1 FILLER_125_126 ();
 sg13g2_fill_2 FILLER_125_132 ();
 sg13g2_fill_2 FILLER_125_144 ();
 sg13g2_fill_1 FILLER_125_146 ();
 sg13g2_fill_2 FILLER_125_152 ();
 sg13g2_fill_2 FILLER_125_164 ();
 sg13g2_fill_1 FILLER_125_166 ();
 sg13g2_decap_4 FILLER_125_172 ();
 sg13g2_fill_2 FILLER_125_176 ();
 sg13g2_fill_2 FILLER_125_185 ();
 sg13g2_fill_2 FILLER_125_213 ();
 sg13g2_fill_1 FILLER_125_215 ();
 sg13g2_fill_1 FILLER_125_242 ();
 sg13g2_decap_4 FILLER_125_258 ();
 sg13g2_fill_2 FILLER_125_262 ();
 sg13g2_decap_4 FILLER_125_269 ();
 sg13g2_fill_1 FILLER_125_273 ();
 sg13g2_fill_2 FILLER_125_283 ();
 sg13g2_fill_2 FILLER_125_311 ();
 sg13g2_decap_8 FILLER_125_319 ();
 sg13g2_decap_4 FILLER_125_326 ();
 sg13g2_fill_1 FILLER_125_330 ();
 sg13g2_decap_8 FILLER_125_341 ();
 sg13g2_decap_8 FILLER_125_360 ();
 sg13g2_decap_8 FILLER_125_367 ();
 sg13g2_decap_8 FILLER_125_411 ();
 sg13g2_fill_2 FILLER_125_418 ();
 sg13g2_fill_1 FILLER_125_425 ();
 sg13g2_fill_2 FILLER_125_441 ();
 sg13g2_decap_8 FILLER_125_465 ();
 sg13g2_decap_4 FILLER_125_472 ();
 sg13g2_fill_1 FILLER_125_476 ();
 sg13g2_fill_1 FILLER_125_482 ();
 sg13g2_decap_8 FILLER_125_488 ();
 sg13g2_decap_8 FILLER_125_495 ();
 sg13g2_fill_2 FILLER_125_502 ();
 sg13g2_decap_4 FILLER_125_559 ();
 sg13g2_fill_1 FILLER_125_563 ();
 sg13g2_fill_1 FILLER_125_625 ();
 sg13g2_decap_8 FILLER_125_630 ();
 sg13g2_decap_4 FILLER_125_670 ();
 sg13g2_fill_2 FILLER_125_674 ();
 sg13g2_decap_4 FILLER_125_706 ();
 sg13g2_decap_4 FILLER_125_724 ();
 sg13g2_fill_2 FILLER_125_741 ();
 sg13g2_fill_1 FILLER_125_743 ();
 sg13g2_decap_8 FILLER_125_749 ();
 sg13g2_decap_4 FILLER_125_781 ();
 sg13g2_fill_2 FILLER_125_785 ();
 sg13g2_decap_8 FILLER_125_822 ();
 sg13g2_decap_8 FILLER_125_829 ();
 sg13g2_fill_2 FILLER_125_836 ();
 sg13g2_fill_1 FILLER_125_838 ();
 sg13g2_fill_2 FILLER_125_847 ();
 sg13g2_decap_4 FILLER_125_858 ();
 sg13g2_decap_4 FILLER_125_868 ();
 sg13g2_fill_1 FILLER_125_893 ();
 sg13g2_decap_8 FILLER_125_920 ();
 sg13g2_decap_4 FILLER_125_927 ();
 sg13g2_fill_1 FILLER_125_931 ();
 sg13g2_decap_8 FILLER_125_944 ();
 sg13g2_decap_8 FILLER_125_951 ();
 sg13g2_fill_1 FILLER_125_958 ();
 sg13g2_decap_8 FILLER_125_963 ();
 sg13g2_fill_2 FILLER_125_970 ();
 sg13g2_decap_8 FILLER_125_1032 ();
 sg13g2_decap_8 FILLER_125_1039 ();
 sg13g2_decap_8 FILLER_125_1046 ();
 sg13g2_decap_8 FILLER_125_1053 ();
 sg13g2_fill_2 FILLER_125_1060 ();
 sg13g2_decap_8 FILLER_125_1070 ();
 sg13g2_fill_2 FILLER_125_1127 ();
 sg13g2_decap_8 FILLER_125_1134 ();
 sg13g2_decap_8 FILLER_125_1141 ();
 sg13g2_decap_8 FILLER_125_1148 ();
 sg13g2_decap_8 FILLER_125_1155 ();
 sg13g2_decap_4 FILLER_125_1162 ();
 sg13g2_fill_2 FILLER_125_1166 ();
 sg13g2_decap_8 FILLER_125_1173 ();
 sg13g2_decap_4 FILLER_125_1180 ();
 sg13g2_fill_1 FILLER_125_1197 ();
 sg13g2_fill_1 FILLER_125_1203 ();
 sg13g2_fill_1 FILLER_125_1211 ();
 sg13g2_fill_2 FILLER_125_1217 ();
 sg13g2_decap_8 FILLER_125_1234 ();
 sg13g2_decap_8 FILLER_125_1241 ();
 sg13g2_decap_8 FILLER_125_1248 ();
 sg13g2_fill_2 FILLER_125_1255 ();
 sg13g2_fill_1 FILLER_125_1257 ();
 sg13g2_decap_8 FILLER_125_1265 ();
 sg13g2_decap_8 FILLER_125_1272 ();
 sg13g2_decap_8 FILLER_125_1279 ();
 sg13g2_fill_1 FILLER_125_1291 ();
 sg13g2_fill_2 FILLER_125_1302 ();
 sg13g2_fill_1 FILLER_125_1309 ();
 sg13g2_decap_8 FILLER_125_1315 ();
 sg13g2_fill_2 FILLER_125_1340 ();
 sg13g2_fill_1 FILLER_125_1353 ();
 sg13g2_decap_8 FILLER_125_1362 ();
 sg13g2_decap_8 FILLER_125_1369 ();
 sg13g2_decap_8 FILLER_125_1376 ();
 sg13g2_fill_1 FILLER_125_1383 ();
 sg13g2_decap_8 FILLER_125_1388 ();
 sg13g2_decap_8 FILLER_125_1395 ();
 sg13g2_decap_8 FILLER_125_1402 ();
 sg13g2_decap_8 FILLER_125_1409 ();
 sg13g2_decap_8 FILLER_125_1416 ();
 sg13g2_decap_8 FILLER_125_1423 ();
 sg13g2_decap_8 FILLER_125_1430 ();
 sg13g2_decap_8 FILLER_125_1437 ();
 sg13g2_decap_8 FILLER_125_1444 ();
 sg13g2_decap_8 FILLER_125_1451 ();
 sg13g2_decap_8 FILLER_125_1458 ();
 sg13g2_decap_8 FILLER_125_1465 ();
 sg13g2_decap_8 FILLER_125_1472 ();
 sg13g2_decap_8 FILLER_125_1479 ();
 sg13g2_decap_8 FILLER_125_1486 ();
 sg13g2_decap_8 FILLER_125_1493 ();
 sg13g2_decap_8 FILLER_125_1500 ();
 sg13g2_decap_8 FILLER_125_1507 ();
 sg13g2_decap_8 FILLER_125_1514 ();
 sg13g2_decap_8 FILLER_125_1521 ();
 sg13g2_decap_8 FILLER_125_1528 ();
 sg13g2_decap_8 FILLER_125_1535 ();
 sg13g2_decap_8 FILLER_125_1542 ();
 sg13g2_decap_8 FILLER_125_1549 ();
 sg13g2_decap_8 FILLER_125_1556 ();
 sg13g2_decap_8 FILLER_125_1563 ();
 sg13g2_decap_8 FILLER_125_1570 ();
 sg13g2_decap_8 FILLER_125_1577 ();
 sg13g2_decap_8 FILLER_125_1584 ();
 sg13g2_decap_8 FILLER_125_1591 ();
 sg13g2_decap_8 FILLER_125_1598 ();
 sg13g2_decap_8 FILLER_125_1605 ();
 sg13g2_decap_8 FILLER_125_1612 ();
 sg13g2_decap_4 FILLER_125_1619 ();
 sg13g2_fill_2 FILLER_125_1623 ();
 sg13g2_decap_8 FILLER_126_0 ();
 sg13g2_decap_8 FILLER_126_7 ();
 sg13g2_decap_8 FILLER_126_14 ();
 sg13g2_fill_2 FILLER_126_21 ();
 sg13g2_fill_1 FILLER_126_23 ();
 sg13g2_decap_8 FILLER_126_53 ();
 sg13g2_decap_4 FILLER_126_60 ();
 sg13g2_fill_1 FILLER_126_72 ();
 sg13g2_fill_2 FILLER_126_81 ();
 sg13g2_decap_4 FILLER_126_100 ();
 sg13g2_decap_4 FILLER_126_109 ();
 sg13g2_decap_4 FILLER_126_134 ();
 sg13g2_fill_1 FILLER_126_160 ();
 sg13g2_fill_1 FILLER_126_166 ();
 sg13g2_decap_8 FILLER_126_172 ();
 sg13g2_decap_4 FILLER_126_179 ();
 sg13g2_fill_2 FILLER_126_183 ();
 sg13g2_decap_8 FILLER_126_190 ();
 sg13g2_decap_8 FILLER_126_197 ();
 sg13g2_fill_2 FILLER_126_204 ();
 sg13g2_fill_1 FILLER_126_206 ();
 sg13g2_decap_8 FILLER_126_221 ();
 sg13g2_decap_4 FILLER_126_228 ();
 sg13g2_fill_2 FILLER_126_232 ();
 sg13g2_decap_8 FILLER_126_237 ();
 sg13g2_decap_8 FILLER_126_261 ();
 sg13g2_fill_1 FILLER_126_268 ();
 sg13g2_decap_8 FILLER_126_279 ();
 sg13g2_decap_4 FILLER_126_286 ();
 sg13g2_fill_1 FILLER_126_290 ();
 sg13g2_decap_8 FILLER_126_295 ();
 sg13g2_decap_8 FILLER_126_302 ();
 sg13g2_fill_2 FILLER_126_309 ();
 sg13g2_fill_1 FILLER_126_311 ();
 sg13g2_fill_2 FILLER_126_343 ();
 sg13g2_fill_1 FILLER_126_345 ();
 sg13g2_decap_8 FILLER_126_382 ();
 sg13g2_decap_4 FILLER_126_389 ();
 sg13g2_decap_4 FILLER_126_415 ();
 sg13g2_fill_1 FILLER_126_429 ();
 sg13g2_decap_8 FILLER_126_443 ();
 sg13g2_decap_8 FILLER_126_457 ();
 sg13g2_decap_4 FILLER_126_464 ();
 sg13g2_fill_1 FILLER_126_468 ();
 sg13g2_decap_8 FILLER_126_486 ();
 sg13g2_decap_8 FILLER_126_493 ();
 sg13g2_decap_8 FILLER_126_500 ();
 sg13g2_decap_4 FILLER_126_507 ();
 sg13g2_fill_1 FILLER_126_511 ();
 sg13g2_decap_8 FILLER_126_516 ();
 sg13g2_decap_8 FILLER_126_523 ();
 sg13g2_decap_8 FILLER_126_530 ();
 sg13g2_fill_1 FILLER_126_537 ();
 sg13g2_decap_8 FILLER_126_602 ();
 sg13g2_decap_8 FILLER_126_609 ();
 sg13g2_decap_4 FILLER_126_616 ();
 sg13g2_fill_2 FILLER_126_620 ();
 sg13g2_decap_4 FILLER_126_673 ();
 sg13g2_fill_2 FILLER_126_677 ();
 sg13g2_fill_2 FILLER_126_714 ();
 sg13g2_fill_1 FILLER_126_716 ();
 sg13g2_decap_8 FILLER_126_725 ();
 sg13g2_fill_2 FILLER_126_732 ();
 sg13g2_decap_8 FILLER_126_790 ();
 sg13g2_decap_8 FILLER_126_797 ();
 sg13g2_decap_4 FILLER_126_804 ();
 sg13g2_fill_2 FILLER_126_808 ();
 sg13g2_decap_8 FILLER_126_815 ();
 sg13g2_fill_2 FILLER_126_822 ();
 sg13g2_fill_1 FILLER_126_824 ();
 sg13g2_decap_8 FILLER_126_829 ();
 sg13g2_decap_8 FILLER_126_836 ();
 sg13g2_decap_8 FILLER_126_843 ();
 sg13g2_decap_8 FILLER_126_863 ();
 sg13g2_decap_8 FILLER_126_870 ();
 sg13g2_decap_8 FILLER_126_877 ();
 sg13g2_fill_2 FILLER_126_884 ();
 sg13g2_fill_1 FILLER_126_890 ();
 sg13g2_fill_1 FILLER_126_904 ();
 sg13g2_decap_8 FILLER_126_934 ();
 sg13g2_decap_8 FILLER_126_941 ();
 sg13g2_decap_4 FILLER_126_948 ();
 sg13g2_decap_4 FILLER_126_978 ();
 sg13g2_fill_1 FILLER_126_982 ();
 sg13g2_fill_1 FILLER_126_988 ();
 sg13g2_decap_8 FILLER_126_1040 ();
 sg13g2_fill_1 FILLER_126_1047 ();
 sg13g2_decap_8 FILLER_126_1052 ();
 sg13g2_decap_8 FILLER_126_1059 ();
 sg13g2_decap_8 FILLER_126_1066 ();
 sg13g2_decap_8 FILLER_126_1073 ();
 sg13g2_decap_8 FILLER_126_1080 ();
 sg13g2_decap_8 FILLER_126_1087 ();
 sg13g2_decap_8 FILLER_126_1094 ();
 sg13g2_decap_8 FILLER_126_1101 ();
 sg13g2_decap_8 FILLER_126_1108 ();
 sg13g2_decap_8 FILLER_126_1115 ();
 sg13g2_decap_8 FILLER_126_1122 ();
 sg13g2_decap_8 FILLER_126_1129 ();
 sg13g2_decap_4 FILLER_126_1136 ();
 sg13g2_fill_2 FILLER_126_1140 ();
 sg13g2_fill_1 FILLER_126_1146 ();
 sg13g2_fill_2 FILLER_126_1152 ();
 sg13g2_fill_1 FILLER_126_1154 ();
 sg13g2_decap_8 FILLER_126_1165 ();
 sg13g2_fill_2 FILLER_126_1172 ();
 sg13g2_fill_1 FILLER_126_1174 ();
 sg13g2_decap_8 FILLER_126_1181 ();
 sg13g2_decap_4 FILLER_126_1188 ();
 sg13g2_fill_1 FILLER_126_1192 ();
 sg13g2_fill_2 FILLER_126_1198 ();
 sg13g2_fill_1 FILLER_126_1200 ();
 sg13g2_decap_4 FILLER_126_1207 ();
 sg13g2_fill_1 FILLER_126_1211 ();
 sg13g2_fill_1 FILLER_126_1225 ();
 sg13g2_fill_1 FILLER_126_1231 ();
 sg13g2_fill_1 FILLER_126_1241 ();
 sg13g2_fill_1 FILLER_126_1247 ();
 sg13g2_fill_1 FILLER_126_1253 ();
 sg13g2_fill_1 FILLER_126_1259 ();
 sg13g2_fill_2 FILLER_126_1265 ();
 sg13g2_fill_2 FILLER_126_1272 ();
 sg13g2_decap_4 FILLER_126_1282 ();
 sg13g2_fill_1 FILLER_126_1286 ();
 sg13g2_decap_8 FILLER_126_1292 ();
 sg13g2_fill_2 FILLER_126_1299 ();
 sg13g2_decap_4 FILLER_126_1306 ();
 sg13g2_decap_8 FILLER_126_1321 ();
 sg13g2_fill_2 FILLER_126_1328 ();
 sg13g2_fill_1 FILLER_126_1330 ();
 sg13g2_fill_1 FILLER_126_1336 ();
 sg13g2_fill_1 FILLER_126_1340 ();
 sg13g2_decap_4 FILLER_126_1347 ();
 sg13g2_decap_8 FILLER_126_1365 ();
 sg13g2_decap_4 FILLER_126_1372 ();
 sg13g2_fill_1 FILLER_126_1376 ();
 sg13g2_decap_8 FILLER_126_1403 ();
 sg13g2_decap_8 FILLER_126_1410 ();
 sg13g2_decap_8 FILLER_126_1417 ();
 sg13g2_decap_8 FILLER_126_1424 ();
 sg13g2_decap_8 FILLER_126_1431 ();
 sg13g2_decap_8 FILLER_126_1438 ();
 sg13g2_decap_8 FILLER_126_1445 ();
 sg13g2_decap_8 FILLER_126_1452 ();
 sg13g2_decap_8 FILLER_126_1459 ();
 sg13g2_decap_8 FILLER_126_1466 ();
 sg13g2_decap_8 FILLER_126_1473 ();
 sg13g2_decap_8 FILLER_126_1480 ();
 sg13g2_decap_8 FILLER_126_1487 ();
 sg13g2_decap_8 FILLER_126_1494 ();
 sg13g2_decap_8 FILLER_126_1501 ();
 sg13g2_decap_8 FILLER_126_1508 ();
 sg13g2_decap_8 FILLER_126_1515 ();
 sg13g2_decap_8 FILLER_126_1522 ();
 sg13g2_decap_8 FILLER_126_1529 ();
 sg13g2_decap_8 FILLER_126_1536 ();
 sg13g2_decap_8 FILLER_126_1543 ();
 sg13g2_decap_8 FILLER_126_1550 ();
 sg13g2_decap_8 FILLER_126_1557 ();
 sg13g2_decap_8 FILLER_126_1564 ();
 sg13g2_decap_8 FILLER_126_1571 ();
 sg13g2_decap_8 FILLER_126_1578 ();
 sg13g2_decap_8 FILLER_126_1585 ();
 sg13g2_decap_8 FILLER_126_1592 ();
 sg13g2_decap_8 FILLER_126_1599 ();
 sg13g2_decap_8 FILLER_126_1606 ();
 sg13g2_decap_8 FILLER_126_1613 ();
 sg13g2_decap_4 FILLER_126_1620 ();
 sg13g2_fill_1 FILLER_126_1624 ();
 sg13g2_decap_8 FILLER_127_0 ();
 sg13g2_fill_1 FILLER_127_11 ();
 sg13g2_fill_2 FILLER_127_16 ();
 sg13g2_fill_1 FILLER_127_28 ();
 sg13g2_decap_4 FILLER_127_43 ();
 sg13g2_fill_2 FILLER_127_47 ();
 sg13g2_decap_8 FILLER_127_61 ();
 sg13g2_fill_2 FILLER_127_68 ();
 sg13g2_fill_1 FILLER_127_70 ();
 sg13g2_decap_8 FILLER_127_76 ();
 sg13g2_decap_4 FILLER_127_83 ();
 sg13g2_fill_1 FILLER_127_87 ();
 sg13g2_fill_1 FILLER_127_93 ();
 sg13g2_decap_4 FILLER_127_99 ();
 sg13g2_fill_2 FILLER_127_103 ();
 sg13g2_fill_2 FILLER_127_131 ();
 sg13g2_decap_4 FILLER_127_138 ();
 sg13g2_decap_8 FILLER_127_146 ();
 sg13g2_decap_4 FILLER_127_153 ();
 sg13g2_fill_1 FILLER_127_157 ();
 sg13g2_decap_8 FILLER_127_184 ();
 sg13g2_decap_8 FILLER_127_191 ();
 sg13g2_decap_8 FILLER_127_198 ();
 sg13g2_decap_8 FILLER_127_205 ();
 sg13g2_decap_8 FILLER_127_212 ();
 sg13g2_decap_8 FILLER_127_219 ();
 sg13g2_fill_2 FILLER_127_226 ();
 sg13g2_fill_1 FILLER_127_228 ();
 sg13g2_fill_1 FILLER_127_259 ();
 sg13g2_fill_2 FILLER_127_270 ();
 sg13g2_decap_8 FILLER_127_284 ();
 sg13g2_decap_8 FILLER_127_291 ();
 sg13g2_decap_8 FILLER_127_298 ();
 sg13g2_fill_2 FILLER_127_305 ();
 sg13g2_decap_8 FILLER_127_311 ();
 sg13g2_decap_8 FILLER_127_322 ();
 sg13g2_decap_4 FILLER_127_329 ();
 sg13g2_fill_1 FILLER_127_333 ();
 sg13g2_decap_8 FILLER_127_355 ();
 sg13g2_fill_1 FILLER_127_362 ();
 sg13g2_fill_1 FILLER_127_368 ();
 sg13g2_fill_2 FILLER_127_373 ();
 sg13g2_fill_1 FILLER_127_375 ();
 sg13g2_fill_2 FILLER_127_383 ();
 sg13g2_decap_4 FILLER_127_390 ();
 sg13g2_fill_1 FILLER_127_394 ();
 sg13g2_decap_8 FILLER_127_407 ();
 sg13g2_fill_2 FILLER_127_414 ();
 sg13g2_fill_1 FILLER_127_416 ();
 sg13g2_fill_1 FILLER_127_423 ();
 sg13g2_fill_2 FILLER_127_429 ();
 sg13g2_fill_1 FILLER_127_431 ();
 sg13g2_decap_8 FILLER_127_437 ();
 sg13g2_decap_4 FILLER_127_452 ();
 sg13g2_decap_8 FILLER_127_459 ();
 sg13g2_decap_8 FILLER_127_466 ();
 sg13g2_fill_2 FILLER_127_486 ();
 sg13g2_decap_8 FILLER_127_494 ();
 sg13g2_decap_4 FILLER_127_501 ();
 sg13g2_decap_8 FILLER_127_513 ();
 sg13g2_decap_8 FILLER_127_520 ();
 sg13g2_decap_8 FILLER_127_527 ();
 sg13g2_fill_2 FILLER_127_534 ();
 sg13g2_decap_4 FILLER_127_540 ();
 sg13g2_fill_1 FILLER_127_544 ();
 sg13g2_decap_8 FILLER_127_550 ();
 sg13g2_fill_1 FILLER_127_557 ();
 sg13g2_fill_2 FILLER_127_616 ();
 sg13g2_fill_1 FILLER_127_618 ();
 sg13g2_fill_2 FILLER_127_645 ();
 sg13g2_decap_8 FILLER_127_718 ();
 sg13g2_decap_8 FILLER_127_725 ();
 sg13g2_decap_4 FILLER_127_732 ();
 sg13g2_fill_2 FILLER_127_736 ();
 sg13g2_fill_2 FILLER_127_742 ();
 sg13g2_fill_1 FILLER_127_744 ();
 sg13g2_decap_8 FILLER_127_749 ();
 sg13g2_decap_8 FILLER_127_756 ();
 sg13g2_decap_8 FILLER_127_763 ();
 sg13g2_fill_2 FILLER_127_770 ();
 sg13g2_decap_8 FILLER_127_776 ();
 sg13g2_decap_4 FILLER_127_783 ();
 sg13g2_decap_8 FILLER_127_791 ();
 sg13g2_decap_4 FILLER_127_802 ();
 sg13g2_fill_2 FILLER_127_815 ();
 sg13g2_decap_8 FILLER_127_843 ();
 sg13g2_decap_4 FILLER_127_850 ();
 sg13g2_decap_8 FILLER_127_858 ();
 sg13g2_decap_8 FILLER_127_865 ();
 sg13g2_decap_8 FILLER_127_872 ();
 sg13g2_fill_1 FILLER_127_879 ();
 sg13g2_decap_4 FILLER_127_898 ();
 sg13g2_decap_4 FILLER_127_910 ();
 sg13g2_fill_1 FILLER_127_914 ();
 sg13g2_decap_8 FILLER_127_931 ();
 sg13g2_decap_4 FILLER_127_938 ();
 sg13g2_fill_2 FILLER_127_942 ();
 sg13g2_decap_8 FILLER_127_948 ();
 sg13g2_decap_8 FILLER_127_955 ();
 sg13g2_decap_8 FILLER_127_962 ();
 sg13g2_decap_4 FILLER_127_969 ();
 sg13g2_fill_2 FILLER_127_976 ();
 sg13g2_fill_1 FILLER_127_978 ();
 sg13g2_fill_1 FILLER_127_988 ();
 sg13g2_fill_1 FILLER_127_1014 ();
 sg13g2_fill_2 FILLER_127_1028 ();
 sg13g2_fill_2 FILLER_127_1084 ();
 sg13g2_fill_1 FILLER_127_1114 ();
 sg13g2_fill_2 FILLER_127_1120 ();
 sg13g2_decap_8 FILLER_127_1126 ();
 sg13g2_fill_2 FILLER_127_1133 ();
 sg13g2_decap_8 FILLER_127_1161 ();
 sg13g2_decap_8 FILLER_127_1168 ();
 sg13g2_fill_2 FILLER_127_1175 ();
 sg13g2_decap_8 FILLER_127_1181 ();
 sg13g2_decap_8 FILLER_127_1188 ();
 sg13g2_decap_8 FILLER_127_1195 ();
 sg13g2_fill_2 FILLER_127_1202 ();
 sg13g2_decap_4 FILLER_127_1210 ();
 sg13g2_fill_1 FILLER_127_1223 ();
 sg13g2_decap_8 FILLER_127_1229 ();
 sg13g2_decap_8 FILLER_127_1236 ();
 sg13g2_fill_2 FILLER_127_1243 ();
 sg13g2_fill_1 FILLER_127_1245 ();
 sg13g2_decap_4 FILLER_127_1251 ();
 sg13g2_fill_2 FILLER_127_1255 ();
 sg13g2_fill_1 FILLER_127_1263 ();
 sg13g2_decap_8 FILLER_127_1268 ();
 sg13g2_decap_4 FILLER_127_1275 ();
 sg13g2_decap_8 FILLER_127_1284 ();
 sg13g2_decap_8 FILLER_127_1291 ();
 sg13g2_decap_8 FILLER_127_1298 ();
 sg13g2_fill_2 FILLER_127_1305 ();
 sg13g2_fill_1 FILLER_127_1311 ();
 sg13g2_fill_1 FILLER_127_1317 ();
 sg13g2_fill_2 FILLER_127_1339 ();
 sg13g2_fill_1 FILLER_127_1341 ();
 sg13g2_fill_2 FILLER_127_1355 ();
 sg13g2_fill_1 FILLER_127_1357 ();
 sg13g2_decap_8 FILLER_127_1362 ();
 sg13g2_fill_2 FILLER_127_1369 ();
 sg13g2_fill_1 FILLER_127_1371 ();
 sg13g2_decap_8 FILLER_127_1404 ();
 sg13g2_decap_8 FILLER_127_1411 ();
 sg13g2_decap_8 FILLER_127_1418 ();
 sg13g2_decap_8 FILLER_127_1425 ();
 sg13g2_decap_8 FILLER_127_1432 ();
 sg13g2_decap_8 FILLER_127_1439 ();
 sg13g2_decap_8 FILLER_127_1446 ();
 sg13g2_decap_8 FILLER_127_1453 ();
 sg13g2_decap_8 FILLER_127_1460 ();
 sg13g2_decap_8 FILLER_127_1467 ();
 sg13g2_decap_8 FILLER_127_1474 ();
 sg13g2_decap_8 FILLER_127_1481 ();
 sg13g2_decap_8 FILLER_127_1488 ();
 sg13g2_decap_8 FILLER_127_1495 ();
 sg13g2_decap_8 FILLER_127_1502 ();
 sg13g2_decap_8 FILLER_127_1509 ();
 sg13g2_decap_8 FILLER_127_1516 ();
 sg13g2_decap_8 FILLER_127_1523 ();
 sg13g2_decap_8 FILLER_127_1530 ();
 sg13g2_decap_8 FILLER_127_1537 ();
 sg13g2_decap_8 FILLER_127_1544 ();
 sg13g2_decap_8 FILLER_127_1551 ();
 sg13g2_decap_8 FILLER_127_1558 ();
 sg13g2_decap_8 FILLER_127_1565 ();
 sg13g2_decap_8 FILLER_127_1572 ();
 sg13g2_decap_8 FILLER_127_1579 ();
 sg13g2_decap_8 FILLER_127_1586 ();
 sg13g2_decap_8 FILLER_127_1593 ();
 sg13g2_decap_8 FILLER_127_1600 ();
 sg13g2_decap_8 FILLER_127_1607 ();
 sg13g2_decap_8 FILLER_127_1614 ();
 sg13g2_decap_4 FILLER_127_1621 ();
 sg13g2_fill_1 FILLER_128_31 ();
 sg13g2_fill_2 FILLER_128_67 ();
 sg13g2_fill_1 FILLER_128_69 ();
 sg13g2_decap_4 FILLER_128_75 ();
 sg13g2_fill_1 FILLER_128_79 ();
 sg13g2_decap_8 FILLER_128_106 ();
 sg13g2_decap_8 FILLER_128_113 ();
 sg13g2_decap_8 FILLER_128_120 ();
 sg13g2_decap_8 FILLER_128_127 ();
 sg13g2_decap_4 FILLER_128_134 ();
 sg13g2_fill_2 FILLER_128_164 ();
 sg13g2_fill_1 FILLER_128_166 ();
 sg13g2_fill_1 FILLER_128_171 ();
 sg13g2_decap_8 FILLER_128_175 ();
 sg13g2_fill_1 FILLER_128_187 ();
 sg13g2_decap_4 FILLER_128_198 ();
 sg13g2_fill_1 FILLER_128_202 ();
 sg13g2_decap_8 FILLER_128_214 ();
 sg13g2_decap_4 FILLER_128_221 ();
 sg13g2_fill_2 FILLER_128_225 ();
 sg13g2_fill_1 FILLER_128_253 ();
 sg13g2_fill_2 FILLER_128_286 ();
 sg13g2_fill_1 FILLER_128_288 ();
 sg13g2_fill_2 FILLER_128_293 ();
 sg13g2_fill_1 FILLER_128_298 ();
 sg13g2_fill_1 FILLER_128_325 ();
 sg13g2_fill_1 FILLER_128_334 ();
 sg13g2_decap_8 FILLER_128_340 ();
 sg13g2_fill_2 FILLER_128_347 ();
 sg13g2_fill_1 FILLER_128_349 ();
 sg13g2_fill_1 FILLER_128_357 ();
 sg13g2_fill_2 FILLER_128_381 ();
 sg13g2_fill_1 FILLER_128_390 ();
 sg13g2_decap_8 FILLER_128_403 ();
 sg13g2_decap_8 FILLER_128_410 ();
 sg13g2_fill_2 FILLER_128_417 ();
 sg13g2_decap_8 FILLER_128_446 ();
 sg13g2_decap_8 FILLER_128_453 ();
 sg13g2_fill_2 FILLER_128_465 ();
 sg13g2_fill_2 FILLER_128_480 ();
 sg13g2_fill_1 FILLER_128_497 ();
 sg13g2_fill_1 FILLER_128_509 ();
 sg13g2_decap_4 FILLER_128_517 ();
 sg13g2_fill_1 FILLER_128_521 ();
 sg13g2_fill_2 FILLER_128_597 ();
 sg13g2_decap_4 FILLER_128_633 ();
 sg13g2_decap_4 FILLER_128_641 ();
 sg13g2_fill_1 FILLER_128_645 ();
 sg13g2_decap_8 FILLER_128_675 ();
 sg13g2_decap_4 FILLER_128_682 ();
 sg13g2_fill_1 FILLER_128_686 ();
 sg13g2_decap_8 FILLER_128_691 ();
 sg13g2_fill_2 FILLER_128_698 ();
 sg13g2_fill_1 FILLER_128_700 ();
 sg13g2_decap_4 FILLER_128_709 ();
 sg13g2_fill_2 FILLER_128_713 ();
 sg13g2_decap_8 FILLER_128_719 ();
 sg13g2_decap_4 FILLER_128_726 ();
 sg13g2_fill_1 FILLER_128_730 ();
 sg13g2_fill_2 FILLER_128_757 ();
 sg13g2_fill_1 FILLER_128_759 ();
 sg13g2_decap_8 FILLER_128_799 ();
 sg13g2_decap_4 FILLER_128_806 ();
 sg13g2_fill_1 FILLER_128_810 ();
 sg13g2_decap_8 FILLER_128_816 ();
 sg13g2_decap_8 FILLER_128_872 ();
 sg13g2_decap_8 FILLER_128_887 ();
 sg13g2_decap_8 FILLER_128_894 ();
 sg13g2_decap_8 FILLER_128_901 ();
 sg13g2_fill_1 FILLER_128_908 ();
 sg13g2_decap_4 FILLER_128_913 ();
 sg13g2_decap_8 FILLER_128_922 ();
 sg13g2_decap_8 FILLER_128_929 ();
 sg13g2_fill_1 FILLER_128_936 ();
 sg13g2_decap_4 FILLER_128_1078 ();
 sg13g2_fill_1 FILLER_128_1082 ();
 sg13g2_fill_1 FILLER_128_1140 ();
 sg13g2_decap_4 FILLER_128_1145 ();
 sg13g2_fill_1 FILLER_128_1149 ();
 sg13g2_fill_2 FILLER_128_1159 ();
 sg13g2_decap_4 FILLER_128_1171 ();
 sg13g2_decap_8 FILLER_128_1193 ();
 sg13g2_decap_8 FILLER_128_1204 ();
 sg13g2_decap_4 FILLER_128_1211 ();
 sg13g2_fill_2 FILLER_128_1215 ();
 sg13g2_decap_8 FILLER_128_1229 ();
 sg13g2_decap_8 FILLER_128_1236 ();
 sg13g2_decap_8 FILLER_128_1243 ();
 sg13g2_decap_8 FILLER_128_1250 ();
 sg13g2_decap_8 FILLER_128_1257 ();
 sg13g2_decap_8 FILLER_128_1264 ();
 sg13g2_decap_8 FILLER_128_1271 ();
 sg13g2_decap_8 FILLER_128_1278 ();
 sg13g2_decap_8 FILLER_128_1285 ();
 sg13g2_fill_2 FILLER_128_1297 ();
 sg13g2_decap_4 FILLER_128_1326 ();
 sg13g2_fill_1 FILLER_128_1330 ();
 sg13g2_fill_2 FILLER_128_1349 ();
 sg13g2_decap_8 FILLER_128_1360 ();
 sg13g2_decap_4 FILLER_128_1367 ();
 sg13g2_fill_1 FILLER_128_1371 ();
 sg13g2_decap_8 FILLER_128_1398 ();
 sg13g2_decap_8 FILLER_128_1405 ();
 sg13g2_decap_8 FILLER_128_1412 ();
 sg13g2_decap_8 FILLER_128_1419 ();
 sg13g2_decap_8 FILLER_128_1426 ();
 sg13g2_decap_8 FILLER_128_1433 ();
 sg13g2_decap_8 FILLER_128_1440 ();
 sg13g2_decap_8 FILLER_128_1447 ();
 sg13g2_decap_8 FILLER_128_1454 ();
 sg13g2_decap_8 FILLER_128_1461 ();
 sg13g2_decap_8 FILLER_128_1468 ();
 sg13g2_decap_8 FILLER_128_1475 ();
 sg13g2_decap_8 FILLER_128_1482 ();
 sg13g2_decap_8 FILLER_128_1489 ();
 sg13g2_decap_8 FILLER_128_1496 ();
 sg13g2_decap_8 FILLER_128_1503 ();
 sg13g2_decap_8 FILLER_128_1510 ();
 sg13g2_decap_8 FILLER_128_1517 ();
 sg13g2_decap_8 FILLER_128_1524 ();
 sg13g2_decap_8 FILLER_128_1531 ();
 sg13g2_decap_8 FILLER_128_1538 ();
 sg13g2_decap_8 FILLER_128_1545 ();
 sg13g2_decap_8 FILLER_128_1552 ();
 sg13g2_decap_8 FILLER_128_1559 ();
 sg13g2_decap_8 FILLER_128_1566 ();
 sg13g2_decap_8 FILLER_128_1573 ();
 sg13g2_decap_8 FILLER_128_1580 ();
 sg13g2_decap_8 FILLER_128_1587 ();
 sg13g2_decap_8 FILLER_128_1594 ();
 sg13g2_decap_8 FILLER_128_1601 ();
 sg13g2_decap_8 FILLER_128_1608 ();
 sg13g2_decap_8 FILLER_128_1615 ();
 sg13g2_fill_2 FILLER_128_1622 ();
 sg13g2_fill_1 FILLER_128_1624 ();
 sg13g2_decap_8 FILLER_129_0 ();
 sg13g2_decap_8 FILLER_129_7 ();
 sg13g2_decap_8 FILLER_129_14 ();
 sg13g2_decap_8 FILLER_129_21 ();
 sg13g2_decap_8 FILLER_129_28 ();
 sg13g2_decap_4 FILLER_129_35 ();
 sg13g2_fill_1 FILLER_129_39 ();
 sg13g2_fill_2 FILLER_129_56 ();
 sg13g2_fill_2 FILLER_129_68 ();
 sg13g2_fill_1 FILLER_129_70 ();
 sg13g2_fill_2 FILLER_129_76 ();
 sg13g2_fill_1 FILLER_129_78 ();
 sg13g2_decap_4 FILLER_129_83 ();
 sg13g2_fill_1 FILLER_129_87 ();
 sg13g2_decap_8 FILLER_129_92 ();
 sg13g2_decap_8 FILLER_129_99 ();
 sg13g2_decap_8 FILLER_129_106 ();
 sg13g2_decap_8 FILLER_129_113 ();
 sg13g2_decap_8 FILLER_129_120 ();
 sg13g2_decap_8 FILLER_129_127 ();
 sg13g2_decap_8 FILLER_129_134 ();
 sg13g2_fill_2 FILLER_129_141 ();
 sg13g2_fill_2 FILLER_129_201 ();
 sg13g2_fill_2 FILLER_129_234 ();
 sg13g2_fill_1 FILLER_129_245 ();
 sg13g2_decap_8 FILLER_129_338 ();
 sg13g2_decap_8 FILLER_129_345 ();
 sg13g2_fill_1 FILLER_129_352 ();
 sg13g2_decap_8 FILLER_129_397 ();
 sg13g2_decap_4 FILLER_129_404 ();
 sg13g2_fill_1 FILLER_129_408 ();
 sg13g2_decap_8 FILLER_129_414 ();
 sg13g2_fill_1 FILLER_129_425 ();
 sg13g2_fill_1 FILLER_129_430 ();
 sg13g2_decap_8 FILLER_129_437 ();
 sg13g2_decap_4 FILLER_129_444 ();
 sg13g2_fill_2 FILLER_129_457 ();
 sg13g2_fill_1 FILLER_129_459 ();
 sg13g2_decap_8 FILLER_129_466 ();
 sg13g2_fill_2 FILLER_129_473 ();
 sg13g2_fill_1 FILLER_129_475 ();
 sg13g2_fill_2 FILLER_129_481 ();
 sg13g2_decap_4 FILLER_129_488 ();
 sg13g2_fill_2 FILLER_129_492 ();
 sg13g2_decap_8 FILLER_129_499 ();
 sg13g2_fill_2 FILLER_129_506 ();
 sg13g2_fill_1 FILLER_129_508 ();
 sg13g2_decap_4 FILLER_129_513 ();
 sg13g2_decap_8 FILLER_129_522 ();
 sg13g2_fill_2 FILLER_129_529 ();
 sg13g2_fill_1 FILLER_129_531 ();
 sg13g2_decap_8 FILLER_129_541 ();
 sg13g2_decap_4 FILLER_129_548 ();
 sg13g2_fill_1 FILLER_129_552 ();
 sg13g2_decap_8 FILLER_129_596 ();
 sg13g2_fill_1 FILLER_129_603 ();
 sg13g2_fill_2 FILLER_129_655 ();
 sg13g2_decap_8 FILLER_129_661 ();
 sg13g2_decap_8 FILLER_129_696 ();
 sg13g2_decap_4 FILLER_129_703 ();
 sg13g2_fill_1 FILLER_129_707 ();
 sg13g2_decap_8 FILLER_129_734 ();
 sg13g2_fill_1 FILLER_129_741 ();
 sg13g2_decap_4 FILLER_129_755 ();
 sg13g2_decap_8 FILLER_129_773 ();
 sg13g2_decap_4 FILLER_129_780 ();
 sg13g2_fill_2 FILLER_129_810 ();
 sg13g2_fill_1 FILLER_129_812 ();
 sg13g2_decap_4 FILLER_129_821 ();
 sg13g2_fill_2 FILLER_129_825 ();
 sg13g2_decap_8 FILLER_129_835 ();
 sg13g2_decap_4 FILLER_129_842 ();
 sg13g2_fill_2 FILLER_129_846 ();
 sg13g2_decap_8 FILLER_129_853 ();
 sg13g2_fill_1 FILLER_129_860 ();
 sg13g2_fill_2 FILLER_129_875 ();
 sg13g2_fill_1 FILLER_129_877 ();
 sg13g2_decap_8 FILLER_129_883 ();
 sg13g2_fill_2 FILLER_129_894 ();
 sg13g2_decap_8 FILLER_129_927 ();
 sg13g2_fill_2 FILLER_129_934 ();
 sg13g2_decap_8 FILLER_129_944 ();
 sg13g2_decap_4 FILLER_129_951 ();
 sg13g2_fill_1 FILLER_129_955 ();
 sg13g2_fill_2 FILLER_129_966 ();
 sg13g2_fill_1 FILLER_129_968 ();
 sg13g2_decap_8 FILLER_129_1074 ();
 sg13g2_decap_4 FILLER_129_1081 ();
 sg13g2_fill_2 FILLER_129_1089 ();
 sg13g2_fill_2 FILLER_129_1120 ();
 sg13g2_fill_1 FILLER_129_1122 ();
 sg13g2_fill_2 FILLER_129_1151 ();
 sg13g2_fill_1 FILLER_129_1166 ();
 sg13g2_decap_4 FILLER_129_1180 ();
 sg13g2_fill_1 FILLER_129_1184 ();
 sg13g2_decap_8 FILLER_129_1202 ();
 sg13g2_decap_4 FILLER_129_1209 ();
 sg13g2_fill_1 FILLER_129_1225 ();
 sg13g2_decap_8 FILLER_129_1242 ();
 sg13g2_decap_4 FILLER_129_1249 ();
 sg13g2_fill_2 FILLER_129_1278 ();
 sg13g2_decap_4 FILLER_129_1284 ();
 sg13g2_decap_8 FILLER_129_1298 ();
 sg13g2_decap_8 FILLER_129_1305 ();
 sg13g2_decap_8 FILLER_129_1321 ();
 sg13g2_decap_8 FILLER_129_1328 ();
 sg13g2_decap_8 FILLER_129_1335 ();
 sg13g2_fill_2 FILLER_129_1342 ();
 sg13g2_fill_1 FILLER_129_1344 ();
 sg13g2_fill_2 FILLER_129_1349 ();
 sg13g2_fill_1 FILLER_129_1351 ();
 sg13g2_decap_8 FILLER_129_1371 ();
 sg13g2_decap_8 FILLER_129_1378 ();
 sg13g2_decap_8 FILLER_129_1385 ();
 sg13g2_decap_8 FILLER_129_1392 ();
 sg13g2_decap_8 FILLER_129_1399 ();
 sg13g2_decap_8 FILLER_129_1406 ();
 sg13g2_decap_8 FILLER_129_1413 ();
 sg13g2_decap_8 FILLER_129_1420 ();
 sg13g2_decap_8 FILLER_129_1427 ();
 sg13g2_decap_8 FILLER_129_1434 ();
 sg13g2_decap_8 FILLER_129_1441 ();
 sg13g2_decap_8 FILLER_129_1448 ();
 sg13g2_decap_8 FILLER_129_1455 ();
 sg13g2_decap_8 FILLER_129_1462 ();
 sg13g2_decap_8 FILLER_129_1469 ();
 sg13g2_decap_8 FILLER_129_1476 ();
 sg13g2_decap_8 FILLER_129_1483 ();
 sg13g2_decap_8 FILLER_129_1490 ();
 sg13g2_decap_8 FILLER_129_1497 ();
 sg13g2_decap_8 FILLER_129_1504 ();
 sg13g2_decap_8 FILLER_129_1511 ();
 sg13g2_decap_8 FILLER_129_1518 ();
 sg13g2_decap_8 FILLER_129_1525 ();
 sg13g2_decap_8 FILLER_129_1532 ();
 sg13g2_decap_8 FILLER_129_1539 ();
 sg13g2_decap_8 FILLER_129_1546 ();
 sg13g2_decap_8 FILLER_129_1553 ();
 sg13g2_decap_8 FILLER_129_1560 ();
 sg13g2_decap_8 FILLER_129_1567 ();
 sg13g2_decap_8 FILLER_129_1574 ();
 sg13g2_decap_8 FILLER_129_1581 ();
 sg13g2_decap_8 FILLER_129_1588 ();
 sg13g2_decap_8 FILLER_129_1595 ();
 sg13g2_decap_8 FILLER_129_1602 ();
 sg13g2_decap_8 FILLER_129_1609 ();
 sg13g2_decap_8 FILLER_129_1616 ();
 sg13g2_fill_2 FILLER_129_1623 ();
 sg13g2_fill_2 FILLER_130_0 ();
 sg13g2_decap_4 FILLER_130_30 ();
 sg13g2_fill_1 FILLER_130_34 ();
 sg13g2_fill_2 FILLER_130_72 ();
 sg13g2_decap_8 FILLER_130_104 ();
 sg13g2_decap_8 FILLER_130_111 ();
 sg13g2_decap_8 FILLER_130_118 ();
 sg13g2_fill_2 FILLER_130_125 ();
 sg13g2_fill_1 FILLER_130_127 ();
 sg13g2_decap_8 FILLER_130_132 ();
 sg13g2_fill_1 FILLER_130_175 ();
 sg13g2_decap_8 FILLER_130_207 ();
 sg13g2_fill_2 FILLER_130_214 ();
 sg13g2_fill_2 FILLER_130_245 ();
 sg13g2_decap_4 FILLER_130_287 ();
 sg13g2_fill_1 FILLER_130_300 ();
 sg13g2_fill_2 FILLER_130_360 ();
 sg13g2_fill_1 FILLER_130_362 ();
 sg13g2_decap_4 FILLER_130_388 ();
 sg13g2_decap_4 FILLER_130_396 ();
 sg13g2_fill_2 FILLER_130_400 ();
 sg13g2_fill_1 FILLER_130_426 ();
 sg13g2_fill_2 FILLER_130_437 ();
 sg13g2_fill_2 FILLER_130_470 ();
 sg13g2_fill_1 FILLER_130_472 ();
 sg13g2_fill_1 FILLER_130_492 ();
 sg13g2_fill_2 FILLER_130_502 ();
 sg13g2_fill_1 FILLER_130_504 ();
 sg13g2_decap_8 FILLER_130_510 ();
 sg13g2_fill_2 FILLER_130_517 ();
 sg13g2_decap_8 FILLER_130_523 ();
 sg13g2_decap_8 FILLER_130_530 ();
 sg13g2_decap_8 FILLER_130_537 ();
 sg13g2_decap_8 FILLER_130_544 ();
 sg13g2_decap_4 FILLER_130_551 ();
 sg13g2_fill_1 FILLER_130_555 ();
 sg13g2_decap_4 FILLER_130_587 ();
 sg13g2_decap_8 FILLER_130_595 ();
 sg13g2_decap_8 FILLER_130_602 ();
 sg13g2_decap_4 FILLER_130_609 ();
 sg13g2_fill_2 FILLER_130_622 ();
 sg13g2_fill_1 FILLER_130_624 ();
 sg13g2_fill_2 FILLER_130_676 ();
 sg13g2_fill_1 FILLER_130_678 ();
 sg13g2_decap_4 FILLER_130_711 ();
 sg13g2_decap_8 FILLER_130_844 ();
 sg13g2_decap_8 FILLER_130_851 ();
 sg13g2_decap_4 FILLER_130_858 ();
 sg13g2_fill_2 FILLER_130_862 ();
 sg13g2_decap_8 FILLER_130_870 ();
 sg13g2_fill_2 FILLER_130_877 ();
 sg13g2_fill_1 FILLER_130_879 ();
 sg13g2_decap_8 FILLER_130_885 ();
 sg13g2_decap_8 FILLER_130_892 ();
 sg13g2_decap_8 FILLER_130_899 ();
 sg13g2_decap_4 FILLER_130_906 ();
 sg13g2_decap_4 FILLER_130_914 ();
 sg13g2_decap_8 FILLER_130_922 ();
 sg13g2_fill_1 FILLER_130_960 ();
 sg13g2_fill_1 FILLER_130_994 ();
 sg13g2_decap_4 FILLER_130_1034 ();
 sg13g2_fill_2 FILLER_130_1077 ();
 sg13g2_decap_8 FILLER_130_1087 ();
 sg13g2_fill_1 FILLER_130_1094 ();
 sg13g2_decap_4 FILLER_130_1104 ();
 sg13g2_fill_1 FILLER_130_1119 ();
 sg13g2_decap_4 FILLER_130_1171 ();
 sg13g2_fill_1 FILLER_130_1189 ();
 sg13g2_fill_1 FILLER_130_1204 ();
 sg13g2_decap_8 FILLER_130_1209 ();
 sg13g2_decap_8 FILLER_130_1216 ();
 sg13g2_decap_4 FILLER_130_1223 ();
 sg13g2_fill_1 FILLER_130_1227 ();
 sg13g2_fill_2 FILLER_130_1259 ();
 sg13g2_fill_1 FILLER_130_1261 ();
 sg13g2_fill_2 FILLER_130_1275 ();
 sg13g2_decap_8 FILLER_130_1287 ();
 sg13g2_decap_8 FILLER_130_1294 ();
 sg13g2_decap_8 FILLER_130_1301 ();
 sg13g2_decap_4 FILLER_130_1308 ();
 sg13g2_fill_1 FILLER_130_1317 ();
 sg13g2_decap_8 FILLER_130_1326 ();
 sg13g2_decap_8 FILLER_130_1333 ();
 sg13g2_decap_8 FILLER_130_1340 ();
 sg13g2_fill_1 FILLER_130_1347 ();
 sg13g2_decap_8 FILLER_130_1357 ();
 sg13g2_fill_2 FILLER_130_1364 ();
 sg13g2_fill_1 FILLER_130_1366 ();
 sg13g2_decap_8 FILLER_130_1372 ();
 sg13g2_fill_2 FILLER_130_1379 ();
 sg13g2_decap_8 FILLER_130_1385 ();
 sg13g2_decap_8 FILLER_130_1392 ();
 sg13g2_decap_8 FILLER_130_1399 ();
 sg13g2_decap_8 FILLER_130_1406 ();
 sg13g2_decap_8 FILLER_130_1413 ();
 sg13g2_decap_8 FILLER_130_1420 ();
 sg13g2_decap_8 FILLER_130_1427 ();
 sg13g2_decap_8 FILLER_130_1434 ();
 sg13g2_decap_8 FILLER_130_1441 ();
 sg13g2_decap_8 FILLER_130_1448 ();
 sg13g2_decap_8 FILLER_130_1455 ();
 sg13g2_decap_8 FILLER_130_1462 ();
 sg13g2_decap_8 FILLER_130_1469 ();
 sg13g2_decap_8 FILLER_130_1476 ();
 sg13g2_decap_8 FILLER_130_1483 ();
 sg13g2_decap_8 FILLER_130_1490 ();
 sg13g2_decap_8 FILLER_130_1497 ();
 sg13g2_decap_8 FILLER_130_1504 ();
 sg13g2_decap_8 FILLER_130_1511 ();
 sg13g2_decap_8 FILLER_130_1518 ();
 sg13g2_decap_8 FILLER_130_1525 ();
 sg13g2_decap_8 FILLER_130_1532 ();
 sg13g2_decap_8 FILLER_130_1539 ();
 sg13g2_decap_8 FILLER_130_1546 ();
 sg13g2_decap_8 FILLER_130_1553 ();
 sg13g2_decap_8 FILLER_130_1560 ();
 sg13g2_decap_8 FILLER_130_1567 ();
 sg13g2_decap_8 FILLER_130_1574 ();
 sg13g2_decap_8 FILLER_130_1581 ();
 sg13g2_decap_8 FILLER_130_1588 ();
 sg13g2_decap_8 FILLER_130_1595 ();
 sg13g2_decap_8 FILLER_130_1602 ();
 sg13g2_decap_8 FILLER_130_1609 ();
 sg13g2_decap_8 FILLER_130_1616 ();
 sg13g2_fill_2 FILLER_130_1623 ();
 sg13g2_fill_2 FILLER_131_31 ();
 sg13g2_fill_1 FILLER_131_33 ();
 sg13g2_decap_8 FILLER_131_94 ();
 sg13g2_fill_2 FILLER_131_101 ();
 sg13g2_fill_2 FILLER_131_107 ();
 sg13g2_fill_1 FILLER_131_109 ();
 sg13g2_decap_4 FILLER_131_114 ();
 sg13g2_fill_1 FILLER_131_118 ();
 sg13g2_fill_1 FILLER_131_123 ();
 sg13g2_fill_2 FILLER_131_178 ();
 sg13g2_fill_2 FILLER_131_185 ();
 sg13g2_decap_8 FILLER_131_191 ();
 sg13g2_fill_1 FILLER_131_198 ();
 sg13g2_fill_2 FILLER_131_209 ();
 sg13g2_fill_1 FILLER_131_211 ();
 sg13g2_fill_2 FILLER_131_243 ();
 sg13g2_fill_1 FILLER_131_278 ();
 sg13g2_decap_4 FILLER_131_412 ();
 sg13g2_fill_1 FILLER_131_416 ();
 sg13g2_decap_8 FILLER_131_422 ();
 sg13g2_decap_8 FILLER_131_429 ();
 sg13g2_fill_2 FILLER_131_436 ();
 sg13g2_fill_1 FILLER_131_438 ();
 sg13g2_decap_8 FILLER_131_450 ();
 sg13g2_decap_8 FILLER_131_457 ();
 sg13g2_decap_8 FILLER_131_464 ();
 sg13g2_decap_8 FILLER_131_471 ();
 sg13g2_fill_2 FILLER_131_478 ();
 sg13g2_decap_4 FILLER_131_484 ();
 sg13g2_decap_4 FILLER_131_499 ();
 sg13g2_fill_1 FILLER_131_544 ();
 sg13g2_decap_4 FILLER_131_551 ();
 sg13g2_fill_2 FILLER_131_560 ();
 sg13g2_fill_2 FILLER_131_568 ();
 sg13g2_decap_8 FILLER_131_574 ();
 sg13g2_fill_2 FILLER_131_581 ();
 sg13g2_fill_1 FILLER_131_583 ();
 sg13g2_decap_8 FILLER_131_678 ();
 sg13g2_decap_8 FILLER_131_685 ();
 sg13g2_decap_8 FILLER_131_692 ();
 sg13g2_decap_8 FILLER_131_699 ();
 sg13g2_fill_2 FILLER_131_706 ();
 sg13g2_fill_1 FILLER_131_708 ();
 sg13g2_fill_2 FILLER_131_735 ();
 sg13g2_fill_2 FILLER_131_747 ();
 sg13g2_fill_1 FILLER_131_754 ();
 sg13g2_fill_2 FILLER_131_781 ();
 sg13g2_fill_1 FILLER_131_783 ();
 sg13g2_fill_1 FILLER_131_813 ();
 sg13g2_decap_8 FILLER_131_818 ();
 sg13g2_decap_4 FILLER_131_829 ();
 sg13g2_fill_1 FILLER_131_833 ();
 sg13g2_fill_1 FILLER_131_844 ();
 sg13g2_decap_4 FILLER_131_871 ();
 sg13g2_decap_8 FILLER_131_907 ();
 sg13g2_decap_8 FILLER_131_914 ();
 sg13g2_fill_1 FILLER_131_921 ();
 sg13g2_fill_1 FILLER_131_964 ();
 sg13g2_fill_2 FILLER_131_1001 ();
 sg13g2_decap_8 FILLER_131_1022 ();
 sg13g2_decap_8 FILLER_131_1029 ();
 sg13g2_decap_8 FILLER_131_1036 ();
 sg13g2_decap_8 FILLER_131_1043 ();
 sg13g2_decap_8 FILLER_131_1050 ();
 sg13g2_decap_8 FILLER_131_1057 ();
 sg13g2_decap_8 FILLER_131_1064 ();
 sg13g2_fill_1 FILLER_131_1071 ();
 sg13g2_decap_8 FILLER_131_1076 ();
 sg13g2_decap_8 FILLER_131_1083 ();
 sg13g2_fill_2 FILLER_131_1116 ();
 sg13g2_fill_2 FILLER_131_1148 ();
 sg13g2_decap_4 FILLER_131_1154 ();
 sg13g2_decap_4 FILLER_131_1191 ();
 sg13g2_fill_2 FILLER_131_1195 ();
 sg13g2_fill_1 FILLER_131_1223 ();
 sg13g2_fill_1 FILLER_131_1242 ();
 sg13g2_fill_2 FILLER_131_1247 ();
 sg13g2_fill_1 FILLER_131_1249 ();
 sg13g2_fill_1 FILLER_131_1258 ();
 sg13g2_decap_8 FILLER_131_1270 ();
 sg13g2_fill_2 FILLER_131_1277 ();
 sg13g2_fill_1 FILLER_131_1279 ();
 sg13g2_fill_1 FILLER_131_1284 ();
 sg13g2_fill_2 FILLER_131_1290 ();
 sg13g2_decap_8 FILLER_131_1297 ();
 sg13g2_decap_8 FILLER_131_1304 ();
 sg13g2_fill_2 FILLER_131_1311 ();
 sg13g2_fill_1 FILLER_131_1313 ();
 sg13g2_fill_1 FILLER_131_1319 ();
 sg13g2_fill_2 FILLER_131_1326 ();
 sg13g2_fill_2 FILLER_131_1337 ();
 sg13g2_fill_1 FILLER_131_1339 ();
 sg13g2_fill_2 FILLER_131_1344 ();
 sg13g2_fill_1 FILLER_131_1346 ();
 sg13g2_decap_8 FILLER_131_1355 ();
 sg13g2_decap_8 FILLER_131_1362 ();
 sg13g2_fill_2 FILLER_131_1369 ();
 sg13g2_fill_1 FILLER_131_1371 ();
 sg13g2_decap_8 FILLER_131_1398 ();
 sg13g2_decap_8 FILLER_131_1405 ();
 sg13g2_decap_8 FILLER_131_1412 ();
 sg13g2_decap_8 FILLER_131_1419 ();
 sg13g2_decap_8 FILLER_131_1426 ();
 sg13g2_decap_8 FILLER_131_1433 ();
 sg13g2_decap_8 FILLER_131_1440 ();
 sg13g2_decap_8 FILLER_131_1447 ();
 sg13g2_decap_8 FILLER_131_1454 ();
 sg13g2_decap_8 FILLER_131_1461 ();
 sg13g2_decap_8 FILLER_131_1468 ();
 sg13g2_decap_8 FILLER_131_1475 ();
 sg13g2_decap_8 FILLER_131_1482 ();
 sg13g2_decap_8 FILLER_131_1489 ();
 sg13g2_decap_8 FILLER_131_1496 ();
 sg13g2_decap_8 FILLER_131_1503 ();
 sg13g2_decap_8 FILLER_131_1510 ();
 sg13g2_decap_8 FILLER_131_1517 ();
 sg13g2_decap_8 FILLER_131_1524 ();
 sg13g2_decap_8 FILLER_131_1531 ();
 sg13g2_decap_8 FILLER_131_1538 ();
 sg13g2_decap_8 FILLER_131_1545 ();
 sg13g2_decap_8 FILLER_131_1552 ();
 sg13g2_decap_8 FILLER_131_1559 ();
 sg13g2_decap_8 FILLER_131_1566 ();
 sg13g2_decap_8 FILLER_131_1573 ();
 sg13g2_decap_8 FILLER_131_1580 ();
 sg13g2_decap_8 FILLER_131_1587 ();
 sg13g2_decap_8 FILLER_131_1594 ();
 sg13g2_decap_8 FILLER_131_1601 ();
 sg13g2_decap_8 FILLER_131_1608 ();
 sg13g2_decap_8 FILLER_131_1615 ();
 sg13g2_fill_2 FILLER_131_1622 ();
 sg13g2_fill_1 FILLER_131_1624 ();
 sg13g2_decap_8 FILLER_132_0 ();
 sg13g2_decap_4 FILLER_132_11 ();
 sg13g2_fill_2 FILLER_132_19 ();
 sg13g2_fill_1 FILLER_132_21 ();
 sg13g2_decap_8 FILLER_132_32 ();
 sg13g2_decap_8 FILLER_132_39 ();
 sg13g2_fill_1 FILLER_132_46 ();
 sg13g2_fill_2 FILLER_132_51 ();
 sg13g2_fill_2 FILLER_132_61 ();
 sg13g2_decap_4 FILLER_132_92 ();
 sg13g2_decap_8 FILLER_132_148 ();
 sg13g2_fill_2 FILLER_132_155 ();
 sg13g2_fill_1 FILLER_132_157 ();
 sg13g2_decap_8 FILLER_132_172 ();
 sg13g2_decap_4 FILLER_132_198 ();
 sg13g2_decap_8 FILLER_132_213 ();
 sg13g2_decap_8 FILLER_132_223 ();
 sg13g2_decap_4 FILLER_132_230 ();
 sg13g2_fill_1 FILLER_132_234 ();
 sg13g2_decap_8 FILLER_132_244 ();
 sg13g2_decap_8 FILLER_132_251 ();
 sg13g2_fill_1 FILLER_132_258 ();
 sg13g2_decap_8 FILLER_132_263 ();
 sg13g2_decap_8 FILLER_132_270 ();
 sg13g2_decap_8 FILLER_132_277 ();
 sg13g2_decap_4 FILLER_132_284 ();
 sg13g2_fill_2 FILLER_132_293 ();
 sg13g2_fill_2 FILLER_132_321 ();
 sg13g2_fill_2 FILLER_132_332 ();
 sg13g2_decap_8 FILLER_132_339 ();
 sg13g2_fill_2 FILLER_132_346 ();
 sg13g2_fill_1 FILLER_132_348 ();
 sg13g2_decap_8 FILLER_132_381 ();
 sg13g2_decap_4 FILLER_132_388 ();
 sg13g2_decap_8 FILLER_132_397 ();
 sg13g2_fill_2 FILLER_132_404 ();
 sg13g2_fill_1 FILLER_132_406 ();
 sg13g2_decap_8 FILLER_132_412 ();
 sg13g2_decap_8 FILLER_132_419 ();
 sg13g2_decap_8 FILLER_132_426 ();
 sg13g2_fill_2 FILLER_132_455 ();
 sg13g2_fill_1 FILLER_132_457 ();
 sg13g2_fill_2 FILLER_132_465 ();
 sg13g2_decap_8 FILLER_132_472 ();
 sg13g2_fill_2 FILLER_132_479 ();
 sg13g2_fill_1 FILLER_132_481 ();
 sg13g2_decap_8 FILLER_132_497 ();
 sg13g2_decap_4 FILLER_132_504 ();
 sg13g2_fill_1 FILLER_132_508 ();
 sg13g2_decap_8 FILLER_132_513 ();
 sg13g2_decap_8 FILLER_132_520 ();
 sg13g2_decap_8 FILLER_132_527 ();
 sg13g2_fill_2 FILLER_132_534 ();
 sg13g2_fill_1 FILLER_132_536 ();
 sg13g2_decap_8 FILLER_132_543 ();
 sg13g2_fill_1 FILLER_132_550 ();
 sg13g2_fill_2 FILLER_132_556 ();
 sg13g2_decap_8 FILLER_132_565 ();
 sg13g2_decap_8 FILLER_132_572 ();
 sg13g2_decap_8 FILLER_132_579 ();
 sg13g2_decap_8 FILLER_132_586 ();
 sg13g2_decap_8 FILLER_132_593 ();
 sg13g2_fill_2 FILLER_132_612 ();
 sg13g2_fill_2 FILLER_132_649 ();
 sg13g2_decap_8 FILLER_132_677 ();
 sg13g2_decap_8 FILLER_132_684 ();
 sg13g2_decap_8 FILLER_132_691 ();
 sg13g2_decap_8 FILLER_132_698 ();
 sg13g2_fill_1 FILLER_132_705 ();
 sg13g2_decap_8 FILLER_132_766 ();
 sg13g2_decap_8 FILLER_132_842 ();
 sg13g2_decap_4 FILLER_132_849 ();
 sg13g2_fill_2 FILLER_132_857 ();
 sg13g2_fill_1 FILLER_132_859 ();
 sg13g2_fill_1 FILLER_132_890 ();
 sg13g2_decap_8 FILLER_132_900 ();
 sg13g2_decap_8 FILLER_132_907 ();
 sg13g2_decap_8 FILLER_132_914 ();
 sg13g2_decap_4 FILLER_132_925 ();
 sg13g2_fill_1 FILLER_132_929 ();
 sg13g2_decap_8 FILLER_132_942 ();
 sg13g2_fill_2 FILLER_132_989 ();
 sg13g2_decap_8 FILLER_132_1025 ();
 sg13g2_decap_8 FILLER_132_1032 ();
 sg13g2_decap_4 FILLER_132_1039 ();
 sg13g2_fill_1 FILLER_132_1043 ();
 sg13g2_fill_1 FILLER_132_1048 ();
 sg13g2_decap_8 FILLER_132_1055 ();
 sg13g2_fill_2 FILLER_132_1062 ();
 sg13g2_fill_1 FILLER_132_1064 ();
 sg13g2_fill_1 FILLER_132_1096 ();
 sg13g2_fill_2 FILLER_132_1107 ();
 sg13g2_fill_1 FILLER_132_1109 ();
 sg13g2_decap_4 FILLER_132_1115 ();
 sg13g2_decap_8 FILLER_132_1123 ();
 sg13g2_decap_8 FILLER_132_1130 ();
 sg13g2_decap_8 FILLER_132_1137 ();
 sg13g2_decap_8 FILLER_132_1144 ();
 sg13g2_decap_8 FILLER_132_1151 ();
 sg13g2_decap_8 FILLER_132_1158 ();
 sg13g2_decap_8 FILLER_132_1165 ();
 sg13g2_fill_2 FILLER_132_1193 ();
 sg13g2_fill_1 FILLER_132_1195 ();
 sg13g2_fill_1 FILLER_132_1204 ();
 sg13g2_fill_1 FILLER_132_1243 ();
 sg13g2_fill_1 FILLER_132_1252 ();
 sg13g2_fill_1 FILLER_132_1258 ();
 sg13g2_fill_1 FILLER_132_1271 ();
 sg13g2_decap_8 FILLER_132_1298 ();
 sg13g2_fill_2 FILLER_132_1305 ();
 sg13g2_decap_4 FILLER_132_1313 ();
 sg13g2_decap_4 FILLER_132_1323 ();
 sg13g2_decap_8 FILLER_132_1358 ();
 sg13g2_decap_4 FILLER_132_1365 ();
 sg13g2_decap_8 FILLER_132_1373 ();
 sg13g2_decap_8 FILLER_132_1380 ();
 sg13g2_decap_8 FILLER_132_1387 ();
 sg13g2_decap_8 FILLER_132_1394 ();
 sg13g2_decap_8 FILLER_132_1401 ();
 sg13g2_decap_8 FILLER_132_1408 ();
 sg13g2_decap_8 FILLER_132_1415 ();
 sg13g2_decap_8 FILLER_132_1422 ();
 sg13g2_decap_8 FILLER_132_1429 ();
 sg13g2_decap_8 FILLER_132_1436 ();
 sg13g2_decap_8 FILLER_132_1443 ();
 sg13g2_decap_8 FILLER_132_1450 ();
 sg13g2_decap_8 FILLER_132_1457 ();
 sg13g2_decap_8 FILLER_132_1464 ();
 sg13g2_decap_8 FILLER_132_1471 ();
 sg13g2_decap_8 FILLER_132_1478 ();
 sg13g2_decap_8 FILLER_132_1485 ();
 sg13g2_decap_8 FILLER_132_1492 ();
 sg13g2_decap_8 FILLER_132_1499 ();
 sg13g2_decap_8 FILLER_132_1506 ();
 sg13g2_decap_8 FILLER_132_1513 ();
 sg13g2_decap_8 FILLER_132_1520 ();
 sg13g2_decap_8 FILLER_132_1527 ();
 sg13g2_decap_8 FILLER_132_1534 ();
 sg13g2_decap_8 FILLER_132_1541 ();
 sg13g2_decap_8 FILLER_132_1548 ();
 sg13g2_decap_8 FILLER_132_1555 ();
 sg13g2_decap_8 FILLER_132_1562 ();
 sg13g2_decap_8 FILLER_132_1569 ();
 sg13g2_decap_8 FILLER_132_1576 ();
 sg13g2_decap_8 FILLER_132_1583 ();
 sg13g2_decap_8 FILLER_132_1590 ();
 sg13g2_decap_8 FILLER_132_1597 ();
 sg13g2_decap_8 FILLER_132_1604 ();
 sg13g2_decap_8 FILLER_132_1611 ();
 sg13g2_decap_8 FILLER_132_1618 ();
 sg13g2_decap_8 FILLER_133_0 ();
 sg13g2_decap_8 FILLER_133_7 ();
 sg13g2_decap_8 FILLER_133_14 ();
 sg13g2_decap_8 FILLER_133_21 ();
 sg13g2_decap_8 FILLER_133_28 ();
 sg13g2_decap_8 FILLER_133_35 ();
 sg13g2_decap_8 FILLER_133_42 ();
 sg13g2_fill_1 FILLER_133_49 ();
 sg13g2_decap_8 FILLER_133_54 ();
 sg13g2_fill_1 FILLER_133_61 ();
 sg13g2_fill_1 FILLER_133_90 ();
 sg13g2_fill_2 FILLER_133_165 ();
 sg13g2_decap_4 FILLER_133_171 ();
 sg13g2_decap_8 FILLER_133_207 ();
 sg13g2_fill_1 FILLER_133_214 ();
 sg13g2_fill_2 FILLER_133_220 ();
 sg13g2_fill_1 FILLER_133_222 ();
 sg13g2_decap_8 FILLER_133_241 ();
 sg13g2_decap_8 FILLER_133_248 ();
 sg13g2_decap_8 FILLER_133_255 ();
 sg13g2_decap_4 FILLER_133_275 ();
 sg13g2_fill_1 FILLER_133_279 ();
 sg13g2_fill_2 FILLER_133_289 ();
 sg13g2_decap_8 FILLER_133_303 ();
 sg13g2_fill_2 FILLER_133_310 ();
 sg13g2_fill_1 FILLER_133_312 ();
 sg13g2_fill_2 FILLER_133_354 ();
 sg13g2_fill_2 FILLER_133_363 ();
 sg13g2_fill_1 FILLER_133_365 ();
 sg13g2_decap_8 FILLER_133_379 ();
 sg13g2_decap_8 FILLER_133_386 ();
 sg13g2_decap_4 FILLER_133_393 ();
 sg13g2_fill_2 FILLER_133_401 ();
 sg13g2_fill_1 FILLER_133_403 ();
 sg13g2_fill_2 FILLER_133_415 ();
 sg13g2_decap_8 FILLER_133_443 ();
 sg13g2_decap_4 FILLER_133_450 ();
 sg13g2_fill_2 FILLER_133_454 ();
 sg13g2_decap_8 FILLER_133_481 ();
 sg13g2_decap_8 FILLER_133_488 ();
 sg13g2_fill_2 FILLER_133_495 ();
 sg13g2_fill_1 FILLER_133_497 ();
 sg13g2_fill_2 FILLER_133_502 ();
 sg13g2_decap_8 FILLER_133_542 ();
 sg13g2_fill_1 FILLER_133_561 ();
 sg13g2_decap_4 FILLER_133_568 ();
 sg13g2_fill_2 FILLER_133_572 ();
 sg13g2_decap_8 FILLER_133_586 ();
 sg13g2_decap_4 FILLER_133_593 ();
 sg13g2_fill_1 FILLER_133_597 ();
 sg13g2_decap_8 FILLER_133_602 ();
 sg13g2_fill_1 FILLER_133_622 ();
 sg13g2_fill_1 FILLER_133_628 ();
 sg13g2_decap_8 FILLER_133_633 ();
 sg13g2_decap_8 FILLER_133_640 ();
 sg13g2_decap_8 FILLER_133_647 ();
 sg13g2_decap_8 FILLER_133_654 ();
 sg13g2_decap_4 FILLER_133_661 ();
 sg13g2_fill_1 FILLER_133_665 ();
 sg13g2_decap_8 FILLER_133_675 ();
 sg13g2_decap_8 FILLER_133_682 ();
 sg13g2_decap_8 FILLER_133_689 ();
 sg13g2_decap_8 FILLER_133_696 ();
 sg13g2_decap_4 FILLER_133_703 ();
 sg13g2_fill_1 FILLER_133_707 ();
 sg13g2_decap_8 FILLER_133_712 ();
 sg13g2_decap_4 FILLER_133_719 ();
 sg13g2_fill_2 FILLER_133_723 ();
 sg13g2_fill_1 FILLER_133_781 ();
 sg13g2_decap_8 FILLER_133_833 ();
 sg13g2_decap_8 FILLER_133_840 ();
 sg13g2_fill_2 FILLER_133_847 ();
 sg13g2_fill_2 FILLER_133_858 ();
 sg13g2_decap_8 FILLER_133_864 ();
 sg13g2_decap_8 FILLER_133_871 ();
 sg13g2_fill_2 FILLER_133_893 ();
 sg13g2_decap_4 FILLER_133_899 ();
 sg13g2_fill_1 FILLER_133_903 ();
 sg13g2_decap_4 FILLER_133_909 ();
 sg13g2_decap_4 FILLER_133_939 ();
 sg13g2_decap_4 FILLER_133_955 ();
 sg13g2_fill_1 FILLER_133_959 ();
 sg13g2_decap_4 FILLER_133_964 ();
 sg13g2_fill_1 FILLER_133_968 ();
 sg13g2_fill_1 FILLER_133_974 ();
 sg13g2_decap_8 FILLER_133_993 ();
 sg13g2_decap_8 FILLER_133_1000 ();
 sg13g2_fill_2 FILLER_133_1013 ();
 sg13g2_fill_1 FILLER_133_1024 ();
 sg13g2_fill_1 FILLER_133_1034 ();
 sg13g2_fill_2 FILLER_133_1061 ();
 sg13g2_fill_1 FILLER_133_1063 ();
 sg13g2_decap_4 FILLER_133_1115 ();
 sg13g2_fill_1 FILLER_133_1119 ();
 sg13g2_decap_8 FILLER_133_1125 ();
 sg13g2_decap_8 FILLER_133_1132 ();
 sg13g2_fill_2 FILLER_133_1139 ();
 sg13g2_fill_1 FILLER_133_1141 ();
 sg13g2_decap_8 FILLER_133_1150 ();
 sg13g2_fill_2 FILLER_133_1157 ();
 sg13g2_fill_2 FILLER_133_1249 ();
 sg13g2_fill_1 FILLER_133_1251 ();
 sg13g2_decap_8 FILLER_133_1260 ();
 sg13g2_decap_8 FILLER_133_1267 ();
 sg13g2_decap_4 FILLER_133_1274 ();
 sg13g2_fill_2 FILLER_133_1278 ();
 sg13g2_decap_8 FILLER_133_1304 ();
 sg13g2_fill_1 FILLER_133_1311 ();
 sg13g2_fill_2 FILLER_133_1318 ();
 sg13g2_fill_1 FILLER_133_1320 ();
 sg13g2_decap_8 FILLER_133_1327 ();
 sg13g2_decap_8 FILLER_133_1334 ();
 sg13g2_decap_4 FILLER_133_1341 ();
 sg13g2_fill_1 FILLER_133_1345 ();
 sg13g2_decap_4 FILLER_133_1356 ();
 sg13g2_fill_1 FILLER_133_1360 ();
 sg13g2_decap_8 FILLER_133_1387 ();
 sg13g2_decap_8 FILLER_133_1394 ();
 sg13g2_decap_8 FILLER_133_1401 ();
 sg13g2_decap_8 FILLER_133_1408 ();
 sg13g2_decap_8 FILLER_133_1415 ();
 sg13g2_decap_8 FILLER_133_1422 ();
 sg13g2_decap_8 FILLER_133_1429 ();
 sg13g2_decap_8 FILLER_133_1436 ();
 sg13g2_decap_8 FILLER_133_1443 ();
 sg13g2_decap_8 FILLER_133_1450 ();
 sg13g2_decap_8 FILLER_133_1457 ();
 sg13g2_decap_8 FILLER_133_1464 ();
 sg13g2_decap_8 FILLER_133_1471 ();
 sg13g2_decap_8 FILLER_133_1478 ();
 sg13g2_decap_8 FILLER_133_1485 ();
 sg13g2_decap_8 FILLER_133_1492 ();
 sg13g2_decap_8 FILLER_133_1499 ();
 sg13g2_decap_8 FILLER_133_1506 ();
 sg13g2_decap_8 FILLER_133_1513 ();
 sg13g2_decap_8 FILLER_133_1520 ();
 sg13g2_decap_8 FILLER_133_1527 ();
 sg13g2_decap_8 FILLER_133_1534 ();
 sg13g2_decap_8 FILLER_133_1541 ();
 sg13g2_decap_8 FILLER_133_1548 ();
 sg13g2_decap_8 FILLER_133_1555 ();
 sg13g2_decap_8 FILLER_133_1562 ();
 sg13g2_decap_8 FILLER_133_1569 ();
 sg13g2_decap_8 FILLER_133_1576 ();
 sg13g2_decap_8 FILLER_133_1583 ();
 sg13g2_decap_8 FILLER_133_1590 ();
 sg13g2_decap_8 FILLER_133_1597 ();
 sg13g2_decap_8 FILLER_133_1604 ();
 sg13g2_decap_8 FILLER_133_1611 ();
 sg13g2_decap_8 FILLER_133_1618 ();
 sg13g2_decap_8 FILLER_134_0 ();
 sg13g2_decap_8 FILLER_134_11 ();
 sg13g2_decap_8 FILLER_134_18 ();
 sg13g2_decap_8 FILLER_134_25 ();
 sg13g2_fill_2 FILLER_134_32 ();
 sg13g2_fill_2 FILLER_134_38 ();
 sg13g2_decap_4 FILLER_134_69 ();
 sg13g2_fill_1 FILLER_134_77 ();
 sg13g2_fill_1 FILLER_134_86 ();
 sg13g2_fill_1 FILLER_134_117 ();
 sg13g2_decap_4 FILLER_134_149 ();
 sg13g2_fill_1 FILLER_134_153 ();
 sg13g2_fill_2 FILLER_134_185 ();
 sg13g2_fill_1 FILLER_134_187 ();
 sg13g2_decap_8 FILLER_134_192 ();
 sg13g2_decap_8 FILLER_134_199 ();
 sg13g2_fill_1 FILLER_134_206 ();
 sg13g2_fill_1 FILLER_134_219 ();
 sg13g2_fill_2 FILLER_134_230 ();
 sg13g2_decap_8 FILLER_134_244 ();
 sg13g2_decap_8 FILLER_134_251 ();
 sg13g2_decap_8 FILLER_134_258 ();
 sg13g2_decap_4 FILLER_134_265 ();
 sg13g2_fill_1 FILLER_134_269 ();
 sg13g2_fill_2 FILLER_134_282 ();
 sg13g2_fill_1 FILLER_134_284 ();
 sg13g2_decap_8 FILLER_134_300 ();
 sg13g2_decap_4 FILLER_134_307 ();
 sg13g2_fill_2 FILLER_134_346 ();
 sg13g2_fill_2 FILLER_134_358 ();
 sg13g2_decap_4 FILLER_134_365 ();
 sg13g2_decap_8 FILLER_134_382 ();
 sg13g2_decap_8 FILLER_134_389 ();
 sg13g2_fill_2 FILLER_134_396 ();
 sg13g2_fill_2 FILLER_134_404 ();
 sg13g2_fill_1 FILLER_134_406 ();
 sg13g2_decap_8 FILLER_134_411 ();
 sg13g2_decap_8 FILLER_134_418 ();
 sg13g2_fill_1 FILLER_134_425 ();
 sg13g2_fill_1 FILLER_134_438 ();
 sg13g2_decap_8 FILLER_134_444 ();
 sg13g2_decap_8 FILLER_134_451 ();
 sg13g2_fill_2 FILLER_134_458 ();
 sg13g2_fill_1 FILLER_134_460 ();
 sg13g2_decap_4 FILLER_134_468 ();
 sg13g2_fill_1 FILLER_134_472 ();
 sg13g2_decap_8 FILLER_134_478 ();
 sg13g2_decap_8 FILLER_134_490 ();
 sg13g2_decap_4 FILLER_134_497 ();
 sg13g2_fill_1 FILLER_134_501 ();
 sg13g2_fill_1 FILLER_134_528 ();
 sg13g2_decap_4 FILLER_134_537 ();
 sg13g2_fill_2 FILLER_134_541 ();
 sg13g2_decap_4 FILLER_134_569 ();
 sg13g2_fill_2 FILLER_134_573 ();
 sg13g2_decap_8 FILLER_134_581 ();
 sg13g2_fill_2 FILLER_134_588 ();
 sg13g2_fill_1 FILLER_134_590 ();
 sg13g2_decap_4 FILLER_134_620 ();
 sg13g2_decap_4 FILLER_134_653 ();
 sg13g2_decap_4 FILLER_134_666 ();
 sg13g2_fill_2 FILLER_134_678 ();
 sg13g2_fill_2 FILLER_134_689 ();
 sg13g2_fill_1 FILLER_134_691 ();
 sg13g2_decap_4 FILLER_134_696 ();
 sg13g2_fill_2 FILLER_134_700 ();
 sg13g2_fill_1 FILLER_134_784 ();
 sg13g2_fill_2 FILLER_134_789 ();
 sg13g2_fill_1 FILLER_134_791 ();
 sg13g2_fill_2 FILLER_134_821 ();
 sg13g2_fill_1 FILLER_134_823 ();
 sg13g2_decap_8 FILLER_134_837 ();
 sg13g2_fill_1 FILLER_134_844 ();
 sg13g2_decap_8 FILLER_134_876 ();
 sg13g2_decap_4 FILLER_134_883 ();
 sg13g2_decap_4 FILLER_134_921 ();
 sg13g2_decap_8 FILLER_134_953 ();
 sg13g2_fill_2 FILLER_134_965 ();
 sg13g2_fill_2 FILLER_134_972 ();
 sg13g2_decap_4 FILLER_134_978 ();
 sg13g2_decap_8 FILLER_134_1010 ();
 sg13g2_decap_8 FILLER_134_1017 ();
 sg13g2_decap_8 FILLER_134_1024 ();
 sg13g2_decap_8 FILLER_134_1031 ();
 sg13g2_decap_8 FILLER_134_1038 ();
 sg13g2_decap_8 FILLER_134_1045 ();
 sg13g2_fill_1 FILLER_134_1052 ();
 sg13g2_decap_8 FILLER_134_1057 ();
 sg13g2_fill_2 FILLER_134_1064 ();
 sg13g2_fill_1 FILLER_134_1066 ();
 sg13g2_fill_1 FILLER_134_1076 ();
 sg13g2_fill_2 FILLER_134_1087 ();
 sg13g2_fill_1 FILLER_134_1089 ();
 sg13g2_decap_4 FILLER_134_1094 ();
 sg13g2_fill_1 FILLER_134_1098 ();
 sg13g2_decap_8 FILLER_134_1104 ();
 sg13g2_fill_1 FILLER_134_1111 ();
 sg13g2_fill_2 FILLER_134_1125 ();
 sg13g2_fill_2 FILLER_134_1135 ();
 sg13g2_fill_1 FILLER_134_1137 ();
 sg13g2_decap_8 FILLER_134_1151 ();
 sg13g2_decap_4 FILLER_134_1166 ();
 sg13g2_decap_4 FILLER_134_1174 ();
 sg13g2_fill_2 FILLER_134_1178 ();
 sg13g2_fill_2 FILLER_134_1188 ();
 sg13g2_fill_1 FILLER_134_1190 ();
 sg13g2_fill_2 FILLER_134_1281 ();
 sg13g2_decap_4 FILLER_134_1289 ();
 sg13g2_fill_1 FILLER_134_1293 ();
 sg13g2_decap_4 FILLER_134_1306 ();
 sg13g2_fill_1 FILLER_134_1310 ();
 sg13g2_fill_1 FILLER_134_1316 ();
 sg13g2_decap_8 FILLER_134_1323 ();
 sg13g2_decap_4 FILLER_134_1330 ();
 sg13g2_fill_1 FILLER_134_1334 ();
 sg13g2_fill_1 FILLER_134_1345 ();
 sg13g2_decap_8 FILLER_134_1350 ();
 sg13g2_decap_4 FILLER_134_1357 ();
 sg13g2_fill_1 FILLER_134_1361 ();
 sg13g2_decap_8 FILLER_134_1365 ();
 sg13g2_decap_8 FILLER_134_1372 ();
 sg13g2_decap_8 FILLER_134_1379 ();
 sg13g2_decap_8 FILLER_134_1386 ();
 sg13g2_decap_8 FILLER_134_1393 ();
 sg13g2_decap_8 FILLER_134_1400 ();
 sg13g2_decap_8 FILLER_134_1407 ();
 sg13g2_decap_8 FILLER_134_1414 ();
 sg13g2_decap_8 FILLER_134_1421 ();
 sg13g2_decap_8 FILLER_134_1428 ();
 sg13g2_decap_8 FILLER_134_1435 ();
 sg13g2_decap_8 FILLER_134_1442 ();
 sg13g2_decap_8 FILLER_134_1449 ();
 sg13g2_decap_8 FILLER_134_1456 ();
 sg13g2_decap_8 FILLER_134_1463 ();
 sg13g2_decap_8 FILLER_134_1470 ();
 sg13g2_decap_8 FILLER_134_1477 ();
 sg13g2_decap_8 FILLER_134_1484 ();
 sg13g2_decap_8 FILLER_134_1491 ();
 sg13g2_decap_8 FILLER_134_1498 ();
 sg13g2_decap_8 FILLER_134_1505 ();
 sg13g2_decap_8 FILLER_134_1512 ();
 sg13g2_decap_8 FILLER_134_1519 ();
 sg13g2_decap_8 FILLER_134_1526 ();
 sg13g2_decap_8 FILLER_134_1533 ();
 sg13g2_decap_8 FILLER_134_1540 ();
 sg13g2_decap_8 FILLER_134_1547 ();
 sg13g2_decap_8 FILLER_134_1554 ();
 sg13g2_decap_8 FILLER_134_1561 ();
 sg13g2_decap_8 FILLER_134_1568 ();
 sg13g2_decap_8 FILLER_134_1575 ();
 sg13g2_decap_8 FILLER_134_1582 ();
 sg13g2_decap_8 FILLER_134_1589 ();
 sg13g2_decap_8 FILLER_134_1596 ();
 sg13g2_decap_8 FILLER_134_1603 ();
 sg13g2_decap_8 FILLER_134_1610 ();
 sg13g2_decap_8 FILLER_134_1617 ();
 sg13g2_fill_1 FILLER_134_1624 ();
 sg13g2_fill_1 FILLER_135_0 ();
 sg13g2_fill_1 FILLER_135_60 ();
 sg13g2_fill_1 FILLER_135_120 ();
 sg13g2_decap_8 FILLER_135_155 ();
 sg13g2_fill_2 FILLER_135_162 ();
 sg13g2_decap_4 FILLER_135_173 ();
 sg13g2_decap_8 FILLER_135_202 ();
 sg13g2_fill_2 FILLER_135_209 ();
 sg13g2_fill_1 FILLER_135_211 ();
 sg13g2_fill_1 FILLER_135_217 ();
 sg13g2_fill_2 FILLER_135_227 ();
 sg13g2_fill_1 FILLER_135_234 ();
 sg13g2_fill_2 FILLER_135_243 ();
 sg13g2_fill_1 FILLER_135_255 ();
 sg13g2_fill_2 FILLER_135_264 ();
 sg13g2_fill_2 FILLER_135_299 ();
 sg13g2_fill_1 FILLER_135_301 ();
 sg13g2_decap_8 FILLER_135_307 ();
 sg13g2_decap_8 FILLER_135_314 ();
 sg13g2_decap_8 FILLER_135_321 ();
 sg13g2_decap_8 FILLER_135_328 ();
 sg13g2_fill_2 FILLER_135_335 ();
 sg13g2_fill_1 FILLER_135_337 ();
 sg13g2_decap_8 FILLER_135_344 ();
 sg13g2_decap_8 FILLER_135_361 ();
 sg13g2_fill_2 FILLER_135_368 ();
 sg13g2_decap_8 FILLER_135_382 ();
 sg13g2_decap_4 FILLER_135_389 ();
 sg13g2_fill_1 FILLER_135_393 ();
 sg13g2_decap_4 FILLER_135_430 ();
 sg13g2_decap_8 FILLER_135_439 ();
 sg13g2_fill_2 FILLER_135_446 ();
 sg13g2_fill_2 FILLER_135_457 ();
 sg13g2_fill_1 FILLER_135_469 ();
 sg13g2_decap_8 FILLER_135_475 ();
 sg13g2_fill_1 FILLER_135_482 ();
 sg13g2_decap_8 FILLER_135_488 ();
 sg13g2_decap_8 FILLER_135_495 ();
 sg13g2_decap_4 FILLER_135_502 ();
 sg13g2_decap_4 FILLER_135_511 ();
 sg13g2_fill_2 FILLER_135_532 ();
 sg13g2_fill_2 FILLER_135_537 ();
 sg13g2_fill_1 FILLER_135_539 ();
 sg13g2_fill_1 FILLER_135_546 ();
 sg13g2_fill_2 FILLER_135_559 ();
 sg13g2_fill_1 FILLER_135_561 ();
 sg13g2_decap_8 FILLER_135_579 ();
 sg13g2_fill_2 FILLER_135_586 ();
 sg13g2_fill_2 FILLER_135_596 ();
 sg13g2_fill_1 FILLER_135_598 ();
 sg13g2_decap_4 FILLER_135_604 ();
 sg13g2_decap_4 FILLER_135_612 ();
 sg13g2_decap_8 FILLER_135_625 ();
 sg13g2_fill_2 FILLER_135_632 ();
 sg13g2_fill_1 FILLER_135_634 ();
 sg13g2_fill_1 FILLER_135_661 ();
 sg13g2_decap_4 FILLER_135_678 ();
 sg13g2_fill_1 FILLER_135_682 ();
 sg13g2_decap_4 FILLER_135_709 ();
 sg13g2_fill_2 FILLER_135_804 ();
 sg13g2_decap_8 FILLER_135_811 ();
 sg13g2_decap_8 FILLER_135_818 ();
 sg13g2_fill_1 FILLER_135_825 ();
 sg13g2_decap_4 FILLER_135_852 ();
 sg13g2_fill_1 FILLER_135_856 ();
 sg13g2_decap_8 FILLER_135_861 ();
 sg13g2_fill_1 FILLER_135_868 ();
 sg13g2_decap_8 FILLER_135_874 ();
 sg13g2_decap_8 FILLER_135_881 ();
 sg13g2_decap_4 FILLER_135_888 ();
 sg13g2_fill_1 FILLER_135_892 ();
 sg13g2_decap_4 FILLER_135_897 ();
 sg13g2_fill_2 FILLER_135_901 ();
 sg13g2_fill_1 FILLER_135_916 ();
 sg13g2_decap_8 FILLER_135_961 ();
 sg13g2_fill_2 FILLER_135_968 ();
 sg13g2_fill_1 FILLER_135_970 ();
 sg13g2_fill_1 FILLER_135_976 ();
 sg13g2_decap_4 FILLER_135_1006 ();
 sg13g2_fill_2 FILLER_135_1015 ();
 sg13g2_decap_4 FILLER_135_1029 ();
 sg13g2_fill_2 FILLER_135_1033 ();
 sg13g2_fill_2 FILLER_135_1042 ();
 sg13g2_fill_1 FILLER_135_1044 ();
 sg13g2_fill_2 FILLER_135_1077 ();
 sg13g2_fill_1 FILLER_135_1079 ();
 sg13g2_fill_2 FILLER_135_1087 ();
 sg13g2_decap_8 FILLER_135_1102 ();
 sg13g2_decap_4 FILLER_135_1109 ();
 sg13g2_fill_1 FILLER_135_1162 ();
 sg13g2_decap_8 FILLER_135_1171 ();
 sg13g2_decap_8 FILLER_135_1178 ();
 sg13g2_decap_8 FILLER_135_1244 ();
 sg13g2_fill_2 FILLER_135_1251 ();
 sg13g2_fill_1 FILLER_135_1288 ();
 sg13g2_decap_8 FILLER_135_1293 ();
 sg13g2_decap_8 FILLER_135_1300 ();
 sg13g2_decap_4 FILLER_135_1307 ();
 sg13g2_decap_4 FILLER_135_1315 ();
 sg13g2_decap_8 FILLER_135_1329 ();
 sg13g2_fill_2 FILLER_135_1336 ();
 sg13g2_decap_8 FILLER_135_1389 ();
 sg13g2_decap_8 FILLER_135_1396 ();
 sg13g2_decap_8 FILLER_135_1403 ();
 sg13g2_decap_8 FILLER_135_1410 ();
 sg13g2_decap_8 FILLER_135_1417 ();
 sg13g2_decap_8 FILLER_135_1424 ();
 sg13g2_decap_8 FILLER_135_1431 ();
 sg13g2_decap_8 FILLER_135_1438 ();
 sg13g2_decap_8 FILLER_135_1445 ();
 sg13g2_decap_8 FILLER_135_1452 ();
 sg13g2_decap_8 FILLER_135_1459 ();
 sg13g2_decap_8 FILLER_135_1466 ();
 sg13g2_decap_8 FILLER_135_1473 ();
 sg13g2_decap_8 FILLER_135_1480 ();
 sg13g2_decap_8 FILLER_135_1487 ();
 sg13g2_decap_8 FILLER_135_1494 ();
 sg13g2_decap_8 FILLER_135_1501 ();
 sg13g2_decap_8 FILLER_135_1508 ();
 sg13g2_decap_8 FILLER_135_1515 ();
 sg13g2_decap_8 FILLER_135_1522 ();
 sg13g2_decap_8 FILLER_135_1529 ();
 sg13g2_decap_8 FILLER_135_1536 ();
 sg13g2_decap_8 FILLER_135_1543 ();
 sg13g2_decap_8 FILLER_135_1550 ();
 sg13g2_decap_8 FILLER_135_1557 ();
 sg13g2_decap_8 FILLER_135_1564 ();
 sg13g2_decap_8 FILLER_135_1571 ();
 sg13g2_decap_8 FILLER_135_1578 ();
 sg13g2_decap_8 FILLER_135_1585 ();
 sg13g2_decap_8 FILLER_135_1592 ();
 sg13g2_decap_8 FILLER_135_1599 ();
 sg13g2_decap_8 FILLER_135_1606 ();
 sg13g2_decap_8 FILLER_135_1613 ();
 sg13g2_decap_4 FILLER_135_1620 ();
 sg13g2_fill_1 FILLER_135_1624 ();
 sg13g2_decap_8 FILLER_136_0 ();
 sg13g2_fill_1 FILLER_136_7 ();
 sg13g2_fill_2 FILLER_136_12 ();
 sg13g2_fill_1 FILLER_136_19 ();
 sg13g2_decap_8 FILLER_136_30 ();
 sg13g2_decap_4 FILLER_136_37 ();
 sg13g2_fill_1 FILLER_136_41 ();
 sg13g2_fill_1 FILLER_136_86 ();
 sg13g2_decap_4 FILLER_136_131 ();
 sg13g2_decap_8 FILLER_136_171 ();
 sg13g2_decap_4 FILLER_136_178 ();
 sg13g2_decap_8 FILLER_136_186 ();
 sg13g2_decap_8 FILLER_136_193 ();
 sg13g2_decap_4 FILLER_136_200 ();
 sg13g2_fill_1 FILLER_136_210 ();
 sg13g2_fill_1 FILLER_136_225 ();
 sg13g2_fill_1 FILLER_136_230 ();
 sg13g2_fill_1 FILLER_136_240 ();
 sg13g2_decap_8 FILLER_136_245 ();
 sg13g2_decap_8 FILLER_136_252 ();
 sg13g2_decap_8 FILLER_136_259 ();
 sg13g2_decap_4 FILLER_136_266 ();
 sg13g2_fill_1 FILLER_136_270 ();
 sg13g2_fill_1 FILLER_136_307 ();
 sg13g2_decap_8 FILLER_136_313 ();
 sg13g2_fill_2 FILLER_136_320 ();
 sg13g2_fill_1 FILLER_136_322 ();
 sg13g2_decap_4 FILLER_136_327 ();
 sg13g2_fill_2 FILLER_136_331 ();
 sg13g2_decap_8 FILLER_136_338 ();
 sg13g2_decap_4 FILLER_136_345 ();
 sg13g2_fill_2 FILLER_136_363 ();
 sg13g2_fill_1 FILLER_136_365 ();
 sg13g2_decap_8 FILLER_136_385 ();
 sg13g2_decap_4 FILLER_136_392 ();
 sg13g2_fill_1 FILLER_136_396 ();
 sg13g2_decap_8 FILLER_136_411 ();
 sg13g2_decap_4 FILLER_136_418 ();
 sg13g2_fill_1 FILLER_136_422 ();
 sg13g2_decap_4 FILLER_136_441 ();
 sg13g2_decap_4 FILLER_136_449 ();
 sg13g2_fill_2 FILLER_136_466 ();
 sg13g2_fill_1 FILLER_136_468 ();
 sg13g2_decap_4 FILLER_136_478 ();
 sg13g2_fill_2 FILLER_136_482 ();
 sg13g2_decap_4 FILLER_136_492 ();
 sg13g2_fill_2 FILLER_136_505 ();
 sg13g2_fill_2 FILLER_136_511 ();
 sg13g2_fill_1 FILLER_136_513 ();
 sg13g2_decap_8 FILLER_136_537 ();
 sg13g2_decap_4 FILLER_136_544 ();
 sg13g2_fill_1 FILLER_136_553 ();
 sg13g2_fill_2 FILLER_136_572 ();
 sg13g2_fill_2 FILLER_136_580 ();
 sg13g2_decap_8 FILLER_136_591 ();
 sg13g2_fill_2 FILLER_136_598 ();
 sg13g2_decap_4 FILLER_136_626 ();
 sg13g2_fill_1 FILLER_136_630 ();
 sg13g2_decap_8 FILLER_136_636 ();
 sg13g2_fill_1 FILLER_136_643 ();
 sg13g2_decap_8 FILLER_136_649 ();
 sg13g2_decap_4 FILLER_136_656 ();
 sg13g2_fill_2 FILLER_136_660 ();
 sg13g2_decap_4 FILLER_136_666 ();
 sg13g2_decap_8 FILLER_136_679 ();
 sg13g2_decap_8 FILLER_136_686 ();
 sg13g2_decap_8 FILLER_136_693 ();
 sg13g2_decap_4 FILLER_136_700 ();
 sg13g2_fill_2 FILLER_136_704 ();
 sg13g2_fill_2 FILLER_136_731 ();
 sg13g2_decap_4 FILLER_136_799 ();
 sg13g2_decap_8 FILLER_136_814 ();
 sg13g2_decap_8 FILLER_136_821 ();
 sg13g2_decap_8 FILLER_136_828 ();
 sg13g2_decap_8 FILLER_136_835 ();
 sg13g2_fill_1 FILLER_136_842 ();
 sg13g2_decap_8 FILLER_136_853 ();
 sg13g2_fill_1 FILLER_136_860 ();
 sg13g2_decap_8 FILLER_136_881 ();
 sg13g2_decap_8 FILLER_136_945 ();
 sg13g2_fill_2 FILLER_136_952 ();
 sg13g2_fill_1 FILLER_136_954 ();
 sg13g2_decap_8 FILLER_136_959 ();
 sg13g2_decap_8 FILLER_136_966 ();
 sg13g2_fill_1 FILLER_136_973 ();
 sg13g2_fill_2 FILLER_136_978 ();
 sg13g2_fill_1 FILLER_136_980 ();
 sg13g2_decap_8 FILLER_136_990 ();
 sg13g2_fill_2 FILLER_136_997 ();
 sg13g2_fill_1 FILLER_136_999 ();
 sg13g2_fill_2 FILLER_136_1035 ();
 sg13g2_fill_1 FILLER_136_1037 ();
 sg13g2_decap_8 FILLER_136_1105 ();
 sg13g2_decap_8 FILLER_136_1112 ();
 sg13g2_decap_8 FILLER_136_1119 ();
 sg13g2_fill_1 FILLER_136_1131 ();
 sg13g2_fill_1 FILLER_136_1137 ();
 sg13g2_fill_2 FILLER_136_1167 ();
 sg13g2_fill_1 FILLER_136_1175 ();
 sg13g2_fill_1 FILLER_136_1180 ();
 sg13g2_fill_1 FILLER_136_1189 ();
 sg13g2_fill_2 FILLER_136_1198 ();
 sg13g2_fill_1 FILLER_136_1205 ();
 sg13g2_decap_8 FILLER_136_1243 ();
 sg13g2_fill_2 FILLER_136_1250 ();
 sg13g2_decap_8 FILLER_136_1307 ();
 sg13g2_fill_1 FILLER_136_1314 ();
 sg13g2_decap_8 FILLER_136_1322 ();
 sg13g2_decap_8 FILLER_136_1329 ();
 sg13g2_decap_8 FILLER_136_1336 ();
 sg13g2_decap_8 FILLER_136_1343 ();
 sg13g2_decap_8 FILLER_136_1350 ();
 sg13g2_decap_8 FILLER_136_1357 ();
 sg13g2_decap_8 FILLER_136_1364 ();
 sg13g2_decap_8 FILLER_136_1371 ();
 sg13g2_decap_8 FILLER_136_1378 ();
 sg13g2_decap_8 FILLER_136_1385 ();
 sg13g2_decap_8 FILLER_136_1392 ();
 sg13g2_decap_8 FILLER_136_1399 ();
 sg13g2_decap_8 FILLER_136_1406 ();
 sg13g2_decap_8 FILLER_136_1413 ();
 sg13g2_decap_8 FILLER_136_1420 ();
 sg13g2_decap_8 FILLER_136_1427 ();
 sg13g2_decap_8 FILLER_136_1434 ();
 sg13g2_decap_8 FILLER_136_1441 ();
 sg13g2_decap_8 FILLER_136_1448 ();
 sg13g2_decap_8 FILLER_136_1455 ();
 sg13g2_decap_8 FILLER_136_1462 ();
 sg13g2_decap_8 FILLER_136_1469 ();
 sg13g2_decap_8 FILLER_136_1476 ();
 sg13g2_decap_8 FILLER_136_1483 ();
 sg13g2_decap_8 FILLER_136_1490 ();
 sg13g2_decap_8 FILLER_136_1497 ();
 sg13g2_decap_8 FILLER_136_1504 ();
 sg13g2_decap_8 FILLER_136_1511 ();
 sg13g2_decap_8 FILLER_136_1518 ();
 sg13g2_decap_8 FILLER_136_1525 ();
 sg13g2_decap_8 FILLER_136_1532 ();
 sg13g2_decap_8 FILLER_136_1539 ();
 sg13g2_decap_8 FILLER_136_1546 ();
 sg13g2_decap_8 FILLER_136_1553 ();
 sg13g2_decap_8 FILLER_136_1560 ();
 sg13g2_decap_8 FILLER_136_1567 ();
 sg13g2_decap_8 FILLER_136_1574 ();
 sg13g2_decap_8 FILLER_136_1581 ();
 sg13g2_decap_8 FILLER_136_1588 ();
 sg13g2_decap_8 FILLER_136_1595 ();
 sg13g2_decap_8 FILLER_136_1602 ();
 sg13g2_decap_8 FILLER_136_1609 ();
 sg13g2_decap_8 FILLER_136_1616 ();
 sg13g2_fill_2 FILLER_136_1623 ();
 sg13g2_fill_1 FILLER_137_0 ();
 sg13g2_decap_8 FILLER_137_33 ();
 sg13g2_decap_8 FILLER_137_40 ();
 sg13g2_fill_1 FILLER_137_51 ();
 sg13g2_fill_1 FILLER_137_78 ();
 sg13g2_fill_1 FILLER_137_144 ();
 sg13g2_decap_8 FILLER_137_205 ();
 sg13g2_decap_4 FILLER_137_228 ();
 sg13g2_decap_4 FILLER_137_251 ();
 sg13g2_fill_1 FILLER_137_255 ();
 sg13g2_decap_8 FILLER_137_260 ();
 sg13g2_decap_8 FILLER_137_267 ();
 sg13g2_decap_4 FILLER_137_274 ();
 sg13g2_decap_8 FILLER_137_282 ();
 sg13g2_decap_8 FILLER_137_289 ();
 sg13g2_fill_1 FILLER_137_296 ();
 sg13g2_decap_4 FILLER_137_309 ();
 sg13g2_fill_2 FILLER_137_313 ();
 sg13g2_decap_8 FILLER_137_341 ();
 sg13g2_fill_2 FILLER_137_348 ();
 sg13g2_fill_1 FILLER_137_350 ();
 sg13g2_decap_8 FILLER_137_360 ();
 sg13g2_decap_4 FILLER_137_367 ();
 sg13g2_decap_4 FILLER_137_386 ();
 sg13g2_fill_2 FILLER_137_390 ();
 sg13g2_fill_2 FILLER_137_428 ();
 sg13g2_fill_1 FILLER_137_430 ();
 sg13g2_decap_8 FILLER_137_441 ();
 sg13g2_decap_8 FILLER_137_448 ();
 sg13g2_decap_8 FILLER_137_455 ();
 sg13g2_fill_1 FILLER_137_462 ();
 sg13g2_decap_8 FILLER_137_474 ();
 sg13g2_decap_4 FILLER_137_481 ();
 sg13g2_decap_8 FILLER_137_490 ();
 sg13g2_fill_2 FILLER_137_497 ();
 sg13g2_fill_1 FILLER_137_499 ();
 sg13g2_decap_8 FILLER_137_532 ();
 sg13g2_decap_4 FILLER_137_545 ();
 sg13g2_fill_2 FILLER_137_549 ();
 sg13g2_fill_1 FILLER_137_555 ();
 sg13g2_decap_8 FILLER_137_574 ();
 sg13g2_decap_8 FILLER_137_581 ();
 sg13g2_decap_8 FILLER_137_588 ();
 sg13g2_decap_8 FILLER_137_595 ();
 sg13g2_decap_8 FILLER_137_602 ();
 sg13g2_fill_2 FILLER_137_609 ();
 sg13g2_fill_1 FILLER_137_611 ();
 sg13g2_fill_1 FILLER_137_646 ();
 sg13g2_decap_8 FILLER_137_681 ();
 sg13g2_decap_8 FILLER_137_688 ();
 sg13g2_decap_8 FILLER_137_695 ();
 sg13g2_fill_2 FILLER_137_702 ();
 sg13g2_fill_1 FILLER_137_704 ();
 sg13g2_fill_2 FILLER_137_774 ();
 sg13g2_fill_2 FILLER_137_784 ();
 sg13g2_fill_2 FILLER_137_794 ();
 sg13g2_fill_1 FILLER_137_796 ();
 sg13g2_decap_4 FILLER_137_828 ();
 sg13g2_fill_2 FILLER_137_832 ();
 sg13g2_decap_4 FILLER_137_859 ();
 sg13g2_decap_4 FILLER_137_868 ();
 sg13g2_decap_8 FILLER_137_876 ();
 sg13g2_fill_2 FILLER_137_883 ();
 sg13g2_fill_1 FILLER_137_885 ();
 sg13g2_decap_8 FILLER_137_917 ();
 sg13g2_decap_8 FILLER_137_924 ();
 sg13g2_decap_4 FILLER_137_931 ();
 sg13g2_fill_2 FILLER_137_935 ();
 sg13g2_decap_4 FILLER_137_941 ();
 sg13g2_fill_2 FILLER_137_945 ();
 sg13g2_decap_8 FILLER_137_973 ();
 sg13g2_decap_8 FILLER_137_980 ();
 sg13g2_fill_1 FILLER_137_987 ();
 sg13g2_decap_8 FILLER_137_1016 ();
 sg13g2_decap_8 FILLER_137_1023 ();
 sg13g2_fill_2 FILLER_137_1030 ();
 sg13g2_fill_1 FILLER_137_1032 ();
 sg13g2_decap_4 FILLER_137_1041 ();
 sg13g2_fill_2 FILLER_137_1045 ();
 sg13g2_decap_8 FILLER_137_1116 ();
 sg13g2_fill_2 FILLER_137_1123 ();
 sg13g2_fill_1 FILLER_137_1125 ();
 sg13g2_decap_4 FILLER_137_1132 ();
 sg13g2_fill_1 FILLER_137_1136 ();
 sg13g2_decap_8 FILLER_137_1142 ();
 sg13g2_decap_4 FILLER_137_1149 ();
 sg13g2_fill_2 FILLER_137_1153 ();
 sg13g2_fill_2 FILLER_137_1168 ();
 sg13g2_fill_1 FILLER_137_1170 ();
 sg13g2_decap_4 FILLER_137_1197 ();
 sg13g2_fill_2 FILLER_137_1201 ();
 sg13g2_fill_1 FILLER_137_1229 ();
 sg13g2_fill_1 FILLER_137_1234 ();
 sg13g2_decap_8 FILLER_137_1241 ();
 sg13g2_decap_8 FILLER_137_1303 ();
 sg13g2_decap_8 FILLER_137_1336 ();
 sg13g2_decap_8 FILLER_137_1343 ();
 sg13g2_decap_8 FILLER_137_1350 ();
 sg13g2_decap_8 FILLER_137_1357 ();
 sg13g2_decap_8 FILLER_137_1364 ();
 sg13g2_decap_8 FILLER_137_1371 ();
 sg13g2_decap_8 FILLER_137_1378 ();
 sg13g2_decap_8 FILLER_137_1385 ();
 sg13g2_decap_8 FILLER_137_1392 ();
 sg13g2_decap_8 FILLER_137_1399 ();
 sg13g2_decap_8 FILLER_137_1406 ();
 sg13g2_decap_8 FILLER_137_1413 ();
 sg13g2_decap_8 FILLER_137_1420 ();
 sg13g2_decap_8 FILLER_137_1427 ();
 sg13g2_decap_8 FILLER_137_1434 ();
 sg13g2_decap_8 FILLER_137_1441 ();
 sg13g2_decap_8 FILLER_137_1448 ();
 sg13g2_decap_8 FILLER_137_1455 ();
 sg13g2_decap_8 FILLER_137_1462 ();
 sg13g2_decap_8 FILLER_137_1469 ();
 sg13g2_decap_8 FILLER_137_1476 ();
 sg13g2_decap_8 FILLER_137_1483 ();
 sg13g2_decap_8 FILLER_137_1490 ();
 sg13g2_decap_8 FILLER_137_1497 ();
 sg13g2_decap_8 FILLER_137_1504 ();
 sg13g2_decap_8 FILLER_137_1511 ();
 sg13g2_decap_8 FILLER_137_1518 ();
 sg13g2_decap_8 FILLER_137_1525 ();
 sg13g2_decap_8 FILLER_137_1532 ();
 sg13g2_decap_8 FILLER_137_1539 ();
 sg13g2_decap_8 FILLER_137_1546 ();
 sg13g2_decap_8 FILLER_137_1553 ();
 sg13g2_decap_8 FILLER_137_1560 ();
 sg13g2_decap_8 FILLER_137_1567 ();
 sg13g2_decap_8 FILLER_137_1574 ();
 sg13g2_decap_8 FILLER_137_1581 ();
 sg13g2_decap_8 FILLER_137_1588 ();
 sg13g2_decap_8 FILLER_137_1595 ();
 sg13g2_decap_8 FILLER_137_1602 ();
 sg13g2_decap_8 FILLER_137_1609 ();
 sg13g2_decap_8 FILLER_137_1616 ();
 sg13g2_fill_2 FILLER_137_1623 ();
 sg13g2_fill_2 FILLER_138_0 ();
 sg13g2_fill_2 FILLER_138_32 ();
 sg13g2_fill_1 FILLER_138_34 ();
 sg13g2_fill_2 FILLER_138_84 ();
 sg13g2_fill_1 FILLER_138_103 ();
 sg13g2_decap_8 FILLER_138_108 ();
 sg13g2_decap_8 FILLER_138_115 ();
 sg13g2_decap_4 FILLER_138_122 ();
 sg13g2_decap_4 FILLER_138_130 ();
 sg13g2_decap_4 FILLER_138_175 ();
 sg13g2_decap_8 FILLER_138_192 ();
 sg13g2_decap_4 FILLER_138_199 ();
 sg13g2_fill_1 FILLER_138_203 ();
 sg13g2_decap_8 FILLER_138_211 ();
 sg13g2_fill_2 FILLER_138_218 ();
 sg13g2_fill_1 FILLER_138_220 ();
 sg13g2_decap_8 FILLER_138_233 ();
 sg13g2_fill_1 FILLER_138_240 ();
 sg13g2_fill_1 FILLER_138_246 ();
 sg13g2_decap_8 FILLER_138_273 ();
 sg13g2_fill_1 FILLER_138_280 ();
 sg13g2_decap_8 FILLER_138_286 ();
 sg13g2_decap_4 FILLER_138_318 ();
 sg13g2_decap_8 FILLER_138_327 ();
 sg13g2_decap_8 FILLER_138_334 ();
 sg13g2_decap_8 FILLER_138_341 ();
 sg13g2_fill_1 FILLER_138_374 ();
 sg13g2_fill_1 FILLER_138_380 ();
 sg13g2_fill_2 FILLER_138_426 ();
 sg13g2_fill_2 FILLER_138_443 ();
 sg13g2_fill_1 FILLER_138_445 ();
 sg13g2_decap_8 FILLER_138_451 ();
 sg13g2_decap_4 FILLER_138_458 ();
 sg13g2_fill_2 FILLER_138_462 ();
 sg13g2_decap_4 FILLER_138_479 ();
 sg13g2_fill_2 FILLER_138_483 ();
 sg13g2_fill_1 FILLER_138_495 ();
 sg13g2_decap_8 FILLER_138_506 ();
 sg13g2_decap_8 FILLER_138_513 ();
 sg13g2_decap_8 FILLER_138_520 ();
 sg13g2_decap_8 FILLER_138_527 ();
 sg13g2_decap_8 FILLER_138_534 ();
 sg13g2_decap_8 FILLER_138_541 ();
 sg13g2_decap_8 FILLER_138_563 ();
 sg13g2_decap_8 FILLER_138_570 ();
 sg13g2_decap_4 FILLER_138_577 ();
 sg13g2_decap_4 FILLER_138_586 ();
 sg13g2_fill_1 FILLER_138_590 ();
 sg13g2_fill_2 FILLER_138_600 ();
 sg13g2_fill_1 FILLER_138_635 ();
 sg13g2_fill_2 FILLER_138_668 ();
 sg13g2_fill_1 FILLER_138_670 ();
 sg13g2_decap_4 FILLER_138_691 ();
 sg13g2_fill_1 FILLER_138_695 ();
 sg13g2_decap_8 FILLER_138_754 ();
 sg13g2_decap_4 FILLER_138_761 ();
 sg13g2_fill_1 FILLER_138_765 ();
 sg13g2_decap_8 FILLER_138_785 ();
 sg13g2_decap_8 FILLER_138_792 ();
 sg13g2_decap_8 FILLER_138_799 ();
 sg13g2_decap_8 FILLER_138_816 ();
 sg13g2_decap_4 FILLER_138_823 ();
 sg13g2_fill_1 FILLER_138_827 ();
 sg13g2_fill_2 FILLER_138_854 ();
 sg13g2_fill_2 FILLER_138_874 ();
 sg13g2_fill_1 FILLER_138_876 ();
 sg13g2_fill_2 FILLER_138_884 ();
 sg13g2_decap_8 FILLER_138_896 ();
 sg13g2_decap_8 FILLER_138_903 ();
 sg13g2_decap_8 FILLER_138_914 ();
 sg13g2_decap_8 FILLER_138_921 ();
 sg13g2_decap_8 FILLER_138_928 ();
 sg13g2_fill_2 FILLER_138_935 ();
 sg13g2_fill_1 FILLER_138_937 ();
 sg13g2_decap_8 FILLER_138_943 ();
 sg13g2_fill_2 FILLER_138_954 ();
 sg13g2_fill_2 FILLER_138_990 ();
 sg13g2_decap_8 FILLER_138_1018 ();
 sg13g2_decap_4 FILLER_138_1025 ();
 sg13g2_fill_2 FILLER_138_1029 ();
 sg13g2_fill_2 FILLER_138_1088 ();
 sg13g2_fill_1 FILLER_138_1090 ();
 sg13g2_decap_8 FILLER_138_1117 ();
 sg13g2_fill_1 FILLER_138_1124 ();
 sg13g2_decap_8 FILLER_138_1142 ();
 sg13g2_decap_4 FILLER_138_1149 ();
 sg13g2_fill_2 FILLER_138_1153 ();
 sg13g2_decap_8 FILLER_138_1161 ();
 sg13g2_decap_8 FILLER_138_1168 ();
 sg13g2_decap_8 FILLER_138_1175 ();
 sg13g2_fill_1 FILLER_138_1186 ();
 sg13g2_decap_8 FILLER_138_1191 ();
 sg13g2_decap_8 FILLER_138_1203 ();
 sg13g2_decap_8 FILLER_138_1214 ();
 sg13g2_fill_2 FILLER_138_1221 ();
 sg13g2_decap_4 FILLER_138_1249 ();
 sg13g2_fill_1 FILLER_138_1282 ();
 sg13g2_decap_8 FILLER_138_1287 ();
 sg13g2_decap_8 FILLER_138_1323 ();
 sg13g2_decap_8 FILLER_138_1330 ();
 sg13g2_decap_8 FILLER_138_1337 ();
 sg13g2_decap_8 FILLER_138_1344 ();
 sg13g2_decap_8 FILLER_138_1351 ();
 sg13g2_decap_8 FILLER_138_1358 ();
 sg13g2_decap_8 FILLER_138_1365 ();
 sg13g2_decap_8 FILLER_138_1372 ();
 sg13g2_decap_8 FILLER_138_1379 ();
 sg13g2_decap_8 FILLER_138_1386 ();
 sg13g2_decap_8 FILLER_138_1393 ();
 sg13g2_decap_8 FILLER_138_1400 ();
 sg13g2_decap_8 FILLER_138_1407 ();
 sg13g2_decap_8 FILLER_138_1414 ();
 sg13g2_decap_8 FILLER_138_1421 ();
 sg13g2_decap_8 FILLER_138_1428 ();
 sg13g2_decap_8 FILLER_138_1435 ();
 sg13g2_decap_8 FILLER_138_1442 ();
 sg13g2_decap_8 FILLER_138_1449 ();
 sg13g2_decap_8 FILLER_138_1456 ();
 sg13g2_decap_8 FILLER_138_1463 ();
 sg13g2_decap_8 FILLER_138_1470 ();
 sg13g2_decap_8 FILLER_138_1477 ();
 sg13g2_decap_8 FILLER_138_1484 ();
 sg13g2_decap_8 FILLER_138_1491 ();
 sg13g2_decap_8 FILLER_138_1498 ();
 sg13g2_decap_8 FILLER_138_1505 ();
 sg13g2_decap_8 FILLER_138_1512 ();
 sg13g2_decap_8 FILLER_138_1519 ();
 sg13g2_decap_8 FILLER_138_1526 ();
 sg13g2_decap_8 FILLER_138_1533 ();
 sg13g2_decap_8 FILLER_138_1540 ();
 sg13g2_decap_8 FILLER_138_1547 ();
 sg13g2_decap_8 FILLER_138_1554 ();
 sg13g2_decap_8 FILLER_138_1561 ();
 sg13g2_decap_8 FILLER_138_1568 ();
 sg13g2_decap_8 FILLER_138_1575 ();
 sg13g2_decap_8 FILLER_138_1582 ();
 sg13g2_decap_8 FILLER_138_1589 ();
 sg13g2_decap_8 FILLER_138_1596 ();
 sg13g2_decap_8 FILLER_138_1603 ();
 sg13g2_decap_8 FILLER_138_1610 ();
 sg13g2_decap_8 FILLER_138_1617 ();
 sg13g2_fill_1 FILLER_138_1624 ();
 sg13g2_decap_8 FILLER_139_0 ();
 sg13g2_decap_4 FILLER_139_7 ();
 sg13g2_decap_8 FILLER_139_19 ();
 sg13g2_decap_8 FILLER_139_26 ();
 sg13g2_decap_8 FILLER_139_33 ();
 sg13g2_decap_4 FILLER_139_44 ();
 sg13g2_fill_1 FILLER_139_48 ();
 sg13g2_decap_8 FILLER_139_53 ();
 sg13g2_fill_1 FILLER_139_64 ();
 sg13g2_fill_1 FILLER_139_70 ();
 sg13g2_fill_1 FILLER_139_79 ();
 sg13g2_fill_1 FILLER_139_86 ();
 sg13g2_decap_8 FILLER_139_91 ();
 sg13g2_decap_8 FILLER_139_98 ();
 sg13g2_decap_8 FILLER_139_105 ();
 sg13g2_decap_8 FILLER_139_112 ();
 sg13g2_decap_8 FILLER_139_119 ();
 sg13g2_fill_2 FILLER_139_126 ();
 sg13g2_decap_8 FILLER_139_132 ();
 sg13g2_fill_1 FILLER_139_139 ();
 sg13g2_decap_8 FILLER_139_171 ();
 sg13g2_decap_8 FILLER_139_178 ();
 sg13g2_fill_2 FILLER_139_185 ();
 sg13g2_fill_1 FILLER_139_187 ();
 sg13g2_decap_8 FILLER_139_193 ();
 sg13g2_fill_1 FILLER_139_200 ();
 sg13g2_decap_8 FILLER_139_205 ();
 sg13g2_decap_8 FILLER_139_212 ();
 sg13g2_decap_8 FILLER_139_219 ();
 sg13g2_decap_8 FILLER_139_226 ();
 sg13g2_fill_2 FILLER_139_233 ();
 sg13g2_decap_8 FILLER_139_239 ();
 sg13g2_decap_8 FILLER_139_246 ();
 sg13g2_decap_8 FILLER_139_253 ();
 sg13g2_decap_8 FILLER_139_260 ();
 sg13g2_decap_8 FILLER_139_267 ();
 sg13g2_fill_2 FILLER_139_274 ();
 sg13g2_decap_4 FILLER_139_284 ();
 sg13g2_fill_2 FILLER_139_293 ();
 sg13g2_decap_4 FILLER_139_301 ();
 sg13g2_fill_2 FILLER_139_317 ();
 sg13g2_fill_1 FILLER_139_319 ();
 sg13g2_decap_4 FILLER_139_330 ();
 sg13g2_decap_8 FILLER_139_369 ();
 sg13g2_decap_8 FILLER_139_376 ();
 sg13g2_decap_8 FILLER_139_383 ();
 sg13g2_fill_2 FILLER_139_390 ();
 sg13g2_decap_8 FILLER_139_396 ();
 sg13g2_fill_2 FILLER_139_408 ();
 sg13g2_fill_1 FILLER_139_410 ();
 sg13g2_decap_8 FILLER_139_420 ();
 sg13g2_decap_4 FILLER_139_427 ();
 sg13g2_decap_8 FILLER_139_457 ();
 sg13g2_decap_4 FILLER_139_464 ();
 sg13g2_fill_2 FILLER_139_468 ();
 sg13g2_decap_4 FILLER_139_481 ();
 sg13g2_decap_8 FILLER_139_491 ();
 sg13g2_decap_4 FILLER_139_498 ();
 sg13g2_fill_2 FILLER_139_502 ();
 sg13g2_decap_8 FILLER_139_521 ();
 sg13g2_decap_8 FILLER_139_528 ();
 sg13g2_decap_4 FILLER_139_535 ();
 sg13g2_fill_1 FILLER_139_539 ();
 sg13g2_decap_8 FILLER_139_544 ();
 sg13g2_decap_4 FILLER_139_551 ();
 sg13g2_fill_1 FILLER_139_555 ();
 sg13g2_decap_4 FILLER_139_571 ();
 sg13g2_fill_2 FILLER_139_575 ();
 sg13g2_fill_1 FILLER_139_581 ();
 sg13g2_decap_4 FILLER_139_596 ();
 sg13g2_fill_2 FILLER_139_600 ();
 sg13g2_fill_1 FILLER_139_653 ();
 sg13g2_fill_2 FILLER_139_683 ();
 sg13g2_fill_1 FILLER_139_685 ();
 sg13g2_decap_8 FILLER_139_691 ();
 sg13g2_decap_8 FILLER_139_698 ();
 sg13g2_decap_4 FILLER_139_705 ();
 sg13g2_fill_2 FILLER_139_709 ();
 sg13g2_decap_8 FILLER_139_715 ();
 sg13g2_fill_2 FILLER_139_727 ();
 sg13g2_fill_1 FILLER_139_729 ();
 sg13g2_decap_8 FILLER_139_750 ();
 sg13g2_decap_8 FILLER_139_757 ();
 sg13g2_fill_2 FILLER_139_764 ();
 sg13g2_fill_1 FILLER_139_766 ();
 sg13g2_decap_8 FILLER_139_777 ();
 sg13g2_decap_8 FILLER_139_784 ();
 sg13g2_decap_8 FILLER_139_791 ();
 sg13g2_fill_1 FILLER_139_803 ();
 sg13g2_fill_2 FILLER_139_812 ();
 sg13g2_fill_1 FILLER_139_814 ();
 sg13g2_decap_8 FILLER_139_819 ();
 sg13g2_decap_4 FILLER_139_831 ();
 sg13g2_decap_8 FILLER_139_857 ();
 sg13g2_decap_8 FILLER_139_864 ();
 sg13g2_decap_4 FILLER_139_871 ();
 sg13g2_fill_2 FILLER_139_875 ();
 sg13g2_fill_1 FILLER_139_882 ();
 sg13g2_fill_2 FILLER_139_902 ();
 sg13g2_decap_4 FILLER_139_922 ();
 sg13g2_fill_2 FILLER_139_932 ();
 sg13g2_fill_1 FILLER_139_939 ();
 sg13g2_fill_1 FILLER_139_946 ();
 sg13g2_fill_1 FILLER_139_951 ();
 sg13g2_fill_1 FILLER_139_957 ();
 sg13g2_fill_1 FILLER_139_989 ();
 sg13g2_fill_2 FILLER_139_995 ();
 sg13g2_fill_1 FILLER_139_997 ();
 sg13g2_decap_8 FILLER_139_1003 ();
 sg13g2_fill_1 FILLER_139_1010 ();
 sg13g2_decap_4 FILLER_139_1017 ();
 sg13g2_fill_2 FILLER_139_1021 ();
 sg13g2_decap_8 FILLER_139_1056 ();
 sg13g2_decap_8 FILLER_139_1063 ();
 sg13g2_decap_8 FILLER_139_1074 ();
 sg13g2_fill_2 FILLER_139_1081 ();
 sg13g2_fill_1 FILLER_139_1083 ();
 sg13g2_fill_1 FILLER_139_1115 ();
 sg13g2_decap_8 FILLER_139_1128 ();
 sg13g2_decap_4 FILLER_139_1135 ();
 sg13g2_fill_2 FILLER_139_1146 ();
 sg13g2_fill_1 FILLER_139_1148 ();
 sg13g2_fill_2 FILLER_139_1154 ();
 sg13g2_decap_8 FILLER_139_1160 ();
 sg13g2_fill_2 FILLER_139_1167 ();
 sg13g2_fill_1 FILLER_139_1169 ();
 sg13g2_decap_4 FILLER_139_1205 ();
 sg13g2_fill_1 FILLER_139_1213 ();
 sg13g2_fill_2 FILLER_139_1244 ();
 sg13g2_decap_8 FILLER_139_1277 ();
 sg13g2_decap_8 FILLER_139_1284 ();
 sg13g2_decap_8 FILLER_139_1291 ();
 sg13g2_decap_8 FILLER_139_1298 ();
 sg13g2_decap_8 FILLER_139_1305 ();
 sg13g2_decap_8 FILLER_139_1312 ();
 sg13g2_decap_8 FILLER_139_1319 ();
 sg13g2_decap_8 FILLER_139_1326 ();
 sg13g2_decap_8 FILLER_139_1333 ();
 sg13g2_decap_8 FILLER_139_1340 ();
 sg13g2_decap_8 FILLER_139_1347 ();
 sg13g2_decap_8 FILLER_139_1354 ();
 sg13g2_decap_8 FILLER_139_1361 ();
 sg13g2_decap_8 FILLER_139_1368 ();
 sg13g2_decap_8 FILLER_139_1375 ();
 sg13g2_decap_8 FILLER_139_1382 ();
 sg13g2_decap_8 FILLER_139_1389 ();
 sg13g2_decap_8 FILLER_139_1396 ();
 sg13g2_decap_8 FILLER_139_1403 ();
 sg13g2_decap_8 FILLER_139_1410 ();
 sg13g2_decap_8 FILLER_139_1417 ();
 sg13g2_decap_8 FILLER_139_1424 ();
 sg13g2_decap_8 FILLER_139_1431 ();
 sg13g2_decap_8 FILLER_139_1438 ();
 sg13g2_decap_8 FILLER_139_1445 ();
 sg13g2_decap_8 FILLER_139_1452 ();
 sg13g2_decap_8 FILLER_139_1459 ();
 sg13g2_decap_8 FILLER_139_1466 ();
 sg13g2_decap_8 FILLER_139_1473 ();
 sg13g2_decap_8 FILLER_139_1480 ();
 sg13g2_decap_8 FILLER_139_1487 ();
 sg13g2_decap_8 FILLER_139_1494 ();
 sg13g2_decap_8 FILLER_139_1501 ();
 sg13g2_decap_8 FILLER_139_1508 ();
 sg13g2_decap_8 FILLER_139_1515 ();
 sg13g2_decap_8 FILLER_139_1522 ();
 sg13g2_decap_8 FILLER_139_1529 ();
 sg13g2_decap_8 FILLER_139_1536 ();
 sg13g2_decap_8 FILLER_139_1543 ();
 sg13g2_decap_8 FILLER_139_1550 ();
 sg13g2_decap_8 FILLER_139_1557 ();
 sg13g2_decap_8 FILLER_139_1564 ();
 sg13g2_decap_8 FILLER_139_1571 ();
 sg13g2_decap_8 FILLER_139_1578 ();
 sg13g2_decap_8 FILLER_139_1585 ();
 sg13g2_decap_8 FILLER_139_1592 ();
 sg13g2_decap_8 FILLER_139_1599 ();
 sg13g2_decap_8 FILLER_139_1606 ();
 sg13g2_decap_8 FILLER_139_1613 ();
 sg13g2_decap_4 FILLER_139_1620 ();
 sg13g2_fill_1 FILLER_139_1624 ();
 sg13g2_decap_4 FILLER_140_0 ();
 sg13g2_fill_1 FILLER_140_4 ();
 sg13g2_decap_8 FILLER_140_31 ();
 sg13g2_decap_8 FILLER_140_38 ();
 sg13g2_decap_8 FILLER_140_51 ();
 sg13g2_fill_2 FILLER_140_63 ();
 sg13g2_fill_1 FILLER_140_65 ();
 sg13g2_decap_8 FILLER_140_71 ();
 sg13g2_decap_8 FILLER_140_78 ();
 sg13g2_decap_4 FILLER_140_85 ();
 sg13g2_fill_1 FILLER_140_89 ();
 sg13g2_decap_8 FILLER_140_95 ();
 sg13g2_fill_1 FILLER_140_102 ();
 sg13g2_decap_8 FILLER_140_107 ();
 sg13g2_decap_8 FILLER_140_114 ();
 sg13g2_decap_4 FILLER_140_121 ();
 sg13g2_decap_8 FILLER_140_130 ();
 sg13g2_decap_8 FILLER_140_137 ();
 sg13g2_decap_8 FILLER_140_144 ();
 sg13g2_decap_8 FILLER_140_151 ();
 sg13g2_decap_8 FILLER_140_158 ();
 sg13g2_fill_1 FILLER_140_165 ();
 sg13g2_fill_1 FILLER_140_170 ();
 sg13g2_decap_4 FILLER_140_180 ();
 sg13g2_fill_1 FILLER_140_184 ();
 sg13g2_decap_8 FILLER_140_216 ();
 sg13g2_decap_4 FILLER_140_223 ();
 sg13g2_fill_1 FILLER_140_262 ();
 sg13g2_fill_2 FILLER_140_268 ();
 sg13g2_fill_1 FILLER_140_270 ();
 sg13g2_fill_2 FILLER_140_283 ();
 sg13g2_fill_1 FILLER_140_285 ();
 sg13g2_decap_4 FILLER_140_290 ();
 sg13g2_fill_1 FILLER_140_324 ();
 sg13g2_decap_4 FILLER_140_356 ();
 sg13g2_fill_2 FILLER_140_365 ();
 sg13g2_fill_1 FILLER_140_367 ();
 sg13g2_decap_8 FILLER_140_397 ();
 sg13g2_fill_2 FILLER_140_404 ();
 sg13g2_fill_1 FILLER_140_406 ();
 sg13g2_decap_4 FILLER_140_433 ();
 sg13g2_fill_1 FILLER_140_437 ();
 sg13g2_decap_8 FILLER_140_442 ();
 sg13g2_decap_8 FILLER_140_449 ();
 sg13g2_fill_1 FILLER_140_473 ();
 sg13g2_decap_4 FILLER_140_478 ();
 sg13g2_fill_1 FILLER_140_482 ();
 sg13g2_fill_2 FILLER_140_489 ();
 sg13g2_fill_2 FILLER_140_497 ();
 sg13g2_fill_1 FILLER_140_499 ();
 sg13g2_decap_8 FILLER_140_505 ();
 sg13g2_fill_1 FILLER_140_512 ();
 sg13g2_decap_8 FILLER_140_517 ();
 sg13g2_fill_2 FILLER_140_524 ();
 sg13g2_decap_8 FILLER_140_530 ();
 sg13g2_fill_2 FILLER_140_537 ();
 sg13g2_fill_1 FILLER_140_539 ();
 sg13g2_decap_8 FILLER_140_548 ();
 sg13g2_decap_8 FILLER_140_555 ();
 sg13g2_decap_4 FILLER_140_562 ();
 sg13g2_decap_4 FILLER_140_597 ();
 sg13g2_fill_2 FILLER_140_601 ();
 sg13g2_decap_4 FILLER_140_607 ();
 sg13g2_decap_4 FILLER_140_615 ();
 sg13g2_fill_1 FILLER_140_619 ();
 sg13g2_fill_2 FILLER_140_625 ();
 sg13g2_fill_1 FILLER_140_627 ();
 sg13g2_fill_1 FILLER_140_633 ();
 sg13g2_fill_1 FILLER_140_639 ();
 sg13g2_fill_2 FILLER_140_650 ();
 sg13g2_decap_4 FILLER_140_678 ();
 sg13g2_fill_2 FILLER_140_692 ();
 sg13g2_decap_4 FILLER_140_699 ();
 sg13g2_fill_1 FILLER_140_703 ();
 sg13g2_fill_2 FILLER_140_740 ();
 sg13g2_fill_2 FILLER_140_747 ();
 sg13g2_fill_1 FILLER_140_753 ();
 sg13g2_fill_2 FILLER_140_770 ();
 sg13g2_fill_2 FILLER_140_777 ();
 sg13g2_fill_2 FILLER_140_811 ();
 sg13g2_fill_1 FILLER_140_813 ();
 sg13g2_decap_8 FILLER_140_822 ();
 sg13g2_decap_4 FILLER_140_829 ();
 sg13g2_fill_2 FILLER_140_833 ();
 sg13g2_decap_8 FILLER_140_845 ();
 sg13g2_decap_8 FILLER_140_852 ();
 sg13g2_decap_4 FILLER_140_867 ();
 sg13g2_fill_1 FILLER_140_871 ();
 sg13g2_decap_8 FILLER_140_883 ();
 sg13g2_decap_8 FILLER_140_890 ();
 sg13g2_decap_4 FILLER_140_897 ();
 sg13g2_fill_1 FILLER_140_901 ();
 sg13g2_decap_4 FILLER_140_906 ();
 sg13g2_fill_2 FILLER_140_910 ();
 sg13g2_fill_1 FILLER_140_935 ();
 sg13g2_fill_2 FILLER_140_947 ();
 sg13g2_fill_1 FILLER_140_949 ();
 sg13g2_decap_8 FILLER_140_965 ();
 sg13g2_decap_8 FILLER_140_976 ();
 sg13g2_fill_2 FILLER_140_983 ();
 sg13g2_decap_8 FILLER_140_990 ();
 sg13g2_decap_8 FILLER_140_1001 ();
 sg13g2_decap_8 FILLER_140_1008 ();
 sg13g2_fill_2 FILLER_140_1023 ();
 sg13g2_fill_1 FILLER_140_1025 ();
 sg13g2_fill_2 FILLER_140_1067 ();
 sg13g2_fill_1 FILLER_140_1069 ();
 sg13g2_decap_8 FILLER_140_1074 ();
 sg13g2_decap_8 FILLER_140_1081 ();
 sg13g2_fill_1 FILLER_140_1088 ();
 sg13g2_fill_2 FILLER_140_1099 ();
 sg13g2_fill_1 FILLER_140_1107 ();
 sg13g2_decap_8 FILLER_140_1126 ();
 sg13g2_decap_8 FILLER_140_1137 ();
 sg13g2_decap_4 FILLER_140_1144 ();
 sg13g2_fill_1 FILLER_140_1174 ();
 sg13g2_decap_4 FILLER_140_1253 ();
 sg13g2_fill_2 FILLER_140_1257 ();
 sg13g2_decap_4 FILLER_140_1263 ();
 sg13g2_fill_1 FILLER_140_1267 ();
 sg13g2_decap_4 FILLER_140_1273 ();
 sg13g2_decap_8 FILLER_140_1281 ();
 sg13g2_decap_8 FILLER_140_1288 ();
 sg13g2_decap_8 FILLER_140_1295 ();
 sg13g2_decap_8 FILLER_140_1302 ();
 sg13g2_decap_8 FILLER_140_1309 ();
 sg13g2_decap_8 FILLER_140_1316 ();
 sg13g2_decap_8 FILLER_140_1323 ();
 sg13g2_decap_8 FILLER_140_1330 ();
 sg13g2_decap_8 FILLER_140_1337 ();
 sg13g2_decap_8 FILLER_140_1344 ();
 sg13g2_decap_8 FILLER_140_1351 ();
 sg13g2_decap_8 FILLER_140_1358 ();
 sg13g2_decap_8 FILLER_140_1365 ();
 sg13g2_decap_8 FILLER_140_1372 ();
 sg13g2_decap_8 FILLER_140_1379 ();
 sg13g2_decap_8 FILLER_140_1386 ();
 sg13g2_decap_8 FILLER_140_1393 ();
 sg13g2_decap_8 FILLER_140_1400 ();
 sg13g2_decap_8 FILLER_140_1407 ();
 sg13g2_decap_8 FILLER_140_1414 ();
 sg13g2_decap_8 FILLER_140_1421 ();
 sg13g2_decap_8 FILLER_140_1428 ();
 sg13g2_decap_8 FILLER_140_1435 ();
 sg13g2_decap_8 FILLER_140_1442 ();
 sg13g2_decap_8 FILLER_140_1449 ();
 sg13g2_decap_8 FILLER_140_1456 ();
 sg13g2_decap_8 FILLER_140_1463 ();
 sg13g2_decap_8 FILLER_140_1470 ();
 sg13g2_decap_8 FILLER_140_1477 ();
 sg13g2_decap_8 FILLER_140_1484 ();
 sg13g2_decap_8 FILLER_140_1491 ();
 sg13g2_decap_8 FILLER_140_1498 ();
 sg13g2_decap_8 FILLER_140_1505 ();
 sg13g2_decap_8 FILLER_140_1512 ();
 sg13g2_decap_8 FILLER_140_1519 ();
 sg13g2_decap_8 FILLER_140_1526 ();
 sg13g2_decap_8 FILLER_140_1533 ();
 sg13g2_decap_8 FILLER_140_1540 ();
 sg13g2_decap_8 FILLER_140_1547 ();
 sg13g2_decap_8 FILLER_140_1554 ();
 sg13g2_decap_8 FILLER_140_1561 ();
 sg13g2_decap_8 FILLER_140_1568 ();
 sg13g2_decap_8 FILLER_140_1575 ();
 sg13g2_decap_8 FILLER_140_1582 ();
 sg13g2_decap_8 FILLER_140_1589 ();
 sg13g2_decap_8 FILLER_140_1596 ();
 sg13g2_decap_8 FILLER_140_1603 ();
 sg13g2_decap_8 FILLER_140_1610 ();
 sg13g2_decap_8 FILLER_140_1617 ();
 sg13g2_fill_1 FILLER_140_1624 ();
 sg13g2_decap_8 FILLER_141_0 ();
 sg13g2_fill_2 FILLER_141_17 ();
 sg13g2_fill_1 FILLER_141_19 ();
 sg13g2_fill_1 FILLER_141_23 ();
 sg13g2_decap_4 FILLER_141_45 ();
 sg13g2_fill_1 FILLER_141_49 ();
 sg13g2_decap_4 FILLER_141_55 ();
 sg13g2_fill_1 FILLER_141_59 ();
 sg13g2_fill_1 FILLER_141_69 ();
 sg13g2_decap_8 FILLER_141_78 ();
 sg13g2_fill_2 FILLER_141_85 ();
 sg13g2_fill_1 FILLER_141_87 ();
 sg13g2_fill_2 FILLER_141_190 ();
 sg13g2_fill_2 FILLER_141_196 ();
 sg13g2_fill_1 FILLER_141_198 ();
 sg13g2_fill_1 FILLER_141_221 ();
 sg13g2_decap_8 FILLER_141_238 ();
 sg13g2_fill_2 FILLER_141_245 ();
 sg13g2_fill_1 FILLER_141_247 ();
 sg13g2_fill_1 FILLER_141_253 ();
 sg13g2_fill_1 FILLER_141_259 ();
 sg13g2_decap_4 FILLER_141_266 ();
 sg13g2_decap_4 FILLER_141_275 ();
 sg13g2_fill_2 FILLER_141_305 ();
 sg13g2_fill_1 FILLER_141_307 ();
 sg13g2_decap_4 FILLER_141_358 ();
 sg13g2_decap_8 FILLER_141_394 ();
 sg13g2_decap_4 FILLER_141_401 ();
 sg13g2_fill_1 FILLER_141_405 ();
 sg13g2_decap_8 FILLER_141_411 ();
 sg13g2_decap_4 FILLER_141_418 ();
 sg13g2_decap_8 FILLER_141_425 ();
 sg13g2_decap_8 FILLER_141_432 ();
 sg13g2_decap_8 FILLER_141_439 ();
 sg13g2_fill_1 FILLER_141_446 ();
 sg13g2_decap_8 FILLER_141_451 ();
 sg13g2_fill_2 FILLER_141_458 ();
 sg13g2_decap_8 FILLER_141_467 ();
 sg13g2_decap_8 FILLER_141_474 ();
 sg13g2_decap_4 FILLER_141_486 ();
 sg13g2_fill_1 FILLER_141_490 ();
 sg13g2_fill_2 FILLER_141_501 ();
 sg13g2_decap_8 FILLER_141_544 ();
 sg13g2_fill_2 FILLER_141_551 ();
 sg13g2_fill_1 FILLER_141_561 ();
 sg13g2_decap_8 FILLER_141_565 ();
 sg13g2_decap_8 FILLER_141_572 ();
 sg13g2_decap_8 FILLER_141_579 ();
 sg13g2_decap_4 FILLER_141_586 ();
 sg13g2_decap_8 FILLER_141_597 ();
 sg13g2_decap_8 FILLER_141_604 ();
 sg13g2_decap_8 FILLER_141_611 ();
 sg13g2_decap_8 FILLER_141_618 ();
 sg13g2_fill_1 FILLER_141_629 ();
 sg13g2_fill_2 FILLER_141_655 ();
 sg13g2_fill_1 FILLER_141_657 ();
 sg13g2_fill_2 FILLER_141_661 ();
 sg13g2_decap_8 FILLER_141_667 ();
 sg13g2_decap_8 FILLER_141_674 ();
 sg13g2_fill_2 FILLER_141_681 ();
 sg13g2_fill_1 FILLER_141_683 ();
 sg13g2_decap_4 FILLER_141_689 ();
 sg13g2_decap_4 FILLER_141_699 ();
 sg13g2_fill_1 FILLER_141_708 ();
 sg13g2_fill_1 FILLER_141_719 ();
 sg13g2_fill_2 FILLER_141_761 ();
 sg13g2_fill_1 FILLER_141_763 ();
 sg13g2_decap_4 FILLER_141_769 ();
 sg13g2_decap_4 FILLER_141_778 ();
 sg13g2_fill_1 FILLER_141_782 ();
 sg13g2_decap_8 FILLER_141_793 ();
 sg13g2_decap_8 FILLER_141_805 ();
 sg13g2_decap_8 FILLER_141_812 ();
 sg13g2_fill_2 FILLER_141_819 ();
 sg13g2_fill_1 FILLER_141_821 ();
 sg13g2_decap_8 FILLER_141_848 ();
 sg13g2_fill_1 FILLER_141_855 ();
 sg13g2_decap_8 FILLER_141_861 ();
 sg13g2_fill_2 FILLER_141_868 ();
 sg13g2_decap_8 FILLER_141_874 ();
 sg13g2_decap_8 FILLER_141_881 ();
 sg13g2_fill_1 FILLER_141_888 ();
 sg13g2_decap_8 FILLER_141_892 ();
 sg13g2_decap_4 FILLER_141_899 ();
 sg13g2_fill_1 FILLER_141_903 ();
 sg13g2_decap_4 FILLER_141_916 ();
 sg13g2_fill_2 FILLER_141_920 ();
 sg13g2_decap_4 FILLER_141_939 ();
 sg13g2_fill_1 FILLER_141_943 ();
 sg13g2_decap_8 FILLER_141_948 ();
 sg13g2_fill_1 FILLER_141_955 ();
 sg13g2_decap_8 FILLER_141_959 ();
 sg13g2_decap_8 FILLER_141_966 ();
 sg13g2_decap_8 FILLER_141_973 ();
 sg13g2_decap_8 FILLER_141_980 ();
 sg13g2_fill_2 FILLER_141_987 ();
 sg13g2_decap_4 FILLER_141_1015 ();
 sg13g2_fill_2 FILLER_141_1019 ();
 sg13g2_decap_8 FILLER_141_1027 ();
 sg13g2_fill_2 FILLER_141_1034 ();
 sg13g2_fill_1 FILLER_141_1036 ();
 sg13g2_fill_1 FILLER_141_1046 ();
 sg13g2_decap_8 FILLER_141_1052 ();
 sg13g2_fill_2 FILLER_141_1059 ();
 sg13g2_fill_2 FILLER_141_1087 ();
 sg13g2_decap_4 FILLER_141_1120 ();
 sg13g2_fill_2 FILLER_141_1150 ();
 sg13g2_fill_1 FILLER_141_1190 ();
 sg13g2_fill_2 FILLER_141_1216 ();
 sg13g2_fill_1 FILLER_141_1218 ();
 sg13g2_decap_8 FILLER_141_1222 ();
 sg13g2_decap_4 FILLER_141_1229 ();
 sg13g2_fill_1 FILLER_141_1233 ();
 sg13g2_decap_8 FILLER_141_1238 ();
 sg13g2_fill_2 FILLER_141_1245 ();
 sg13g2_decap_8 FILLER_141_1251 ();
 sg13g2_decap_8 FILLER_141_1258 ();
 sg13g2_decap_4 FILLER_141_1265 ();
 sg13g2_decap_8 FILLER_141_1295 ();
 sg13g2_decap_8 FILLER_141_1302 ();
 sg13g2_decap_8 FILLER_141_1309 ();
 sg13g2_decap_8 FILLER_141_1316 ();
 sg13g2_decap_8 FILLER_141_1323 ();
 sg13g2_decap_8 FILLER_141_1330 ();
 sg13g2_decap_8 FILLER_141_1337 ();
 sg13g2_decap_8 FILLER_141_1344 ();
 sg13g2_decap_8 FILLER_141_1351 ();
 sg13g2_decap_8 FILLER_141_1358 ();
 sg13g2_decap_8 FILLER_141_1365 ();
 sg13g2_decap_8 FILLER_141_1372 ();
 sg13g2_decap_8 FILLER_141_1379 ();
 sg13g2_decap_8 FILLER_141_1386 ();
 sg13g2_decap_8 FILLER_141_1393 ();
 sg13g2_decap_8 FILLER_141_1400 ();
 sg13g2_decap_8 FILLER_141_1407 ();
 sg13g2_decap_8 FILLER_141_1414 ();
 sg13g2_decap_8 FILLER_141_1421 ();
 sg13g2_decap_8 FILLER_141_1428 ();
 sg13g2_decap_8 FILLER_141_1435 ();
 sg13g2_decap_8 FILLER_141_1442 ();
 sg13g2_decap_8 FILLER_141_1449 ();
 sg13g2_decap_8 FILLER_141_1456 ();
 sg13g2_decap_8 FILLER_141_1463 ();
 sg13g2_decap_8 FILLER_141_1470 ();
 sg13g2_decap_8 FILLER_141_1477 ();
 sg13g2_decap_8 FILLER_141_1484 ();
 sg13g2_decap_8 FILLER_141_1491 ();
 sg13g2_decap_8 FILLER_141_1498 ();
 sg13g2_decap_8 FILLER_141_1505 ();
 sg13g2_decap_8 FILLER_141_1512 ();
 sg13g2_decap_8 FILLER_141_1519 ();
 sg13g2_decap_8 FILLER_141_1526 ();
 sg13g2_decap_8 FILLER_141_1533 ();
 sg13g2_decap_8 FILLER_141_1540 ();
 sg13g2_decap_8 FILLER_141_1547 ();
 sg13g2_decap_8 FILLER_141_1554 ();
 sg13g2_decap_8 FILLER_141_1561 ();
 sg13g2_decap_8 FILLER_141_1568 ();
 sg13g2_decap_8 FILLER_141_1575 ();
 sg13g2_decap_8 FILLER_141_1582 ();
 sg13g2_decap_8 FILLER_141_1589 ();
 sg13g2_decap_8 FILLER_141_1596 ();
 sg13g2_decap_8 FILLER_141_1603 ();
 sg13g2_decap_8 FILLER_141_1610 ();
 sg13g2_decap_8 FILLER_141_1617 ();
 sg13g2_fill_1 FILLER_141_1624 ();
 sg13g2_fill_2 FILLER_142_0 ();
 sg13g2_fill_1 FILLER_142_2 ();
 sg13g2_fill_1 FILLER_142_32 ();
 sg13g2_decap_8 FILLER_142_43 ();
 sg13g2_decap_8 FILLER_142_50 ();
 sg13g2_decap_4 FILLER_142_57 ();
 sg13g2_fill_1 FILLER_142_61 ();
 sg13g2_decap_8 FILLER_142_72 ();
 sg13g2_decap_8 FILLER_142_79 ();
 sg13g2_decap_4 FILLER_142_86 ();
 sg13g2_decap_8 FILLER_142_96 ();
 sg13g2_fill_1 FILLER_142_103 ();
 sg13g2_decap_8 FILLER_142_133 ();
 sg13g2_fill_2 FILLER_142_140 ();
 sg13g2_decap_4 FILLER_142_146 ();
 sg13g2_decap_4 FILLER_142_184 ();
 sg13g2_decap_4 FILLER_142_218 ();
 sg13g2_decap_8 FILLER_142_235 ();
 sg13g2_fill_2 FILLER_142_242 ();
 sg13g2_fill_1 FILLER_142_244 ();
 sg13g2_fill_2 FILLER_142_253 ();
 sg13g2_fill_1 FILLER_142_255 ();
 sg13g2_fill_2 FILLER_142_260 ();
 sg13g2_decap_8 FILLER_142_267 ();
 sg13g2_fill_2 FILLER_142_274 ();
 sg13g2_fill_1 FILLER_142_276 ();
 sg13g2_fill_2 FILLER_142_318 ();
 sg13g2_fill_2 FILLER_142_326 ();
 sg13g2_fill_2 FILLER_142_333 ();
 sg13g2_fill_2 FILLER_142_357 ();
 sg13g2_decap_8 FILLER_142_401 ();
 sg13g2_fill_1 FILLER_142_408 ();
 sg13g2_decap_8 FILLER_142_421 ();
 sg13g2_decap_4 FILLER_142_428 ();
 sg13g2_fill_2 FILLER_142_432 ();
 sg13g2_decap_8 FILLER_142_438 ();
 sg13g2_decap_8 FILLER_142_445 ();
 sg13g2_decap_4 FILLER_142_452 ();
 sg13g2_fill_1 FILLER_142_456 ();
 sg13g2_decap_4 FILLER_142_466 ();
 sg13g2_fill_1 FILLER_142_470 ();
 sg13g2_decap_4 FILLER_142_477 ();
 sg13g2_fill_1 FILLER_142_481 ();
 sg13g2_decap_8 FILLER_142_486 ();
 sg13g2_fill_2 FILLER_142_493 ();
 sg13g2_fill_1 FILLER_142_495 ();
 sg13g2_decap_4 FILLER_142_513 ();
 sg13g2_fill_2 FILLER_142_517 ();
 sg13g2_decap_4 FILLER_142_553 ();
 sg13g2_fill_2 FILLER_142_557 ();
 sg13g2_fill_1 FILLER_142_570 ();
 sg13g2_fill_1 FILLER_142_582 ();
 sg13g2_decap_4 FILLER_142_588 ();
 sg13g2_fill_1 FILLER_142_592 ();
 sg13g2_decap_8 FILLER_142_597 ();
 sg13g2_decap_4 FILLER_142_604 ();
 sg13g2_fill_1 FILLER_142_608 ();
 sg13g2_decap_4 FILLER_142_635 ();
 sg13g2_fill_2 FILLER_142_669 ();
 sg13g2_fill_1 FILLER_142_671 ();
 sg13g2_decap_8 FILLER_142_677 ();
 sg13g2_decap_4 FILLER_142_684 ();
 sg13g2_fill_1 FILLER_142_688 ();
 sg13g2_fill_1 FILLER_142_697 ();
 sg13g2_decap_8 FILLER_142_708 ();
 sg13g2_fill_1 FILLER_142_715 ();
 sg13g2_fill_2 FILLER_142_727 ();
 sg13g2_fill_1 FILLER_142_729 ();
 sg13g2_fill_2 FILLER_142_734 ();
 sg13g2_fill_2 FILLER_142_762 ();
 sg13g2_fill_1 FILLER_142_764 ();
 sg13g2_fill_2 FILLER_142_769 ();
 sg13g2_fill_2 FILLER_142_775 ();
 sg13g2_fill_2 FILLER_142_787 ();
 sg13g2_fill_1 FILLER_142_789 ();
 sg13g2_decap_8 FILLER_142_797 ();
 sg13g2_decap_8 FILLER_142_804 ();
 sg13g2_decap_4 FILLER_142_811 ();
 sg13g2_fill_1 FILLER_142_815 ();
 sg13g2_fill_2 FILLER_142_820 ();
 sg13g2_fill_2 FILLER_142_827 ();
 sg13g2_decap_4 FILLER_142_838 ();
 sg13g2_fill_2 FILLER_142_842 ();
 sg13g2_decap_8 FILLER_142_848 ();
 sg13g2_decap_8 FILLER_142_859 ();
 sg13g2_decap_8 FILLER_142_866 ();
 sg13g2_fill_2 FILLER_142_894 ();
 sg13g2_fill_1 FILLER_142_896 ();
 sg13g2_decap_8 FILLER_142_906 ();
 sg13g2_decap_8 FILLER_142_913 ();
 sg13g2_decap_4 FILLER_142_920 ();
 sg13g2_decap_4 FILLER_142_930 ();
 sg13g2_fill_1 FILLER_142_934 ();
 sg13g2_fill_2 FILLER_142_961 ();
 sg13g2_fill_2 FILLER_142_968 ();
 sg13g2_fill_1 FILLER_142_970 ();
 sg13g2_decap_8 FILLER_142_977 ();
 sg13g2_decap_8 FILLER_142_990 ();
 sg13g2_decap_8 FILLER_142_997 ();
 sg13g2_fill_1 FILLER_142_1004 ();
 sg13g2_decap_4 FILLER_142_1069 ();
 sg13g2_fill_2 FILLER_142_1172 ();
 sg13g2_fill_1 FILLER_142_1187 ();
 sg13g2_decap_8 FILLER_142_1196 ();
 sg13g2_fill_2 FILLER_142_1203 ();
 sg13g2_fill_1 FILLER_142_1205 ();
 sg13g2_decap_8 FILLER_142_1290 ();
 sg13g2_decap_8 FILLER_142_1297 ();
 sg13g2_decap_8 FILLER_142_1304 ();
 sg13g2_decap_8 FILLER_142_1311 ();
 sg13g2_decap_8 FILLER_142_1318 ();
 sg13g2_decap_8 FILLER_142_1325 ();
 sg13g2_decap_8 FILLER_142_1332 ();
 sg13g2_decap_8 FILLER_142_1339 ();
 sg13g2_decap_8 FILLER_142_1346 ();
 sg13g2_decap_8 FILLER_142_1353 ();
 sg13g2_decap_8 FILLER_142_1360 ();
 sg13g2_decap_8 FILLER_142_1367 ();
 sg13g2_decap_8 FILLER_142_1374 ();
 sg13g2_decap_8 FILLER_142_1381 ();
 sg13g2_decap_8 FILLER_142_1388 ();
 sg13g2_decap_8 FILLER_142_1395 ();
 sg13g2_decap_8 FILLER_142_1402 ();
 sg13g2_decap_8 FILLER_142_1409 ();
 sg13g2_decap_8 FILLER_142_1416 ();
 sg13g2_decap_8 FILLER_142_1423 ();
 sg13g2_decap_8 FILLER_142_1430 ();
 sg13g2_decap_8 FILLER_142_1437 ();
 sg13g2_decap_8 FILLER_142_1444 ();
 sg13g2_decap_8 FILLER_142_1451 ();
 sg13g2_decap_8 FILLER_142_1458 ();
 sg13g2_decap_8 FILLER_142_1465 ();
 sg13g2_decap_8 FILLER_142_1472 ();
 sg13g2_decap_8 FILLER_142_1479 ();
 sg13g2_decap_8 FILLER_142_1486 ();
 sg13g2_decap_8 FILLER_142_1493 ();
 sg13g2_decap_8 FILLER_142_1500 ();
 sg13g2_decap_8 FILLER_142_1507 ();
 sg13g2_decap_8 FILLER_142_1514 ();
 sg13g2_decap_8 FILLER_142_1521 ();
 sg13g2_decap_8 FILLER_142_1528 ();
 sg13g2_decap_8 FILLER_142_1535 ();
 sg13g2_decap_8 FILLER_142_1542 ();
 sg13g2_decap_8 FILLER_142_1549 ();
 sg13g2_decap_8 FILLER_142_1556 ();
 sg13g2_decap_8 FILLER_142_1563 ();
 sg13g2_decap_8 FILLER_142_1570 ();
 sg13g2_decap_8 FILLER_142_1577 ();
 sg13g2_decap_8 FILLER_142_1584 ();
 sg13g2_decap_8 FILLER_142_1591 ();
 sg13g2_decap_8 FILLER_142_1598 ();
 sg13g2_decap_8 FILLER_142_1605 ();
 sg13g2_decap_8 FILLER_142_1612 ();
 sg13g2_decap_4 FILLER_142_1619 ();
 sg13g2_fill_2 FILLER_142_1623 ();
 sg13g2_decap_8 FILLER_143_0 ();
 sg13g2_fill_2 FILLER_143_11 ();
 sg13g2_fill_1 FILLER_143_13 ();
 sg13g2_fill_2 FILLER_143_19 ();
 sg13g2_fill_2 FILLER_143_26 ();
 sg13g2_fill_1 FILLER_143_28 ();
 sg13g2_decap_8 FILLER_143_39 ();
 sg13g2_decap_8 FILLER_143_46 ();
 sg13g2_decap_8 FILLER_143_53 ();
 sg13g2_decap_8 FILLER_143_60 ();
 sg13g2_fill_2 FILLER_143_67 ();
 sg13g2_fill_1 FILLER_143_73 ();
 sg13g2_decap_8 FILLER_143_82 ();
 sg13g2_fill_1 FILLER_143_120 ();
 sg13g2_fill_1 FILLER_143_126 ();
 sg13g2_decap_4 FILLER_143_132 ();
 sg13g2_fill_2 FILLER_143_162 ();
 sg13g2_decap_8 FILLER_143_169 ();
 sg13g2_decap_8 FILLER_143_176 ();
 sg13g2_fill_2 FILLER_143_183 ();
 sg13g2_decap_8 FILLER_143_222 ();
 sg13g2_decap_4 FILLER_143_229 ();
 sg13g2_decap_8 FILLER_143_240 ();
 sg13g2_decap_8 FILLER_143_247 ();
 sg13g2_fill_1 FILLER_143_263 ();
 sg13g2_decap_8 FILLER_143_304 ();
 sg13g2_decap_4 FILLER_143_311 ();
 sg13g2_decap_8 FILLER_143_320 ();
 sg13g2_decap_8 FILLER_143_327 ();
 sg13g2_fill_1 FILLER_143_334 ();
 sg13g2_fill_1 FILLER_143_344 ();
 sg13g2_decap_4 FILLER_143_360 ();
 sg13g2_fill_1 FILLER_143_364 ();
 sg13g2_fill_2 FILLER_143_372 ();
 sg13g2_fill_2 FILLER_143_413 ();
 sg13g2_fill_2 FILLER_143_454 ();
 sg13g2_fill_2 FILLER_143_482 ();
 sg13g2_decap_8 FILLER_143_491 ();
 sg13g2_fill_2 FILLER_143_498 ();
 sg13g2_fill_1 FILLER_143_500 ();
 sg13g2_fill_2 FILLER_143_510 ();
 sg13g2_decap_8 FILLER_143_554 ();
 sg13g2_decap_8 FILLER_143_561 ();
 sg13g2_decap_8 FILLER_143_576 ();
 sg13g2_fill_1 FILLER_143_583 ();
 sg13g2_fill_1 FILLER_143_614 ();
 sg13g2_decap_8 FILLER_143_623 ();
 sg13g2_fill_1 FILLER_143_648 ();
 sg13g2_decap_8 FILLER_143_680 ();
 sg13g2_decap_8 FILLER_143_687 ();
 sg13g2_fill_2 FILLER_143_694 ();
 sg13g2_fill_2 FILLER_143_703 ();
 sg13g2_decap_8 FILLER_143_710 ();
 sg13g2_fill_2 FILLER_143_717 ();
 sg13g2_fill_1 FILLER_143_719 ();
 sg13g2_fill_1 FILLER_143_725 ();
 sg13g2_fill_2 FILLER_143_736 ();
 sg13g2_fill_1 FILLER_143_742 ();
 sg13g2_decap_8 FILLER_143_754 ();
 sg13g2_decap_8 FILLER_143_761 ();
 sg13g2_fill_2 FILLER_143_768 ();
 sg13g2_fill_1 FILLER_143_781 ();
 sg13g2_fill_2 FILLER_143_792 ();
 sg13g2_fill_2 FILLER_143_799 ();
 sg13g2_decap_8 FILLER_143_806 ();
 sg13g2_decap_8 FILLER_143_813 ();
 sg13g2_fill_2 FILLER_143_820 ();
 sg13g2_fill_1 FILLER_143_822 ();
 sg13g2_fill_2 FILLER_143_874 ();
 sg13g2_fill_1 FILLER_143_876 ();
 sg13g2_fill_2 FILLER_143_898 ();
 sg13g2_fill_1 FILLER_143_900 ();
 sg13g2_fill_2 FILLER_143_942 ();
 sg13g2_decap_8 FILLER_143_949 ();
 sg13g2_fill_1 FILLER_143_956 ();
 sg13g2_decap_8 FILLER_143_964 ();
 sg13g2_fill_2 FILLER_143_992 ();
 sg13g2_fill_1 FILLER_143_998 ();
 sg13g2_fill_1 FILLER_143_1034 ();
 sg13g2_fill_2 FILLER_143_1045 ();
 sg13g2_decap_8 FILLER_143_1130 ();
 sg13g2_decap_4 FILLER_143_1137 ();
 sg13g2_fill_2 FILLER_143_1141 ();
 sg13g2_fill_2 FILLER_143_1175 ();
 sg13g2_fill_1 FILLER_143_1177 ();
 sg13g2_fill_2 FILLER_143_1230 ();
 sg13g2_fill_1 FILLER_143_1232 ();
 sg13g2_decap_8 FILLER_143_1241 ();
 sg13g2_decap_8 FILLER_143_1248 ();
 sg13g2_decap_8 FILLER_143_1255 ();
 sg13g2_fill_2 FILLER_143_1262 ();
 sg13g2_fill_1 FILLER_143_1264 ();
 sg13g2_decap_4 FILLER_143_1273 ();
 sg13g2_fill_2 FILLER_143_1277 ();
 sg13g2_decap_8 FILLER_143_1283 ();
 sg13g2_fill_2 FILLER_143_1290 ();
 sg13g2_decap_8 FILLER_143_1296 ();
 sg13g2_decap_8 FILLER_143_1303 ();
 sg13g2_decap_8 FILLER_143_1310 ();
 sg13g2_decap_8 FILLER_143_1317 ();
 sg13g2_decap_8 FILLER_143_1324 ();
 sg13g2_decap_8 FILLER_143_1331 ();
 sg13g2_decap_8 FILLER_143_1338 ();
 sg13g2_decap_8 FILLER_143_1345 ();
 sg13g2_decap_8 FILLER_143_1352 ();
 sg13g2_decap_8 FILLER_143_1359 ();
 sg13g2_decap_8 FILLER_143_1366 ();
 sg13g2_decap_8 FILLER_143_1373 ();
 sg13g2_decap_8 FILLER_143_1380 ();
 sg13g2_decap_8 FILLER_143_1387 ();
 sg13g2_decap_8 FILLER_143_1394 ();
 sg13g2_decap_8 FILLER_143_1401 ();
 sg13g2_decap_8 FILLER_143_1408 ();
 sg13g2_decap_8 FILLER_143_1415 ();
 sg13g2_decap_8 FILLER_143_1422 ();
 sg13g2_decap_8 FILLER_143_1429 ();
 sg13g2_decap_8 FILLER_143_1436 ();
 sg13g2_decap_8 FILLER_143_1443 ();
 sg13g2_decap_8 FILLER_143_1450 ();
 sg13g2_decap_8 FILLER_143_1457 ();
 sg13g2_decap_8 FILLER_143_1464 ();
 sg13g2_decap_8 FILLER_143_1471 ();
 sg13g2_decap_8 FILLER_143_1478 ();
 sg13g2_decap_8 FILLER_143_1485 ();
 sg13g2_decap_8 FILLER_143_1492 ();
 sg13g2_decap_8 FILLER_143_1499 ();
 sg13g2_decap_8 FILLER_143_1506 ();
 sg13g2_decap_8 FILLER_143_1513 ();
 sg13g2_decap_8 FILLER_143_1520 ();
 sg13g2_decap_8 FILLER_143_1527 ();
 sg13g2_decap_8 FILLER_143_1534 ();
 sg13g2_decap_8 FILLER_143_1541 ();
 sg13g2_decap_8 FILLER_143_1548 ();
 sg13g2_decap_8 FILLER_143_1555 ();
 sg13g2_decap_8 FILLER_143_1562 ();
 sg13g2_decap_8 FILLER_143_1569 ();
 sg13g2_decap_8 FILLER_143_1576 ();
 sg13g2_decap_8 FILLER_143_1583 ();
 sg13g2_decap_8 FILLER_143_1590 ();
 sg13g2_decap_8 FILLER_143_1597 ();
 sg13g2_decap_8 FILLER_143_1604 ();
 sg13g2_decap_8 FILLER_143_1611 ();
 sg13g2_decap_8 FILLER_143_1618 ();
 sg13g2_fill_2 FILLER_144_35 ();
 sg13g2_fill_2 FILLER_144_47 ();
 sg13g2_fill_1 FILLER_144_49 ();
 sg13g2_fill_1 FILLER_144_68 ();
 sg13g2_decap_8 FILLER_144_79 ();
 sg13g2_fill_1 FILLER_144_95 ();
 sg13g2_decap_4 FILLER_144_100 ();
 sg13g2_fill_1 FILLER_144_108 ();
 sg13g2_fill_2 FILLER_144_119 ();
 sg13g2_fill_1 FILLER_144_121 ();
 sg13g2_fill_1 FILLER_144_147 ();
 sg13g2_decap_8 FILLER_144_157 ();
 sg13g2_fill_2 FILLER_144_164 ();
 sg13g2_decap_8 FILLER_144_170 ();
 sg13g2_decap_8 FILLER_144_177 ();
 sg13g2_decap_8 FILLER_144_184 ();
 sg13g2_decap_4 FILLER_144_191 ();
 sg13g2_fill_2 FILLER_144_195 ();
 sg13g2_fill_2 FILLER_144_201 ();
 sg13g2_fill_2 FILLER_144_208 ();
 sg13g2_decap_8 FILLER_144_215 ();
 sg13g2_fill_1 FILLER_144_241 ();
 sg13g2_decap_8 FILLER_144_312 ();
 sg13g2_fill_1 FILLER_144_319 ();
 sg13g2_fill_1 FILLER_144_346 ();
 sg13g2_fill_1 FILLER_144_352 ();
 sg13g2_fill_1 FILLER_144_358 ();
 sg13g2_fill_2 FILLER_144_364 ();
 sg13g2_decap_4 FILLER_144_373 ();
 sg13g2_fill_1 FILLER_144_377 ();
 sg13g2_decap_8 FILLER_144_383 ();
 sg13g2_decap_8 FILLER_144_390 ();
 sg13g2_fill_1 FILLER_144_397 ();
 sg13g2_decap_8 FILLER_144_402 ();
 sg13g2_fill_2 FILLER_144_421 ();
 sg13g2_decap_8 FILLER_144_433 ();
 sg13g2_decap_8 FILLER_144_440 ();
 sg13g2_decap_8 FILLER_144_472 ();
 sg13g2_decap_4 FILLER_144_479 ();
 sg13g2_decap_8 FILLER_144_492 ();
 sg13g2_decap_4 FILLER_144_526 ();
 sg13g2_fill_2 FILLER_144_530 ();
 sg13g2_fill_2 FILLER_144_537 ();
 sg13g2_decap_8 FILLER_144_544 ();
 sg13g2_fill_2 FILLER_144_556 ();
 sg13g2_fill_1 FILLER_144_563 ();
 sg13g2_decap_8 FILLER_144_581 ();
 sg13g2_decap_8 FILLER_144_588 ();
 sg13g2_fill_1 FILLER_144_595 ();
 sg13g2_fill_2 FILLER_144_650 ();
 sg13g2_fill_1 FILLER_144_658 ();
 sg13g2_fill_2 FILLER_144_663 ();
 sg13g2_fill_1 FILLER_144_665 ();
 sg13g2_decap_8 FILLER_144_670 ();
 sg13g2_decap_8 FILLER_144_677 ();
 sg13g2_decap_8 FILLER_144_684 ();
 sg13g2_decap_8 FILLER_144_691 ();
 sg13g2_decap_8 FILLER_144_698 ();
 sg13g2_decap_4 FILLER_144_705 ();
 sg13g2_fill_2 FILLER_144_709 ();
 sg13g2_fill_2 FILLER_144_716 ();
 sg13g2_fill_1 FILLER_144_718 ();
 sg13g2_fill_2 FILLER_144_729 ();
 sg13g2_fill_1 FILLER_144_731 ();
 sg13g2_decap_8 FILLER_144_737 ();
 sg13g2_fill_2 FILLER_144_744 ();
 sg13g2_fill_1 FILLER_144_746 ();
 sg13g2_decap_8 FILLER_144_751 ();
 sg13g2_decap_8 FILLER_144_758 ();
 sg13g2_decap_8 FILLER_144_765 ();
 sg13g2_decap_8 FILLER_144_772 ();
 sg13g2_fill_2 FILLER_144_779 ();
 sg13g2_decap_4 FILLER_144_786 ();
 sg13g2_fill_2 FILLER_144_790 ();
 sg13g2_decap_4 FILLER_144_805 ();
 sg13g2_decap_8 FILLER_144_813 ();
 sg13g2_decap_8 FILLER_144_820 ();
 sg13g2_decap_4 FILLER_144_830 ();
 sg13g2_decap_8 FILLER_144_889 ();
 sg13g2_decap_8 FILLER_144_896 ();
 sg13g2_fill_2 FILLER_144_903 ();
 sg13g2_decap_8 FILLER_144_915 ();
 sg13g2_decap_4 FILLER_144_922 ();
 sg13g2_fill_2 FILLER_144_926 ();
 sg13g2_fill_1 FILLER_144_933 ();
 sg13g2_decap_8 FILLER_144_946 ();
 sg13g2_decap_4 FILLER_144_953 ();
 sg13g2_fill_1 FILLER_144_963 ();
 sg13g2_fill_2 FILLER_144_970 ();
 sg13g2_fill_2 FILLER_144_976 ();
 sg13g2_decap_4 FILLER_144_983 ();
 sg13g2_decap_8 FILLER_144_1017 ();
 sg13g2_decap_8 FILLER_144_1024 ();
 sg13g2_decap_8 FILLER_144_1031 ();
 sg13g2_decap_8 FILLER_144_1038 ();
 sg13g2_fill_2 FILLER_144_1045 ();
 sg13g2_fill_1 FILLER_144_1106 ();
 sg13g2_fill_2 FILLER_144_1138 ();
 sg13g2_decap_8 FILLER_144_1144 ();
 sg13g2_fill_2 FILLER_144_1151 ();
 sg13g2_fill_2 FILLER_144_1183 ();
 sg13g2_fill_2 FILLER_144_1197 ();
 sg13g2_decap_4 FILLER_144_1205 ();
 sg13g2_fill_2 FILLER_144_1209 ();
 sg13g2_decap_4 FILLER_144_1215 ();
 sg13g2_decap_8 FILLER_144_1236 ();
 sg13g2_decap_8 FILLER_144_1243 ();
 sg13g2_decap_8 FILLER_144_1250 ();
 sg13g2_fill_1 FILLER_144_1257 ();
 sg13g2_fill_1 FILLER_144_1263 ();
 sg13g2_fill_1 FILLER_144_1267 ();
 sg13g2_fill_1 FILLER_144_1272 ();
 sg13g2_fill_2 FILLER_144_1281 ();
 sg13g2_fill_1 FILLER_144_1283 ();
 sg13g2_decap_8 FILLER_144_1310 ();
 sg13g2_decap_8 FILLER_144_1317 ();
 sg13g2_decap_8 FILLER_144_1324 ();
 sg13g2_decap_8 FILLER_144_1331 ();
 sg13g2_decap_8 FILLER_144_1338 ();
 sg13g2_decap_8 FILLER_144_1345 ();
 sg13g2_decap_8 FILLER_144_1352 ();
 sg13g2_decap_8 FILLER_144_1359 ();
 sg13g2_decap_8 FILLER_144_1366 ();
 sg13g2_decap_8 FILLER_144_1373 ();
 sg13g2_decap_8 FILLER_144_1380 ();
 sg13g2_decap_8 FILLER_144_1387 ();
 sg13g2_decap_8 FILLER_144_1394 ();
 sg13g2_decap_8 FILLER_144_1401 ();
 sg13g2_decap_8 FILLER_144_1408 ();
 sg13g2_decap_8 FILLER_144_1415 ();
 sg13g2_decap_8 FILLER_144_1422 ();
 sg13g2_decap_8 FILLER_144_1429 ();
 sg13g2_decap_8 FILLER_144_1436 ();
 sg13g2_decap_8 FILLER_144_1443 ();
 sg13g2_decap_8 FILLER_144_1450 ();
 sg13g2_decap_8 FILLER_144_1457 ();
 sg13g2_decap_8 FILLER_144_1464 ();
 sg13g2_decap_8 FILLER_144_1471 ();
 sg13g2_decap_8 FILLER_144_1478 ();
 sg13g2_decap_8 FILLER_144_1485 ();
 sg13g2_decap_8 FILLER_144_1492 ();
 sg13g2_decap_8 FILLER_144_1499 ();
 sg13g2_decap_8 FILLER_144_1506 ();
 sg13g2_decap_8 FILLER_144_1513 ();
 sg13g2_decap_8 FILLER_144_1520 ();
 sg13g2_decap_8 FILLER_144_1527 ();
 sg13g2_decap_8 FILLER_144_1534 ();
 sg13g2_decap_8 FILLER_144_1541 ();
 sg13g2_decap_8 FILLER_144_1548 ();
 sg13g2_decap_8 FILLER_144_1555 ();
 sg13g2_decap_8 FILLER_144_1562 ();
 sg13g2_decap_8 FILLER_144_1569 ();
 sg13g2_decap_8 FILLER_144_1576 ();
 sg13g2_decap_8 FILLER_144_1583 ();
 sg13g2_decap_8 FILLER_144_1590 ();
 sg13g2_decap_8 FILLER_144_1597 ();
 sg13g2_decap_8 FILLER_144_1604 ();
 sg13g2_decap_8 FILLER_144_1611 ();
 sg13g2_decap_8 FILLER_144_1618 ();
 sg13g2_decap_8 FILLER_145_0 ();
 sg13g2_fill_2 FILLER_145_7 ();
 sg13g2_fill_1 FILLER_145_9 ();
 sg13g2_decap_8 FILLER_145_17 ();
 sg13g2_decap_8 FILLER_145_24 ();
 sg13g2_decap_8 FILLER_145_40 ();
 sg13g2_decap_8 FILLER_145_47 ();
 sg13g2_decap_4 FILLER_145_54 ();
 sg13g2_fill_2 FILLER_145_58 ();
 sg13g2_decap_8 FILLER_145_70 ();
 sg13g2_fill_1 FILLER_145_77 ();
 sg13g2_decap_4 FILLER_145_87 ();
 sg13g2_fill_1 FILLER_145_91 ();
 sg13g2_fill_2 FILLER_145_127 ();
 sg13g2_fill_2 FILLER_145_184 ();
 sg13g2_fill_1 FILLER_145_186 ();
 sg13g2_decap_4 FILLER_145_196 ();
 sg13g2_fill_2 FILLER_145_200 ();
 sg13g2_decap_4 FILLER_145_215 ();
 sg13g2_fill_2 FILLER_145_226 ();
 sg13g2_fill_1 FILLER_145_233 ();
 sg13g2_decap_8 FILLER_145_243 ();
 sg13g2_decap_8 FILLER_145_250 ();
 sg13g2_decap_8 FILLER_145_257 ();
 sg13g2_decap_4 FILLER_145_264 ();
 sg13g2_fill_1 FILLER_145_293 ();
 sg13g2_decap_8 FILLER_145_333 ();
 sg13g2_decap_8 FILLER_145_340 ();
 sg13g2_fill_1 FILLER_145_347 ();
 sg13g2_decap_4 FILLER_145_360 ();
 sg13g2_decap_8 FILLER_145_369 ();
 sg13g2_decap_4 FILLER_145_376 ();
 sg13g2_decap_8 FILLER_145_385 ();
 sg13g2_fill_1 FILLER_145_392 ();
 sg13g2_fill_1 FILLER_145_418 ();
 sg13g2_fill_2 FILLER_145_424 ();
 sg13g2_decap_8 FILLER_145_431 ();
 sg13g2_decap_8 FILLER_145_438 ();
 sg13g2_decap_8 FILLER_145_445 ();
 sg13g2_fill_2 FILLER_145_452 ();
 sg13g2_decap_4 FILLER_145_460 ();
 sg13g2_fill_1 FILLER_145_464 ();
 sg13g2_decap_4 FILLER_145_474 ();
 sg13g2_fill_1 FILLER_145_478 ();
 sg13g2_fill_2 FILLER_145_485 ();
 sg13g2_decap_8 FILLER_145_499 ();
 sg13g2_decap_8 FILLER_145_506 ();
 sg13g2_decap_8 FILLER_145_513 ();
 sg13g2_decap_8 FILLER_145_520 ();
 sg13g2_decap_8 FILLER_145_527 ();
 sg13g2_decap_8 FILLER_145_534 ();
 sg13g2_decap_8 FILLER_145_541 ();
 sg13g2_decap_8 FILLER_145_548 ();
 sg13g2_decap_8 FILLER_145_555 ();
 sg13g2_fill_1 FILLER_145_562 ();
 sg13g2_decap_8 FILLER_145_573 ();
 sg13g2_decap_4 FILLER_145_580 ();
 sg13g2_fill_1 FILLER_145_635 ();
 sg13g2_fill_2 FILLER_145_685 ();
 sg13g2_decap_8 FILLER_145_691 ();
 sg13g2_decap_8 FILLER_145_698 ();
 sg13g2_fill_2 FILLER_145_705 ();
 sg13g2_fill_2 FILLER_145_719 ();
 sg13g2_fill_1 FILLER_145_721 ();
 sg13g2_decap_8 FILLER_145_737 ();
 sg13g2_decap_8 FILLER_145_744 ();
 sg13g2_decap_8 FILLER_145_751 ();
 sg13g2_fill_2 FILLER_145_758 ();
 sg13g2_fill_1 FILLER_145_760 ();
 sg13g2_decap_8 FILLER_145_774 ();
 sg13g2_decap_8 FILLER_145_781 ();
 sg13g2_fill_2 FILLER_145_788 ();
 sg13g2_fill_1 FILLER_145_790 ();
 sg13g2_decap_8 FILLER_145_796 ();
 sg13g2_decap_4 FILLER_145_803 ();
 sg13g2_decap_8 FILLER_145_833 ();
 sg13g2_decap_8 FILLER_145_840 ();
 sg13g2_decap_8 FILLER_145_847 ();
 sg13g2_fill_1 FILLER_145_854 ();
 sg13g2_fill_2 FILLER_145_882 ();
 sg13g2_fill_2 FILLER_145_904 ();
 sg13g2_fill_1 FILLER_145_906 ();
 sg13g2_decap_8 FILLER_145_913 ();
 sg13g2_decap_8 FILLER_145_944 ();
 sg13g2_decap_8 FILLER_145_951 ();
 sg13g2_decap_8 FILLER_145_958 ();
 sg13g2_fill_1 FILLER_145_965 ();
 sg13g2_decap_8 FILLER_145_970 ();
 sg13g2_decap_8 FILLER_145_977 ();
 sg13g2_fill_2 FILLER_145_984 ();
 sg13g2_fill_1 FILLER_145_986 ();
 sg13g2_decap_8 FILLER_145_995 ();
 sg13g2_decap_8 FILLER_145_1002 ();
 sg13g2_decap_4 FILLER_145_1009 ();
 sg13g2_fill_1 FILLER_145_1013 ();
 sg13g2_fill_1 FILLER_145_1019 ();
 sg13g2_decap_4 FILLER_145_1024 ();
 sg13g2_fill_2 FILLER_145_1028 ();
 sg13g2_decap_4 FILLER_145_1034 ();
 sg13g2_fill_1 FILLER_145_1038 ();
 sg13g2_decap_4 FILLER_145_1044 ();
 sg13g2_fill_1 FILLER_145_1048 ();
 sg13g2_decap_4 FILLER_145_1055 ();
 sg13g2_fill_1 FILLER_145_1059 ();
 sg13g2_fill_2 FILLER_145_1065 ();
 sg13g2_fill_1 FILLER_145_1067 ();
 sg13g2_decap_8 FILLER_145_1072 ();
 sg13g2_fill_2 FILLER_145_1079 ();
 sg13g2_fill_1 FILLER_145_1081 ();
 sg13g2_fill_2 FILLER_145_1089 ();
 sg13g2_fill_1 FILLER_145_1091 ();
 sg13g2_decap_8 FILLER_145_1224 ();
 sg13g2_fill_2 FILLER_145_1242 ();
 sg13g2_decap_8 FILLER_145_1264 ();
 sg13g2_decap_8 FILLER_145_1316 ();
 sg13g2_decap_8 FILLER_145_1323 ();
 sg13g2_decap_8 FILLER_145_1330 ();
 sg13g2_decap_8 FILLER_145_1337 ();
 sg13g2_decap_8 FILLER_145_1344 ();
 sg13g2_decap_8 FILLER_145_1351 ();
 sg13g2_decap_8 FILLER_145_1358 ();
 sg13g2_decap_8 FILLER_145_1365 ();
 sg13g2_decap_8 FILLER_145_1372 ();
 sg13g2_decap_8 FILLER_145_1379 ();
 sg13g2_decap_8 FILLER_145_1386 ();
 sg13g2_decap_8 FILLER_145_1393 ();
 sg13g2_decap_8 FILLER_145_1400 ();
 sg13g2_decap_8 FILLER_145_1407 ();
 sg13g2_decap_8 FILLER_145_1414 ();
 sg13g2_decap_8 FILLER_145_1421 ();
 sg13g2_decap_8 FILLER_145_1428 ();
 sg13g2_decap_8 FILLER_145_1435 ();
 sg13g2_decap_8 FILLER_145_1442 ();
 sg13g2_decap_8 FILLER_145_1449 ();
 sg13g2_decap_8 FILLER_145_1456 ();
 sg13g2_decap_8 FILLER_145_1463 ();
 sg13g2_decap_8 FILLER_145_1470 ();
 sg13g2_decap_8 FILLER_145_1477 ();
 sg13g2_decap_8 FILLER_145_1484 ();
 sg13g2_decap_8 FILLER_145_1491 ();
 sg13g2_decap_8 FILLER_145_1498 ();
 sg13g2_decap_8 FILLER_145_1505 ();
 sg13g2_decap_8 FILLER_145_1512 ();
 sg13g2_decap_8 FILLER_145_1519 ();
 sg13g2_decap_8 FILLER_145_1526 ();
 sg13g2_decap_8 FILLER_145_1533 ();
 sg13g2_decap_8 FILLER_145_1540 ();
 sg13g2_decap_8 FILLER_145_1547 ();
 sg13g2_decap_8 FILLER_145_1554 ();
 sg13g2_decap_8 FILLER_145_1561 ();
 sg13g2_decap_8 FILLER_145_1568 ();
 sg13g2_decap_8 FILLER_145_1575 ();
 sg13g2_decap_8 FILLER_145_1582 ();
 sg13g2_decap_8 FILLER_145_1589 ();
 sg13g2_decap_8 FILLER_145_1596 ();
 sg13g2_decap_8 FILLER_145_1603 ();
 sg13g2_decap_8 FILLER_145_1610 ();
 sg13g2_decap_8 FILLER_145_1617 ();
 sg13g2_fill_1 FILLER_145_1624 ();
 sg13g2_decap_4 FILLER_146_0 ();
 sg13g2_decap_8 FILLER_146_11 ();
 sg13g2_decap_8 FILLER_146_18 ();
 sg13g2_decap_4 FILLER_146_25 ();
 sg13g2_decap_8 FILLER_146_48 ();
 sg13g2_decap_8 FILLER_146_55 ();
 sg13g2_decap_8 FILLER_146_70 ();
 sg13g2_decap_8 FILLER_146_77 ();
 sg13g2_decap_8 FILLER_146_115 ();
 sg13g2_decap_8 FILLER_146_122 ();
 sg13g2_fill_1 FILLER_146_129 ();
 sg13g2_decap_8 FILLER_146_160 ();
 sg13g2_decap_8 FILLER_146_171 ();
 sg13g2_fill_1 FILLER_146_178 ();
 sg13g2_fill_2 FILLER_146_208 ();
 sg13g2_decap_4 FILLER_146_236 ();
 sg13g2_decap_8 FILLER_146_266 ();
 sg13g2_fill_2 FILLER_146_273 ();
 sg13g2_decap_8 FILLER_146_279 ();
 sg13g2_fill_1 FILLER_146_292 ();
 sg13g2_decap_8 FILLER_146_298 ();
 sg13g2_fill_2 FILLER_146_305 ();
 sg13g2_decap_4 FILLER_146_337 ();
 sg13g2_fill_2 FILLER_146_341 ();
 sg13g2_decap_8 FILLER_146_347 ();
 sg13g2_fill_1 FILLER_146_354 ();
 sg13g2_decap_4 FILLER_146_373 ();
 sg13g2_decap_4 FILLER_146_416 ();
 sg13g2_fill_2 FILLER_146_420 ();
 sg13g2_decap_4 FILLER_146_430 ();
 sg13g2_fill_2 FILLER_146_434 ();
 sg13g2_decap_8 FILLER_146_440 ();
 sg13g2_fill_2 FILLER_146_447 ();
 sg13g2_fill_2 FILLER_146_456 ();
 sg13g2_fill_1 FILLER_146_458 ();
 sg13g2_fill_1 FILLER_146_491 ();
 sg13g2_fill_1 FILLER_146_496 ();
 sg13g2_fill_1 FILLER_146_505 ();
 sg13g2_fill_2 FILLER_146_512 ();
 sg13g2_fill_1 FILLER_146_514 ();
 sg13g2_decap_4 FILLER_146_521 ();
 sg13g2_fill_1 FILLER_146_525 ();
 sg13g2_fill_1 FILLER_146_531 ();
 sg13g2_decap_8 FILLER_146_538 ();
 sg13g2_decap_4 FILLER_146_564 ();
 sg13g2_fill_1 FILLER_146_568 ();
 sg13g2_decap_4 FILLER_146_587 ();
 sg13g2_fill_1 FILLER_146_591 ();
 sg13g2_fill_2 FILLER_146_618 ();
 sg13g2_fill_1 FILLER_146_620 ();
 sg13g2_decap_8 FILLER_146_660 ();
 sg13g2_decap_8 FILLER_146_667 ();
 sg13g2_decap_8 FILLER_146_674 ();
 sg13g2_decap_4 FILLER_146_707 ();
 sg13g2_fill_1 FILLER_146_726 ();
 sg13g2_decap_8 FILLER_146_744 ();
 sg13g2_fill_1 FILLER_146_791 ();
 sg13g2_decap_4 FILLER_146_801 ();
 sg13g2_fill_1 FILLER_146_805 ();
 sg13g2_decap_8 FILLER_146_816 ();
 sg13g2_decap_8 FILLER_146_823 ();
 sg13g2_decap_8 FILLER_146_830 ();
 sg13g2_fill_1 FILLER_146_837 ();
 sg13g2_fill_1 FILLER_146_848 ();
 sg13g2_fill_1 FILLER_146_858 ();
 sg13g2_fill_1 FILLER_146_865 ();
 sg13g2_fill_1 FILLER_146_870 ();
 sg13g2_decap_8 FILLER_146_879 ();
 sg13g2_fill_2 FILLER_146_886 ();
 sg13g2_fill_1 FILLER_146_888 ();
 sg13g2_decap_8 FILLER_146_894 ();
 sg13g2_decap_8 FILLER_146_901 ();
 sg13g2_decap_8 FILLER_146_914 ();
 sg13g2_fill_1 FILLER_146_921 ();
 sg13g2_decap_4 FILLER_146_927 ();
 sg13g2_decap_4 FILLER_146_935 ();
 sg13g2_decap_8 FILLER_146_944 ();
 sg13g2_decap_4 FILLER_146_951 ();
 sg13g2_decap_8 FILLER_146_962 ();
 sg13g2_decap_8 FILLER_146_975 ();
 sg13g2_decap_8 FILLER_146_982 ();
 sg13g2_fill_1 FILLER_146_989 ();
 sg13g2_fill_1 FILLER_146_995 ();
 sg13g2_decap_4 FILLER_146_1000 ();
 sg13g2_fill_1 FILLER_146_1004 ();
 sg13g2_fill_1 FILLER_146_1017 ();
 sg13g2_fill_1 FILLER_146_1049 ();
 sg13g2_decap_8 FILLER_146_1054 ();
 sg13g2_decap_8 FILLER_146_1061 ();
 sg13g2_fill_2 FILLER_146_1068 ();
 sg13g2_fill_1 FILLER_146_1070 ();
 sg13g2_decap_8 FILLER_146_1080 ();
 sg13g2_decap_4 FILLER_146_1087 ();
 sg13g2_fill_2 FILLER_146_1097 ();
 sg13g2_fill_2 FILLER_146_1105 ();
 sg13g2_fill_1 FILLER_146_1107 ();
 sg13g2_fill_1 FILLER_146_1111 ();
 sg13g2_fill_2 FILLER_146_1138 ();
 sg13g2_fill_1 FILLER_146_1140 ();
 sg13g2_decap_8 FILLER_146_1145 ();
 sg13g2_decap_4 FILLER_146_1152 ();
 sg13g2_fill_2 FILLER_146_1156 ();
 sg13g2_fill_2 FILLER_146_1193 ();
 sg13g2_fill_1 FILLER_146_1195 ();
 sg13g2_decap_8 FILLER_146_1206 ();
 sg13g2_decap_4 FILLER_146_1213 ();
 sg13g2_fill_1 FILLER_146_1217 ();
 sg13g2_decap_8 FILLER_146_1239 ();
 sg13g2_decap_8 FILLER_146_1246 ();
 sg13g2_fill_1 FILLER_146_1253 ();
 sg13g2_fill_2 FILLER_146_1265 ();
 sg13g2_decap_8 FILLER_146_1272 ();
 sg13g2_decap_8 FILLER_146_1279 ();
 sg13g2_fill_2 FILLER_146_1286 ();
 sg13g2_decap_8 FILLER_146_1314 ();
 sg13g2_decap_8 FILLER_146_1321 ();
 sg13g2_decap_8 FILLER_146_1328 ();
 sg13g2_decap_8 FILLER_146_1335 ();
 sg13g2_decap_8 FILLER_146_1342 ();
 sg13g2_decap_8 FILLER_146_1349 ();
 sg13g2_decap_8 FILLER_146_1356 ();
 sg13g2_decap_8 FILLER_146_1363 ();
 sg13g2_decap_8 FILLER_146_1370 ();
 sg13g2_decap_8 FILLER_146_1377 ();
 sg13g2_decap_8 FILLER_146_1384 ();
 sg13g2_decap_8 FILLER_146_1391 ();
 sg13g2_decap_8 FILLER_146_1398 ();
 sg13g2_decap_8 FILLER_146_1405 ();
 sg13g2_decap_8 FILLER_146_1412 ();
 sg13g2_decap_8 FILLER_146_1419 ();
 sg13g2_decap_8 FILLER_146_1426 ();
 sg13g2_decap_8 FILLER_146_1433 ();
 sg13g2_decap_8 FILLER_146_1440 ();
 sg13g2_decap_8 FILLER_146_1447 ();
 sg13g2_decap_8 FILLER_146_1454 ();
 sg13g2_decap_8 FILLER_146_1461 ();
 sg13g2_decap_8 FILLER_146_1468 ();
 sg13g2_decap_8 FILLER_146_1475 ();
 sg13g2_decap_8 FILLER_146_1482 ();
 sg13g2_decap_8 FILLER_146_1489 ();
 sg13g2_decap_8 FILLER_146_1496 ();
 sg13g2_decap_8 FILLER_146_1503 ();
 sg13g2_decap_8 FILLER_146_1510 ();
 sg13g2_decap_8 FILLER_146_1517 ();
 sg13g2_decap_8 FILLER_146_1524 ();
 sg13g2_decap_8 FILLER_146_1531 ();
 sg13g2_decap_8 FILLER_146_1538 ();
 sg13g2_decap_8 FILLER_146_1545 ();
 sg13g2_decap_8 FILLER_146_1552 ();
 sg13g2_decap_8 FILLER_146_1559 ();
 sg13g2_decap_8 FILLER_146_1566 ();
 sg13g2_decap_8 FILLER_146_1573 ();
 sg13g2_decap_8 FILLER_146_1580 ();
 sg13g2_decap_8 FILLER_146_1587 ();
 sg13g2_decap_8 FILLER_146_1594 ();
 sg13g2_decap_8 FILLER_146_1601 ();
 sg13g2_decap_8 FILLER_146_1608 ();
 sg13g2_decap_8 FILLER_146_1615 ();
 sg13g2_fill_2 FILLER_146_1622 ();
 sg13g2_fill_1 FILLER_146_1624 ();
 sg13g2_fill_2 FILLER_147_26 ();
 sg13g2_fill_1 FILLER_147_28 ();
 sg13g2_fill_1 FILLER_147_33 ();
 sg13g2_fill_2 FILLER_147_39 ();
 sg13g2_fill_1 FILLER_147_46 ();
 sg13g2_fill_2 FILLER_147_53 ();
 sg13g2_fill_2 FILLER_147_60 ();
 sg13g2_fill_2 FILLER_147_70 ();
 sg13g2_fill_2 FILLER_147_106 ();
 sg13g2_fill_2 FILLER_147_117 ();
 sg13g2_fill_1 FILLER_147_119 ();
 sg13g2_decap_4 FILLER_147_211 ();
 sg13g2_fill_2 FILLER_147_221 ();
 sg13g2_fill_2 FILLER_147_233 ();
 sg13g2_decap_8 FILLER_147_239 ();
 sg13g2_decap_8 FILLER_147_250 ();
 sg13g2_decap_8 FILLER_147_257 ();
 sg13g2_decap_4 FILLER_147_264 ();
 sg13g2_decap_8 FILLER_147_302 ();
 sg13g2_decap_8 FILLER_147_309 ();
 sg13g2_decap_4 FILLER_147_331 ();
 sg13g2_fill_2 FILLER_147_335 ();
 sg13g2_fill_2 FILLER_147_363 ();
 sg13g2_decap_8 FILLER_147_373 ();
 sg13g2_decap_4 FILLER_147_380 ();
 sg13g2_fill_1 FILLER_147_384 ();
 sg13g2_decap_8 FILLER_147_390 ();
 sg13g2_decap_8 FILLER_147_397 ();
 sg13g2_decap_8 FILLER_147_404 ();
 sg13g2_decap_8 FILLER_147_411 ();
 sg13g2_decap_8 FILLER_147_418 ();
 sg13g2_fill_2 FILLER_147_425 ();
 sg13g2_fill_1 FILLER_147_427 ();
 sg13g2_fill_2 FILLER_147_454 ();
 sg13g2_fill_1 FILLER_147_472 ();
 sg13g2_decap_8 FILLER_147_481 ();
 sg13g2_decap_8 FILLER_147_488 ();
 sg13g2_decap_8 FILLER_147_495 ();
 sg13g2_decap_8 FILLER_147_502 ();
 sg13g2_decap_8 FILLER_147_509 ();
 sg13g2_decap_8 FILLER_147_516 ();
 sg13g2_fill_1 FILLER_147_523 ();
 sg13g2_decap_4 FILLER_147_550 ();
 sg13g2_fill_2 FILLER_147_554 ();
 sg13g2_decap_8 FILLER_147_560 ();
 sg13g2_decap_8 FILLER_147_567 ();
 sg13g2_decap_8 FILLER_147_574 ();
 sg13g2_decap_8 FILLER_147_581 ();
 sg13g2_fill_2 FILLER_147_588 ();
 sg13g2_decap_4 FILLER_147_594 ();
 sg13g2_fill_2 FILLER_147_598 ();
 sg13g2_fill_2 FILLER_147_661 ();
 sg13g2_decap_8 FILLER_147_700 ();
 sg13g2_fill_2 FILLER_147_707 ();
 sg13g2_fill_1 FILLER_147_709 ();
 sg13g2_fill_2 FILLER_147_718 ();
 sg13g2_fill_1 FILLER_147_730 ();
 sg13g2_decap_8 FILLER_147_749 ();
 sg13g2_fill_1 FILLER_147_756 ();
 sg13g2_decap_8 FILLER_147_761 ();
 sg13g2_decap_4 FILLER_147_775 ();
 sg13g2_decap_8 FILLER_147_798 ();
 sg13g2_decap_8 FILLER_147_805 ();
 sg13g2_decap_8 FILLER_147_812 ();
 sg13g2_decap_8 FILLER_147_819 ();
 sg13g2_decap_8 FILLER_147_826 ();
 sg13g2_decap_8 FILLER_147_833 ();
 sg13g2_fill_2 FILLER_147_840 ();
 sg13g2_fill_1 FILLER_147_842 ();
 sg13g2_fill_1 FILLER_147_859 ();
 sg13g2_fill_1 FILLER_147_882 ();
 sg13g2_decap_8 FILLER_147_895 ();
 sg13g2_decap_8 FILLER_147_902 ();
 sg13g2_decap_4 FILLER_147_909 ();
 sg13g2_fill_2 FILLER_147_913 ();
 sg13g2_decap_8 FILLER_147_919 ();
 sg13g2_decap_8 FILLER_147_926 ();
 sg13g2_decap_8 FILLER_147_933 ();
 sg13g2_decap_4 FILLER_147_940 ();
 sg13g2_fill_1 FILLER_147_956 ();
 sg13g2_decap_8 FILLER_147_966 ();
 sg13g2_fill_1 FILLER_147_973 ();
 sg13g2_decap_8 FILLER_147_1012 ();
 sg13g2_fill_1 FILLER_147_1024 ();
 sg13g2_fill_2 FILLER_147_1034 ();
 sg13g2_fill_1 FILLER_147_1040 ();
 sg13g2_fill_2 FILLER_147_1067 ();
 sg13g2_fill_1 FILLER_147_1069 ();
 sg13g2_decap_4 FILLER_147_1096 ();
 sg13g2_fill_1 FILLER_147_1100 ();
 sg13g2_decap_8 FILLER_147_1106 ();
 sg13g2_decap_4 FILLER_147_1113 ();
 sg13g2_fill_2 FILLER_147_1117 ();
 sg13g2_decap_4 FILLER_147_1127 ();
 sg13g2_fill_1 FILLER_147_1157 ();
 sg13g2_fill_1 FILLER_147_1161 ();
 sg13g2_decap_8 FILLER_147_1170 ();
 sg13g2_decap_8 FILLER_147_1177 ();
 sg13g2_decap_8 FILLER_147_1184 ();
 sg13g2_decap_4 FILLER_147_1191 ();
 sg13g2_fill_2 FILLER_147_1195 ();
 sg13g2_fill_1 FILLER_147_1227 ();
 sg13g2_fill_1 FILLER_147_1240 ();
 sg13g2_fill_1 FILLER_147_1249 ();
 sg13g2_fill_2 FILLER_147_1254 ();
 sg13g2_decap_8 FILLER_147_1260 ();
 sg13g2_fill_2 FILLER_147_1267 ();
 sg13g2_fill_1 FILLER_147_1269 ();
 sg13g2_decap_8 FILLER_147_1278 ();
 sg13g2_fill_2 FILLER_147_1285 ();
 sg13g2_decap_8 FILLER_147_1291 ();
 sg13g2_decap_8 FILLER_147_1298 ();
 sg13g2_decap_8 FILLER_147_1305 ();
 sg13g2_decap_8 FILLER_147_1312 ();
 sg13g2_decap_8 FILLER_147_1319 ();
 sg13g2_decap_8 FILLER_147_1326 ();
 sg13g2_decap_8 FILLER_147_1333 ();
 sg13g2_decap_8 FILLER_147_1340 ();
 sg13g2_decap_8 FILLER_147_1347 ();
 sg13g2_decap_8 FILLER_147_1354 ();
 sg13g2_decap_8 FILLER_147_1361 ();
 sg13g2_decap_8 FILLER_147_1368 ();
 sg13g2_decap_8 FILLER_147_1375 ();
 sg13g2_decap_8 FILLER_147_1382 ();
 sg13g2_decap_8 FILLER_147_1389 ();
 sg13g2_decap_8 FILLER_147_1396 ();
 sg13g2_decap_8 FILLER_147_1403 ();
 sg13g2_decap_8 FILLER_147_1410 ();
 sg13g2_decap_8 FILLER_147_1417 ();
 sg13g2_decap_8 FILLER_147_1424 ();
 sg13g2_decap_8 FILLER_147_1431 ();
 sg13g2_decap_8 FILLER_147_1438 ();
 sg13g2_decap_8 FILLER_147_1445 ();
 sg13g2_decap_8 FILLER_147_1452 ();
 sg13g2_decap_8 FILLER_147_1459 ();
 sg13g2_decap_8 FILLER_147_1466 ();
 sg13g2_decap_8 FILLER_147_1473 ();
 sg13g2_decap_8 FILLER_147_1480 ();
 sg13g2_decap_8 FILLER_147_1487 ();
 sg13g2_decap_8 FILLER_147_1494 ();
 sg13g2_decap_8 FILLER_147_1501 ();
 sg13g2_decap_8 FILLER_147_1508 ();
 sg13g2_decap_8 FILLER_147_1515 ();
 sg13g2_decap_8 FILLER_147_1522 ();
 sg13g2_decap_8 FILLER_147_1529 ();
 sg13g2_decap_8 FILLER_147_1536 ();
 sg13g2_decap_8 FILLER_147_1543 ();
 sg13g2_decap_8 FILLER_147_1550 ();
 sg13g2_decap_8 FILLER_147_1557 ();
 sg13g2_decap_8 FILLER_147_1564 ();
 sg13g2_decap_8 FILLER_147_1571 ();
 sg13g2_decap_8 FILLER_147_1578 ();
 sg13g2_decap_8 FILLER_147_1585 ();
 sg13g2_decap_8 FILLER_147_1592 ();
 sg13g2_decap_8 FILLER_147_1599 ();
 sg13g2_decap_8 FILLER_147_1606 ();
 sg13g2_decap_8 FILLER_147_1613 ();
 sg13g2_decap_4 FILLER_147_1620 ();
 sg13g2_fill_1 FILLER_147_1624 ();
 sg13g2_decap_8 FILLER_148_0 ();
 sg13g2_decap_4 FILLER_148_7 ();
 sg13g2_fill_1 FILLER_148_11 ();
 sg13g2_fill_1 FILLER_148_30 ();
 sg13g2_fill_1 FILLER_148_42 ();
 sg13g2_fill_1 FILLER_148_48 ();
 sg13g2_fill_1 FILLER_148_53 ();
 sg13g2_decap_8 FILLER_148_58 ();
 sg13g2_fill_2 FILLER_148_65 ();
 sg13g2_fill_1 FILLER_148_67 ();
 sg13g2_decap_8 FILLER_148_110 ();
 sg13g2_decap_4 FILLER_148_117 ();
 sg13g2_fill_2 FILLER_148_125 ();
 sg13g2_fill_1 FILLER_148_127 ();
 sg13g2_decap_4 FILLER_148_166 ();
 sg13g2_decap_8 FILLER_148_175 ();
 sg13g2_decap_8 FILLER_148_182 ();
 sg13g2_fill_1 FILLER_148_189 ();
 sg13g2_decap_4 FILLER_148_194 ();
 sg13g2_decap_8 FILLER_148_202 ();
 sg13g2_decap_4 FILLER_148_209 ();
 sg13g2_decap_4 FILLER_148_218 ();
 sg13g2_fill_2 FILLER_148_222 ();
 sg13g2_decap_8 FILLER_148_254 ();
 sg13g2_decap_8 FILLER_148_261 ();
 sg13g2_decap_8 FILLER_148_268 ();
 sg13g2_decap_4 FILLER_148_275 ();
 sg13g2_fill_2 FILLER_148_279 ();
 sg13g2_decap_8 FILLER_148_285 ();
 sg13g2_decap_8 FILLER_148_292 ();
 sg13g2_decap_4 FILLER_148_299 ();
 sg13g2_fill_1 FILLER_148_303 ();
 sg13g2_decap_8 FILLER_148_332 ();
 sg13g2_decap_8 FILLER_148_339 ();
 sg13g2_decap_8 FILLER_148_346 ();
 sg13g2_decap_4 FILLER_148_353 ();
 sg13g2_fill_2 FILLER_148_361 ();
 sg13g2_decap_8 FILLER_148_390 ();
 sg13g2_fill_2 FILLER_148_397 ();
 sg13g2_decap_8 FILLER_148_403 ();
 sg13g2_decap_8 FILLER_148_410 ();
 sg13g2_decap_4 FILLER_148_422 ();
 sg13g2_fill_1 FILLER_148_426 ();
 sg13g2_decap_8 FILLER_148_452 ();
 sg13g2_decap_4 FILLER_148_459 ();
 sg13g2_fill_2 FILLER_148_463 ();
 sg13g2_decap_8 FILLER_148_472 ();
 sg13g2_decap_8 FILLER_148_479 ();
 sg13g2_fill_2 FILLER_148_486 ();
 sg13g2_decap_8 FILLER_148_495 ();
 sg13g2_fill_2 FILLER_148_502 ();
 sg13g2_decap_8 FILLER_148_508 ();
 sg13g2_decap_8 FILLER_148_515 ();
 sg13g2_decap_8 FILLER_148_522 ();
 sg13g2_fill_2 FILLER_148_529 ();
 sg13g2_decap_8 FILLER_148_535 ();
 sg13g2_fill_1 FILLER_148_542 ();
 sg13g2_fill_2 FILLER_148_574 ();
 sg13g2_fill_2 FILLER_148_606 ();
 sg13g2_fill_1 FILLER_148_664 ();
 sg13g2_fill_2 FILLER_148_699 ();
 sg13g2_fill_2 FILLER_148_710 ();
 sg13g2_decap_8 FILLER_148_796 ();
 sg13g2_decap_4 FILLER_148_803 ();
 sg13g2_fill_2 FILLER_148_807 ();
 sg13g2_decap_8 FILLER_148_814 ();
 sg13g2_decap_8 FILLER_148_829 ();
 sg13g2_decap_4 FILLER_148_836 ();
 sg13g2_fill_1 FILLER_148_840 ();
 sg13g2_decap_8 FILLER_148_845 ();
 sg13g2_decap_8 FILLER_148_852 ();
 sg13g2_fill_1 FILLER_148_859 ();
 sg13g2_fill_1 FILLER_148_888 ();
 sg13g2_decap_8 FILLER_148_894 ();
 sg13g2_fill_1 FILLER_148_901 ();
 sg13g2_fill_2 FILLER_148_906 ();
 sg13g2_decap_8 FILLER_148_934 ();
 sg13g2_decap_4 FILLER_148_941 ();
 sg13g2_fill_1 FILLER_148_945 ();
 sg13g2_decap_8 FILLER_148_961 ();
 sg13g2_fill_1 FILLER_148_977 ();
 sg13g2_fill_1 FILLER_148_986 ();
 sg13g2_decap_8 FILLER_148_991 ();
 sg13g2_decap_4 FILLER_148_998 ();
 sg13g2_decap_8 FILLER_148_1008 ();
 sg13g2_fill_2 FILLER_148_1015 ();
 sg13g2_fill_1 FILLER_148_1017 ();
 sg13g2_fill_1 FILLER_148_1030 ();
 sg13g2_decap_4 FILLER_148_1060 ();
 sg13g2_fill_1 FILLER_148_1064 ();
 sg13g2_fill_1 FILLER_148_1070 ();
 sg13g2_fill_2 FILLER_148_1075 ();
 sg13g2_fill_1 FILLER_148_1081 ();
 sg13g2_fill_2 FILLER_148_1087 ();
 sg13g2_fill_1 FILLER_148_1089 ();
 sg13g2_fill_1 FILLER_148_1095 ();
 sg13g2_decap_8 FILLER_148_1115 ();
 sg13g2_decap_8 FILLER_148_1122 ();
 sg13g2_fill_2 FILLER_148_1129 ();
 sg13g2_fill_1 FILLER_148_1168 ();
 sg13g2_decap_8 FILLER_148_1179 ();
 sg13g2_fill_2 FILLER_148_1186 ();
 sg13g2_fill_1 FILLER_148_1188 ();
 sg13g2_decap_8 FILLER_148_1193 ();
 sg13g2_fill_2 FILLER_148_1200 ();
 sg13g2_fill_1 FILLER_148_1202 ();
 sg13g2_decap_4 FILLER_148_1207 ();
 sg13g2_decap_4 FILLER_148_1215 ();
 sg13g2_fill_2 FILLER_148_1219 ();
 sg13g2_decap_8 FILLER_148_1226 ();
 sg13g2_decap_8 FILLER_148_1233 ();
 sg13g2_decap_4 FILLER_148_1240 ();
 sg13g2_fill_1 FILLER_148_1274 ();
 sg13g2_decap_8 FILLER_148_1305 ();
 sg13g2_decap_8 FILLER_148_1312 ();
 sg13g2_decap_8 FILLER_148_1319 ();
 sg13g2_decap_8 FILLER_148_1326 ();
 sg13g2_decap_8 FILLER_148_1333 ();
 sg13g2_decap_8 FILLER_148_1340 ();
 sg13g2_decap_8 FILLER_148_1347 ();
 sg13g2_decap_8 FILLER_148_1354 ();
 sg13g2_decap_8 FILLER_148_1361 ();
 sg13g2_decap_8 FILLER_148_1368 ();
 sg13g2_decap_8 FILLER_148_1375 ();
 sg13g2_decap_8 FILLER_148_1382 ();
 sg13g2_decap_8 FILLER_148_1389 ();
 sg13g2_decap_8 FILLER_148_1396 ();
 sg13g2_decap_8 FILLER_148_1403 ();
 sg13g2_decap_8 FILLER_148_1410 ();
 sg13g2_decap_8 FILLER_148_1417 ();
 sg13g2_decap_8 FILLER_148_1424 ();
 sg13g2_decap_8 FILLER_148_1431 ();
 sg13g2_decap_8 FILLER_148_1438 ();
 sg13g2_decap_8 FILLER_148_1445 ();
 sg13g2_decap_8 FILLER_148_1452 ();
 sg13g2_decap_8 FILLER_148_1459 ();
 sg13g2_decap_8 FILLER_148_1466 ();
 sg13g2_decap_8 FILLER_148_1473 ();
 sg13g2_decap_8 FILLER_148_1480 ();
 sg13g2_decap_8 FILLER_148_1487 ();
 sg13g2_decap_8 FILLER_148_1494 ();
 sg13g2_decap_8 FILLER_148_1501 ();
 sg13g2_decap_8 FILLER_148_1508 ();
 sg13g2_decap_8 FILLER_148_1515 ();
 sg13g2_decap_8 FILLER_148_1522 ();
 sg13g2_decap_8 FILLER_148_1529 ();
 sg13g2_decap_8 FILLER_148_1536 ();
 sg13g2_decap_8 FILLER_148_1543 ();
 sg13g2_decap_8 FILLER_148_1550 ();
 sg13g2_decap_8 FILLER_148_1557 ();
 sg13g2_decap_8 FILLER_148_1564 ();
 sg13g2_decap_8 FILLER_148_1571 ();
 sg13g2_decap_8 FILLER_148_1578 ();
 sg13g2_decap_8 FILLER_148_1585 ();
 sg13g2_decap_8 FILLER_148_1592 ();
 sg13g2_decap_8 FILLER_148_1599 ();
 sg13g2_decap_8 FILLER_148_1606 ();
 sg13g2_decap_8 FILLER_148_1613 ();
 sg13g2_decap_4 FILLER_148_1620 ();
 sg13g2_fill_1 FILLER_148_1624 ();
 sg13g2_decap_8 FILLER_149_0 ();
 sg13g2_decap_4 FILLER_149_7 ();
 sg13g2_fill_2 FILLER_149_16 ();
 sg13g2_decap_4 FILLER_149_23 ();
 sg13g2_fill_2 FILLER_149_41 ();
 sg13g2_fill_2 FILLER_149_61 ();
 sg13g2_fill_2 FILLER_149_82 ();
 sg13g2_fill_2 FILLER_149_171 ();
 sg13g2_fill_1 FILLER_149_178 ();
 sg13g2_decap_8 FILLER_149_185 ();
 sg13g2_decap_4 FILLER_149_192 ();
 sg13g2_decap_8 FILLER_149_205 ();
 sg13g2_decap_8 FILLER_149_212 ();
 sg13g2_fill_2 FILLER_149_219 ();
 sg13g2_decap_8 FILLER_149_238 ();
 sg13g2_decap_8 FILLER_149_245 ();
 sg13g2_decap_4 FILLER_149_252 ();
 sg13g2_decap_8 FILLER_149_260 ();
 sg13g2_decap_4 FILLER_149_267 ();
 sg13g2_fill_2 FILLER_149_271 ();
 sg13g2_fill_1 FILLER_149_301 ();
 sg13g2_fill_1 FILLER_149_313 ();
 sg13g2_fill_1 FILLER_149_318 ();
 sg13g2_decap_4 FILLER_149_331 ();
 sg13g2_fill_2 FILLER_149_340 ();
 sg13g2_decap_8 FILLER_149_371 ();
 sg13g2_fill_2 FILLER_149_378 ();
 sg13g2_fill_2 FILLER_149_383 ();
 sg13g2_fill_1 FILLER_149_385 ();
 sg13g2_fill_1 FILLER_149_390 ();
 sg13g2_decap_8 FILLER_149_443 ();
 sg13g2_decap_8 FILLER_149_450 ();
 sg13g2_decap_8 FILLER_149_457 ();
 sg13g2_decap_8 FILLER_149_464 ();
 sg13g2_decap_8 FILLER_149_471 ();
 sg13g2_fill_1 FILLER_149_478 ();
 sg13g2_fill_2 FILLER_149_489 ();
 sg13g2_fill_2 FILLER_149_522 ();
 sg13g2_fill_1 FILLER_149_524 ();
 sg13g2_decap_4 FILLER_149_560 ();
 sg13g2_decap_4 FILLER_149_568 ();
 sg13g2_decap_4 FILLER_149_575 ();
 sg13g2_fill_2 FILLER_149_646 ();
 sg13g2_fill_1 FILLER_149_653 ();
 sg13g2_decap_8 FILLER_149_664 ();
 sg13g2_fill_1 FILLER_149_674 ();
 sg13g2_decap_8 FILLER_149_679 ();
 sg13g2_decap_8 FILLER_149_686 ();
 sg13g2_fill_1 FILLER_149_693 ();
 sg13g2_fill_2 FILLER_149_699 ();
 sg13g2_fill_1 FILLER_149_716 ();
 sg13g2_decap_4 FILLER_149_742 ();
 sg13g2_decap_8 FILLER_149_756 ();
 sg13g2_fill_2 FILLER_149_763 ();
 sg13g2_decap_8 FILLER_149_791 ();
 sg13g2_decap_8 FILLER_149_798 ();
 sg13g2_fill_2 FILLER_149_814 ();
 sg13g2_decap_8 FILLER_149_842 ();
 sg13g2_fill_1 FILLER_149_855 ();
 sg13g2_decap_8 FILLER_149_866 ();
 sg13g2_fill_1 FILLER_149_873 ();
 sg13g2_decap_4 FILLER_149_879 ();
 sg13g2_fill_1 FILLER_149_883 ();
 sg13g2_decap_8 FILLER_149_900 ();
 sg13g2_decap_8 FILLER_149_907 ();
 sg13g2_fill_1 FILLER_149_914 ();
 sg13g2_fill_2 FILLER_149_920 ();
 sg13g2_decap_8 FILLER_149_932 ();
 sg13g2_fill_1 FILLER_149_939 ();
 sg13g2_decap_8 FILLER_149_944 ();
 sg13g2_fill_2 FILLER_149_951 ();
 sg13g2_fill_1 FILLER_149_953 ();
 sg13g2_decap_8 FILLER_149_964 ();
 sg13g2_decap_4 FILLER_149_971 ();
 sg13g2_fill_1 FILLER_149_975 ();
 sg13g2_decap_8 FILLER_149_1006 ();
 sg13g2_decap_8 FILLER_149_1013 ();
 sg13g2_fill_2 FILLER_149_1020 ();
 sg13g2_fill_1 FILLER_149_1022 ();
 sg13g2_decap_8 FILLER_149_1052 ();
 sg13g2_decap_4 FILLER_149_1059 ();
 sg13g2_fill_2 FILLER_149_1067 ();
 sg13g2_fill_1 FILLER_149_1074 ();
 sg13g2_fill_1 FILLER_149_1105 ();
 sg13g2_decap_8 FILLER_149_1111 ();
 sg13g2_fill_2 FILLER_149_1118 ();
 sg13g2_decap_4 FILLER_149_1127 ();
 sg13g2_decap_8 FILLER_149_1135 ();
 sg13g2_fill_1 FILLER_149_1142 ();
 sg13g2_decap_4 FILLER_149_1168 ();
 sg13g2_fill_1 FILLER_149_1180 ();
 sg13g2_decap_8 FILLER_149_1236 ();
 sg13g2_decap_8 FILLER_149_1243 ();
 sg13g2_decap_8 FILLER_149_1250 ();
 sg13g2_decap_8 FILLER_149_1257 ();
 sg13g2_fill_2 FILLER_149_1268 ();
 sg13g2_fill_1 FILLER_149_1270 ();
 sg13g2_decap_8 FILLER_149_1275 ();
 sg13g2_decap_8 FILLER_149_1282 ();
 sg13g2_decap_8 FILLER_149_1289 ();
 sg13g2_fill_1 FILLER_149_1296 ();
 sg13g2_decap_8 FILLER_149_1301 ();
 sg13g2_decap_8 FILLER_149_1308 ();
 sg13g2_decap_8 FILLER_149_1315 ();
 sg13g2_decap_8 FILLER_149_1322 ();
 sg13g2_decap_8 FILLER_149_1329 ();
 sg13g2_decap_8 FILLER_149_1336 ();
 sg13g2_decap_8 FILLER_149_1343 ();
 sg13g2_decap_8 FILLER_149_1350 ();
 sg13g2_decap_8 FILLER_149_1357 ();
 sg13g2_decap_8 FILLER_149_1364 ();
 sg13g2_decap_8 FILLER_149_1371 ();
 sg13g2_decap_8 FILLER_149_1378 ();
 sg13g2_decap_8 FILLER_149_1385 ();
 sg13g2_decap_8 FILLER_149_1392 ();
 sg13g2_decap_8 FILLER_149_1399 ();
 sg13g2_decap_8 FILLER_149_1406 ();
 sg13g2_decap_8 FILLER_149_1413 ();
 sg13g2_decap_8 FILLER_149_1420 ();
 sg13g2_decap_8 FILLER_149_1427 ();
 sg13g2_decap_8 FILLER_149_1434 ();
 sg13g2_decap_8 FILLER_149_1441 ();
 sg13g2_decap_8 FILLER_149_1448 ();
 sg13g2_decap_8 FILLER_149_1455 ();
 sg13g2_decap_8 FILLER_149_1462 ();
 sg13g2_decap_8 FILLER_149_1469 ();
 sg13g2_decap_8 FILLER_149_1476 ();
 sg13g2_decap_8 FILLER_149_1483 ();
 sg13g2_decap_8 FILLER_149_1490 ();
 sg13g2_decap_8 FILLER_149_1497 ();
 sg13g2_decap_8 FILLER_149_1504 ();
 sg13g2_decap_8 FILLER_149_1511 ();
 sg13g2_decap_8 FILLER_149_1518 ();
 sg13g2_decap_8 FILLER_149_1525 ();
 sg13g2_decap_8 FILLER_149_1532 ();
 sg13g2_decap_8 FILLER_149_1539 ();
 sg13g2_decap_8 FILLER_149_1546 ();
 sg13g2_decap_8 FILLER_149_1553 ();
 sg13g2_decap_8 FILLER_149_1560 ();
 sg13g2_decap_8 FILLER_149_1567 ();
 sg13g2_decap_8 FILLER_149_1574 ();
 sg13g2_decap_8 FILLER_149_1581 ();
 sg13g2_decap_8 FILLER_149_1588 ();
 sg13g2_decap_8 FILLER_149_1595 ();
 sg13g2_decap_8 FILLER_149_1602 ();
 sg13g2_decap_8 FILLER_149_1609 ();
 sg13g2_decap_8 FILLER_149_1616 ();
 sg13g2_fill_2 FILLER_149_1623 ();
 sg13g2_decap_8 FILLER_150_0 ();
 sg13g2_decap_8 FILLER_150_7 ();
 sg13g2_fill_2 FILLER_150_14 ();
 sg13g2_fill_1 FILLER_150_16 ();
 sg13g2_fill_2 FILLER_150_32 ();
 sg13g2_fill_2 FILLER_150_42 ();
 sg13g2_decap_8 FILLER_150_56 ();
 sg13g2_decap_8 FILLER_150_63 ();
 sg13g2_decap_4 FILLER_150_70 ();
 sg13g2_decap_4 FILLER_150_122 ();
 sg13g2_fill_2 FILLER_150_126 ();
 sg13g2_fill_2 FILLER_150_133 ();
 sg13g2_fill_1 FILLER_150_140 ();
 sg13g2_fill_1 FILLER_150_186 ();
 sg13g2_fill_1 FILLER_150_194 ();
 sg13g2_fill_1 FILLER_150_221 ();
 sg13g2_fill_1 FILLER_150_227 ();
 sg13g2_fill_1 FILLER_150_232 ();
 sg13g2_fill_1 FILLER_150_274 ();
 sg13g2_fill_2 FILLER_150_301 ();
 sg13g2_fill_1 FILLER_150_309 ();
 sg13g2_fill_1 FILLER_150_315 ();
 sg13g2_fill_1 FILLER_150_327 ();
 sg13g2_fill_2 FILLER_150_334 ();
 sg13g2_fill_1 FILLER_150_336 ();
 sg13g2_decap_4 FILLER_150_341 ();
 sg13g2_decap_8 FILLER_150_349 ();
 sg13g2_fill_1 FILLER_150_356 ();
 sg13g2_decap_8 FILLER_150_383 ();
 sg13g2_decap_4 FILLER_150_398 ();
 sg13g2_fill_1 FILLER_150_402 ();
 sg13g2_fill_1 FILLER_150_408 ();
 sg13g2_decap_8 FILLER_150_430 ();
 sg13g2_decap_4 FILLER_150_437 ();
 sg13g2_decap_8 FILLER_150_450 ();
 sg13g2_decap_8 FILLER_150_457 ();
 sg13g2_decap_8 FILLER_150_464 ();
 sg13g2_fill_2 FILLER_150_471 ();
 sg13g2_fill_1 FILLER_150_473 ();
 sg13g2_fill_2 FILLER_150_479 ();
 sg13g2_fill_1 FILLER_150_481 ();
 sg13g2_decap_4 FILLER_150_487 ();
 sg13g2_fill_1 FILLER_150_491 ();
 sg13g2_decap_8 FILLER_150_496 ();
 sg13g2_decap_8 FILLER_150_503 ();
 sg13g2_decap_8 FILLER_150_510 ();
 sg13g2_fill_2 FILLER_150_523 ();
 sg13g2_decap_4 FILLER_150_553 ();
 sg13g2_fill_1 FILLER_150_637 ();
 sg13g2_fill_2 FILLER_150_655 ();
 sg13g2_fill_1 FILLER_150_665 ();
 sg13g2_fill_1 FILLER_150_670 ();
 sg13g2_decap_8 FILLER_150_696 ();
 sg13g2_fill_2 FILLER_150_713 ();
 sg13g2_fill_2 FILLER_150_720 ();
 sg13g2_fill_1 FILLER_150_744 ();
 sg13g2_fill_2 FILLER_150_750 ();
 sg13g2_decap_8 FILLER_150_791 ();
 sg13g2_fill_1 FILLER_150_798 ();
 sg13g2_fill_2 FILLER_150_806 ();
 sg13g2_decap_4 FILLER_150_819 ();
 sg13g2_decap_8 FILLER_150_861 ();
 sg13g2_decap_8 FILLER_150_868 ();
 sg13g2_decap_8 FILLER_150_875 ();
 sg13g2_fill_2 FILLER_150_882 ();
 sg13g2_fill_1 FILLER_150_884 ();
 sg13g2_decap_8 FILLER_150_923 ();
 sg13g2_decap_4 FILLER_150_930 ();
 sg13g2_decap_4 FILLER_150_973 ();
 sg13g2_fill_2 FILLER_150_977 ();
 sg13g2_fill_1 FILLER_150_1018 ();
 sg13g2_decap_8 FILLER_150_1025 ();
 sg13g2_decap_8 FILLER_150_1032 ();
 sg13g2_decap_8 FILLER_150_1039 ();
 sg13g2_decap_8 FILLER_150_1046 ();
 sg13g2_fill_2 FILLER_150_1053 ();
 sg13g2_fill_1 FILLER_150_1110 ();
 sg13g2_fill_2 FILLER_150_1116 ();
 sg13g2_fill_1 FILLER_150_1118 ();
 sg13g2_fill_1 FILLER_150_1123 ();
 sg13g2_fill_2 FILLER_150_1150 ();
 sg13g2_decap_8 FILLER_150_1187 ();
 sg13g2_fill_2 FILLER_150_1194 ();
 sg13g2_fill_1 FILLER_150_1196 ();
 sg13g2_fill_1 FILLER_150_1202 ();
 sg13g2_decap_4 FILLER_150_1241 ();
 sg13g2_fill_1 FILLER_150_1245 ();
 sg13g2_decap_4 FILLER_150_1250 ();
 sg13g2_fill_1 FILLER_150_1254 ();
 sg13g2_decap_8 FILLER_150_1314 ();
 sg13g2_decap_8 FILLER_150_1321 ();
 sg13g2_decap_8 FILLER_150_1328 ();
 sg13g2_decap_8 FILLER_150_1335 ();
 sg13g2_decap_8 FILLER_150_1342 ();
 sg13g2_decap_8 FILLER_150_1349 ();
 sg13g2_decap_8 FILLER_150_1356 ();
 sg13g2_decap_8 FILLER_150_1363 ();
 sg13g2_decap_8 FILLER_150_1370 ();
 sg13g2_decap_8 FILLER_150_1377 ();
 sg13g2_decap_8 FILLER_150_1384 ();
 sg13g2_decap_8 FILLER_150_1391 ();
 sg13g2_decap_8 FILLER_150_1398 ();
 sg13g2_decap_8 FILLER_150_1405 ();
 sg13g2_decap_8 FILLER_150_1412 ();
 sg13g2_decap_8 FILLER_150_1419 ();
 sg13g2_decap_8 FILLER_150_1426 ();
 sg13g2_decap_8 FILLER_150_1433 ();
 sg13g2_decap_8 FILLER_150_1440 ();
 sg13g2_decap_8 FILLER_150_1447 ();
 sg13g2_decap_8 FILLER_150_1454 ();
 sg13g2_decap_8 FILLER_150_1461 ();
 sg13g2_decap_8 FILLER_150_1468 ();
 sg13g2_decap_8 FILLER_150_1475 ();
 sg13g2_decap_8 FILLER_150_1482 ();
 sg13g2_decap_8 FILLER_150_1489 ();
 sg13g2_decap_8 FILLER_150_1496 ();
 sg13g2_decap_8 FILLER_150_1503 ();
 sg13g2_decap_8 FILLER_150_1510 ();
 sg13g2_decap_8 FILLER_150_1517 ();
 sg13g2_decap_8 FILLER_150_1524 ();
 sg13g2_decap_8 FILLER_150_1531 ();
 sg13g2_decap_8 FILLER_150_1538 ();
 sg13g2_decap_8 FILLER_150_1545 ();
 sg13g2_decap_8 FILLER_150_1552 ();
 sg13g2_decap_8 FILLER_150_1559 ();
 sg13g2_decap_8 FILLER_150_1566 ();
 sg13g2_decap_8 FILLER_150_1573 ();
 sg13g2_decap_8 FILLER_150_1580 ();
 sg13g2_decap_8 FILLER_150_1587 ();
 sg13g2_decap_8 FILLER_150_1594 ();
 sg13g2_decap_8 FILLER_150_1601 ();
 sg13g2_decap_8 FILLER_150_1608 ();
 sg13g2_decap_8 FILLER_150_1615 ();
 sg13g2_fill_2 FILLER_150_1622 ();
 sg13g2_fill_1 FILLER_150_1624 ();
 sg13g2_decap_8 FILLER_151_0 ();
 sg13g2_decap_8 FILLER_151_7 ();
 sg13g2_decap_4 FILLER_151_14 ();
 sg13g2_fill_2 FILLER_151_18 ();
 sg13g2_decap_4 FILLER_151_30 ();
 sg13g2_fill_1 FILLER_151_34 ();
 sg13g2_decap_8 FILLER_151_51 ();
 sg13g2_decap_8 FILLER_151_58 ();
 sg13g2_decap_8 FILLER_151_65 ();
 sg13g2_decap_8 FILLER_151_72 ();
 sg13g2_fill_2 FILLER_151_79 ();
 sg13g2_fill_1 FILLER_151_81 ();
 sg13g2_decap_4 FILLER_151_86 ();
 sg13g2_decap_8 FILLER_151_121 ();
 sg13g2_decap_8 FILLER_151_128 ();
 sg13g2_fill_2 FILLER_151_135 ();
 sg13g2_fill_2 FILLER_151_181 ();
 sg13g2_decap_4 FILLER_151_217 ();
 sg13g2_fill_1 FILLER_151_221 ();
 sg13g2_decap_8 FILLER_151_237 ();
 sg13g2_decap_8 FILLER_151_244 ();
 sg13g2_fill_1 FILLER_151_251 ();
 sg13g2_decap_8 FILLER_151_277 ();
 sg13g2_decap_8 FILLER_151_284 ();
 sg13g2_decap_8 FILLER_151_291 ();
 sg13g2_fill_2 FILLER_151_298 ();
 sg13g2_decap_4 FILLER_151_304 ();
 sg13g2_decap_8 FILLER_151_328 ();
 sg13g2_fill_2 FILLER_151_335 ();
 sg13g2_fill_1 FILLER_151_337 ();
 sg13g2_decap_8 FILLER_151_364 ();
 sg13g2_decap_8 FILLER_151_371 ();
 sg13g2_decap_8 FILLER_151_378 ();
 sg13g2_fill_2 FILLER_151_430 ();
 sg13g2_fill_1 FILLER_151_432 ();
 sg13g2_fill_1 FILLER_151_437 ();
 sg13g2_fill_2 FILLER_151_464 ();
 sg13g2_fill_1 FILLER_151_466 ();
 sg13g2_fill_2 FILLER_151_473 ();
 sg13g2_fill_1 FILLER_151_475 ();
 sg13g2_decap_8 FILLER_151_481 ();
 sg13g2_fill_2 FILLER_151_491 ();
 sg13g2_fill_1 FILLER_151_493 ();
 sg13g2_decap_8 FILLER_151_499 ();
 sg13g2_decap_8 FILLER_151_506 ();
 sg13g2_decap_4 FILLER_151_513 ();
 sg13g2_decap_8 FILLER_151_522 ();
 sg13g2_fill_1 FILLER_151_529 ();
 sg13g2_decap_8 FILLER_151_540 ();
 sg13g2_fill_1 FILLER_151_592 ();
 sg13g2_fill_1 FILLER_151_622 ();
 sg13g2_decap_8 FILLER_151_627 ();
 sg13g2_fill_1 FILLER_151_634 ();
 sg13g2_fill_2 FILLER_151_640 ();
 sg13g2_fill_1 FILLER_151_642 ();
 sg13g2_fill_2 FILLER_151_652 ();
 sg13g2_fill_1 FILLER_151_654 ();
 sg13g2_fill_2 FILLER_151_685 ();
 sg13g2_fill_1 FILLER_151_687 ();
 sg13g2_decap_4 FILLER_151_694 ();
 sg13g2_fill_2 FILLER_151_718 ();
 sg13g2_fill_1 FILLER_151_730 ();
 sg13g2_fill_2 FILLER_151_759 ();
 sg13g2_decap_4 FILLER_151_801 ();
 sg13g2_decap_4 FILLER_151_810 ();
 sg13g2_fill_2 FILLER_151_814 ();
 sg13g2_fill_2 FILLER_151_855 ();
 sg13g2_decap_8 FILLER_151_862 ();
 sg13g2_decap_8 FILLER_151_869 ();
 sg13g2_decap_8 FILLER_151_876 ();
 sg13g2_decap_4 FILLER_151_883 ();
 sg13g2_fill_1 FILLER_151_887 ();
 sg13g2_fill_2 FILLER_151_914 ();
 sg13g2_fill_1 FILLER_151_916 ();
 sg13g2_decap_8 FILLER_151_921 ();
 sg13g2_decap_8 FILLER_151_928 ();
 sg13g2_decap_4 FILLER_151_935 ();
 sg13g2_fill_2 FILLER_151_939 ();
 sg13g2_fill_2 FILLER_151_945 ();
 sg13g2_decap_8 FILLER_151_976 ();
 sg13g2_fill_1 FILLER_151_983 ();
 sg13g2_decap_8 FILLER_151_988 ();
 sg13g2_decap_8 FILLER_151_995 ();
 sg13g2_decap_8 FILLER_151_1002 ();
 sg13g2_fill_1 FILLER_151_1009 ();
 sg13g2_fill_2 FILLER_151_1016 ();
 sg13g2_fill_1 FILLER_151_1018 ();
 sg13g2_fill_2 FILLER_151_1024 ();
 sg13g2_fill_1 FILLER_151_1026 ();
 sg13g2_decap_8 FILLER_151_1031 ();
 sg13g2_decap_8 FILLER_151_1057 ();
 sg13g2_decap_8 FILLER_151_1064 ();
 sg13g2_decap_8 FILLER_151_1071 ();
 sg13g2_decap_8 FILLER_151_1078 ();
 sg13g2_decap_4 FILLER_151_1085 ();
 sg13g2_fill_1 FILLER_151_1089 ();
 sg13g2_fill_2 FILLER_151_1094 ();
 sg13g2_fill_1 FILLER_151_1096 ();
 sg13g2_decap_8 FILLER_151_1101 ();
 sg13g2_decap_8 FILLER_151_1108 ();
 sg13g2_decap_8 FILLER_151_1127 ();
 sg13g2_decap_8 FILLER_151_1134 ();
 sg13g2_fill_2 FILLER_151_1141 ();
 sg13g2_decap_8 FILLER_151_1146 ();
 sg13g2_fill_2 FILLER_151_1157 ();
 sg13g2_decap_8 FILLER_151_1163 ();
 sg13g2_decap_8 FILLER_151_1170 ();
 sg13g2_decap_4 FILLER_151_1177 ();
 sg13g2_fill_2 FILLER_151_1181 ();
 sg13g2_decap_4 FILLER_151_1191 ();
 sg13g2_fill_2 FILLER_151_1195 ();
 sg13g2_decap_4 FILLER_151_1206 ();
 sg13g2_fill_2 FILLER_151_1210 ();
 sg13g2_decap_8 FILLER_151_1217 ();
 sg13g2_decap_8 FILLER_151_1224 ();
 sg13g2_fill_2 FILLER_151_1231 ();
 sg13g2_fill_1 FILLER_151_1233 ();
 sg13g2_decap_8 FILLER_151_1316 ();
 sg13g2_decap_8 FILLER_151_1323 ();
 sg13g2_decap_8 FILLER_151_1330 ();
 sg13g2_decap_8 FILLER_151_1337 ();
 sg13g2_decap_8 FILLER_151_1344 ();
 sg13g2_decap_8 FILLER_151_1351 ();
 sg13g2_decap_8 FILLER_151_1358 ();
 sg13g2_decap_8 FILLER_151_1365 ();
 sg13g2_decap_8 FILLER_151_1372 ();
 sg13g2_decap_8 FILLER_151_1379 ();
 sg13g2_decap_8 FILLER_151_1386 ();
 sg13g2_decap_8 FILLER_151_1393 ();
 sg13g2_decap_8 FILLER_151_1400 ();
 sg13g2_decap_8 FILLER_151_1407 ();
 sg13g2_decap_8 FILLER_151_1414 ();
 sg13g2_decap_8 FILLER_151_1421 ();
 sg13g2_decap_8 FILLER_151_1428 ();
 sg13g2_decap_8 FILLER_151_1435 ();
 sg13g2_decap_8 FILLER_151_1442 ();
 sg13g2_decap_8 FILLER_151_1449 ();
 sg13g2_decap_8 FILLER_151_1456 ();
 sg13g2_decap_8 FILLER_151_1463 ();
 sg13g2_decap_8 FILLER_151_1470 ();
 sg13g2_decap_8 FILLER_151_1477 ();
 sg13g2_decap_8 FILLER_151_1484 ();
 sg13g2_decap_8 FILLER_151_1491 ();
 sg13g2_decap_8 FILLER_151_1498 ();
 sg13g2_decap_8 FILLER_151_1505 ();
 sg13g2_decap_8 FILLER_151_1512 ();
 sg13g2_decap_8 FILLER_151_1519 ();
 sg13g2_decap_8 FILLER_151_1526 ();
 sg13g2_decap_8 FILLER_151_1533 ();
 sg13g2_decap_8 FILLER_151_1540 ();
 sg13g2_decap_8 FILLER_151_1547 ();
 sg13g2_decap_8 FILLER_151_1554 ();
 sg13g2_decap_8 FILLER_151_1561 ();
 sg13g2_decap_8 FILLER_151_1568 ();
 sg13g2_decap_8 FILLER_151_1575 ();
 sg13g2_decap_8 FILLER_151_1582 ();
 sg13g2_decap_8 FILLER_151_1589 ();
 sg13g2_decap_8 FILLER_151_1596 ();
 sg13g2_decap_8 FILLER_151_1603 ();
 sg13g2_decap_8 FILLER_151_1610 ();
 sg13g2_decap_8 FILLER_151_1617 ();
 sg13g2_fill_1 FILLER_151_1624 ();
 sg13g2_decap_8 FILLER_152_0 ();
 sg13g2_decap_4 FILLER_152_11 ();
 sg13g2_fill_2 FILLER_152_15 ();
 sg13g2_fill_2 FILLER_152_38 ();
 sg13g2_fill_1 FILLER_152_40 ();
 sg13g2_decap_8 FILLER_152_46 ();
 sg13g2_decap_8 FILLER_152_53 ();
 sg13g2_decap_4 FILLER_152_60 ();
 sg13g2_decap_4 FILLER_152_67 ();
 sg13g2_fill_2 FILLER_152_71 ();
 sg13g2_decap_8 FILLER_152_81 ();
 sg13g2_decap_8 FILLER_152_88 ();
 sg13g2_fill_2 FILLER_152_95 ();
 sg13g2_fill_2 FILLER_152_100 ();
 sg13g2_fill_1 FILLER_152_111 ();
 sg13g2_fill_1 FILLER_152_134 ();
 sg13g2_decap_8 FILLER_152_140 ();
 sg13g2_decap_8 FILLER_152_147 ();
 sg13g2_decap_4 FILLER_152_154 ();
 sg13g2_decap_8 FILLER_152_166 ();
 sg13g2_decap_8 FILLER_152_173 ();
 sg13g2_decap_8 FILLER_152_180 ();
 sg13g2_fill_2 FILLER_152_198 ();
 sg13g2_fill_2 FILLER_152_205 ();
 sg13g2_decap_8 FILLER_152_215 ();
 sg13g2_decap_8 FILLER_152_222 ();
 sg13g2_decap_4 FILLER_152_229 ();
 sg13g2_decap_8 FILLER_152_274 ();
 sg13g2_decap_4 FILLER_152_281 ();
 sg13g2_fill_1 FILLER_152_285 ();
 sg13g2_decap_8 FILLER_152_291 ();
 sg13g2_decap_8 FILLER_152_298 ();
 sg13g2_decap_8 FILLER_152_305 ();
 sg13g2_decap_8 FILLER_152_312 ();
 sg13g2_decap_8 FILLER_152_319 ();
 sg13g2_decap_8 FILLER_152_326 ();
 sg13g2_fill_2 FILLER_152_333 ();
 sg13g2_decap_8 FILLER_152_340 ();
 sg13g2_decap_8 FILLER_152_347 ();
 sg13g2_fill_2 FILLER_152_354 ();
 sg13g2_fill_1 FILLER_152_356 ();
 sg13g2_decap_4 FILLER_152_386 ();
 sg13g2_decap_8 FILLER_152_425 ();
 sg13g2_fill_2 FILLER_152_432 ();
 sg13g2_fill_2 FILLER_152_438 ();
 sg13g2_decap_4 FILLER_152_445 ();
 sg13g2_fill_2 FILLER_152_449 ();
 sg13g2_fill_2 FILLER_152_458 ();
 sg13g2_fill_1 FILLER_152_490 ();
 sg13g2_decap_8 FILLER_152_499 ();
 sg13g2_decap_8 FILLER_152_506 ();
 sg13g2_decap_4 FILLER_152_513 ();
 sg13g2_fill_2 FILLER_152_517 ();
 sg13g2_decap_4 FILLER_152_549 ();
 sg13g2_decap_8 FILLER_152_566 ();
 sg13g2_fill_2 FILLER_152_583 ();
 sg13g2_fill_1 FILLER_152_589 ();
 sg13g2_decap_8 FILLER_152_642 ();
 sg13g2_decap_8 FILLER_152_649 ();
 sg13g2_decap_8 FILLER_152_660 ();
 sg13g2_decap_8 FILLER_152_667 ();
 sg13g2_decap_8 FILLER_152_674 ();
 sg13g2_decap_4 FILLER_152_681 ();
 sg13g2_fill_2 FILLER_152_685 ();
 sg13g2_decap_4 FILLER_152_692 ();
 sg13g2_fill_1 FILLER_152_696 ();
 sg13g2_fill_2 FILLER_152_727 ();
 sg13g2_decap_8 FILLER_152_738 ();
 sg13g2_decap_4 FILLER_152_752 ();
 sg13g2_fill_2 FILLER_152_792 ();
 sg13g2_fill_1 FILLER_152_794 ();
 sg13g2_fill_1 FILLER_152_806 ();
 sg13g2_fill_1 FILLER_152_812 ();
 sg13g2_fill_2 FILLER_152_829 ();
 sg13g2_fill_2 FILLER_152_849 ();
 sg13g2_fill_1 FILLER_152_851 ();
 sg13g2_fill_2 FILLER_152_861 ();
 sg13g2_fill_1 FILLER_152_863 ();
 sg13g2_fill_1 FILLER_152_895 ();
 sg13g2_decap_4 FILLER_152_903 ();
 sg13g2_fill_2 FILLER_152_907 ();
 sg13g2_fill_2 FILLER_152_961 ();
 sg13g2_fill_1 FILLER_152_963 ();
 sg13g2_fill_2 FILLER_152_969 ();
 sg13g2_decap_4 FILLER_152_1002 ();
 sg13g2_fill_2 FILLER_152_1011 ();
 sg13g2_fill_2 FILLER_152_1019 ();
 sg13g2_decap_4 FILLER_152_1065 ();
 sg13g2_decap_4 FILLER_152_1073 ();
 sg13g2_fill_1 FILLER_152_1077 ();
 sg13g2_decap_8 FILLER_152_1087 ();
 sg13g2_decap_8 FILLER_152_1094 ();
 sg13g2_decap_8 FILLER_152_1101 ();
 sg13g2_decap_8 FILLER_152_1108 ();
 sg13g2_decap_4 FILLER_152_1115 ();
 sg13g2_fill_1 FILLER_152_1119 ();
 sg13g2_decap_8 FILLER_152_1125 ();
 sg13g2_decap_4 FILLER_152_1132 ();
 sg13g2_fill_2 FILLER_152_1136 ();
 sg13g2_fill_1 FILLER_152_1142 ();
 sg13g2_decap_8 FILLER_152_1148 ();
 sg13g2_decap_8 FILLER_152_1155 ();
 sg13g2_decap_8 FILLER_152_1162 ();
 sg13g2_decap_8 FILLER_152_1169 ();
 sg13g2_decap_4 FILLER_152_1176 ();
 sg13g2_fill_1 FILLER_152_1180 ();
 sg13g2_decap_8 FILLER_152_1215 ();
 sg13g2_decap_8 FILLER_152_1222 ();
 sg13g2_fill_2 FILLER_152_1229 ();
 sg13g2_fill_1 FILLER_152_1231 ();
 sg13g2_decap_4 FILLER_152_1255 ();
 sg13g2_fill_2 FILLER_152_1259 ();
 sg13g2_decap_8 FILLER_152_1269 ();
 sg13g2_decap_8 FILLER_152_1276 ();
 sg13g2_fill_2 FILLER_152_1283 ();
 sg13g2_decap_8 FILLER_152_1293 ();
 sg13g2_decap_8 FILLER_152_1304 ();
 sg13g2_decap_8 FILLER_152_1311 ();
 sg13g2_decap_8 FILLER_152_1318 ();
 sg13g2_decap_8 FILLER_152_1325 ();
 sg13g2_decap_8 FILLER_152_1332 ();
 sg13g2_decap_8 FILLER_152_1339 ();
 sg13g2_decap_8 FILLER_152_1346 ();
 sg13g2_decap_8 FILLER_152_1353 ();
 sg13g2_decap_8 FILLER_152_1360 ();
 sg13g2_decap_8 FILLER_152_1367 ();
 sg13g2_decap_8 FILLER_152_1374 ();
 sg13g2_decap_8 FILLER_152_1381 ();
 sg13g2_decap_8 FILLER_152_1388 ();
 sg13g2_decap_8 FILLER_152_1395 ();
 sg13g2_decap_8 FILLER_152_1402 ();
 sg13g2_decap_8 FILLER_152_1409 ();
 sg13g2_decap_8 FILLER_152_1416 ();
 sg13g2_decap_8 FILLER_152_1423 ();
 sg13g2_decap_8 FILLER_152_1430 ();
 sg13g2_decap_8 FILLER_152_1437 ();
 sg13g2_decap_8 FILLER_152_1444 ();
 sg13g2_decap_8 FILLER_152_1451 ();
 sg13g2_decap_8 FILLER_152_1458 ();
 sg13g2_decap_8 FILLER_152_1465 ();
 sg13g2_decap_8 FILLER_152_1472 ();
 sg13g2_decap_8 FILLER_152_1479 ();
 sg13g2_decap_8 FILLER_152_1486 ();
 sg13g2_decap_8 FILLER_152_1493 ();
 sg13g2_decap_8 FILLER_152_1500 ();
 sg13g2_decap_8 FILLER_152_1507 ();
 sg13g2_decap_8 FILLER_152_1514 ();
 sg13g2_decap_8 FILLER_152_1521 ();
 sg13g2_decap_8 FILLER_152_1528 ();
 sg13g2_decap_8 FILLER_152_1535 ();
 sg13g2_decap_8 FILLER_152_1542 ();
 sg13g2_decap_8 FILLER_152_1549 ();
 sg13g2_decap_8 FILLER_152_1556 ();
 sg13g2_decap_8 FILLER_152_1563 ();
 sg13g2_decap_8 FILLER_152_1570 ();
 sg13g2_decap_8 FILLER_152_1577 ();
 sg13g2_decap_8 FILLER_152_1584 ();
 sg13g2_decap_8 FILLER_152_1591 ();
 sg13g2_decap_8 FILLER_152_1598 ();
 sg13g2_decap_8 FILLER_152_1605 ();
 sg13g2_decap_8 FILLER_152_1612 ();
 sg13g2_decap_4 FILLER_152_1619 ();
 sg13g2_fill_2 FILLER_152_1623 ();
 sg13g2_fill_1 FILLER_153_0 ();
 sg13g2_decap_8 FILLER_153_27 ();
 sg13g2_decap_8 FILLER_153_49 ();
 sg13g2_decap_4 FILLER_153_56 ();
 sg13g2_fill_1 FILLER_153_60 ();
 sg13g2_fill_1 FILLER_153_72 ();
 sg13g2_decap_4 FILLER_153_78 ();
 sg13g2_decap_8 FILLER_153_100 ();
 sg13g2_fill_2 FILLER_153_107 ();
 sg13g2_fill_2 FILLER_153_114 ();
 sg13g2_fill_2 FILLER_153_121 ();
 sg13g2_decap_8 FILLER_153_136 ();
 sg13g2_decap_8 FILLER_153_143 ();
 sg13g2_decap_8 FILLER_153_150 ();
 sg13g2_decap_8 FILLER_153_157 ();
 sg13g2_decap_4 FILLER_153_164 ();
 sg13g2_fill_1 FILLER_153_168 ();
 sg13g2_decap_8 FILLER_153_173 ();
 sg13g2_decap_8 FILLER_153_180 ();
 sg13g2_fill_2 FILLER_153_201 ();
 sg13g2_fill_1 FILLER_153_203 ();
 sg13g2_fill_1 FILLER_153_230 ();
 sg13g2_decap_8 FILLER_153_235 ();
 sg13g2_decap_8 FILLER_153_242 ();
 sg13g2_decap_8 FILLER_153_249 ();
 sg13g2_decap_4 FILLER_153_260 ();
 sg13g2_fill_2 FILLER_153_303 ();
 sg13g2_decap_4 FILLER_153_309 ();
 sg13g2_fill_1 FILLER_153_313 ();
 sg13g2_fill_2 FILLER_153_324 ();
 sg13g2_fill_2 FILLER_153_381 ();
 sg13g2_decap_4 FILLER_153_386 ();
 sg13g2_decap_4 FILLER_153_395 ();
 sg13g2_fill_2 FILLER_153_404 ();
 sg13g2_fill_1 FILLER_153_406 ();
 sg13g2_decap_8 FILLER_153_411 ();
 sg13g2_fill_2 FILLER_153_453 ();
 sg13g2_fill_1 FILLER_153_455 ();
 sg13g2_decap_8 FILLER_153_539 ();
 sg13g2_decap_8 FILLER_153_546 ();
 sg13g2_decap_8 FILLER_153_553 ();
 sg13g2_decap_8 FILLER_153_560 ();
 sg13g2_decap_8 FILLER_153_567 ();
 sg13g2_decap_8 FILLER_153_574 ();
 sg13g2_fill_1 FILLER_153_581 ();
 sg13g2_decap_8 FILLER_153_592 ();
 sg13g2_decap_8 FILLER_153_599 ();
 sg13g2_decap_8 FILLER_153_606 ();
 sg13g2_decap_8 FILLER_153_613 ();
 sg13g2_decap_8 FILLER_153_620 ();
 sg13g2_decap_8 FILLER_153_627 ();
 sg13g2_decap_4 FILLER_153_634 ();
 sg13g2_fill_2 FILLER_153_638 ();
 sg13g2_decap_8 FILLER_153_676 ();
 sg13g2_decap_8 FILLER_153_683 ();
 sg13g2_decap_4 FILLER_153_690 ();
 sg13g2_fill_2 FILLER_153_699 ();
 sg13g2_fill_2 FILLER_153_710 ();
 sg13g2_fill_1 FILLER_153_712 ();
 sg13g2_fill_2 FILLER_153_737 ();
 sg13g2_fill_1 FILLER_153_739 ();
 sg13g2_decap_4 FILLER_153_803 ();
 sg13g2_fill_1 FILLER_153_807 ();
 sg13g2_fill_1 FILLER_153_811 ();
 sg13g2_decap_8 FILLER_153_817 ();
 sg13g2_decap_8 FILLER_153_824 ();
 sg13g2_decap_8 FILLER_153_831 ();
 sg13g2_fill_2 FILLER_153_843 ();
 sg13g2_fill_1 FILLER_153_845 ();
 sg13g2_decap_8 FILLER_153_876 ();
 sg13g2_fill_2 FILLER_153_883 ();
 sg13g2_fill_1 FILLER_153_915 ();
 sg13g2_decap_8 FILLER_153_920 ();
 sg13g2_decap_4 FILLER_153_927 ();
 sg13g2_fill_1 FILLER_153_931 ();
 sg13g2_fill_1 FILLER_153_962 ();
 sg13g2_fill_1 FILLER_153_968 ();
 sg13g2_decap_8 FILLER_153_975 ();
 sg13g2_decap_8 FILLER_153_982 ();
 sg13g2_decap_8 FILLER_153_989 ();
 sg13g2_decap_8 FILLER_153_996 ();
 sg13g2_decap_8 FILLER_153_1016 ();
 sg13g2_fill_2 FILLER_153_1028 ();
 sg13g2_fill_1 FILLER_153_1030 ();
 sg13g2_fill_2 FILLER_153_1057 ();
 sg13g2_fill_1 FILLER_153_1059 ();
 sg13g2_fill_2 FILLER_153_1114 ();
 sg13g2_fill_1 FILLER_153_1116 ();
 sg13g2_fill_1 FILLER_153_1121 ();
 sg13g2_decap_8 FILLER_153_1155 ();
 sg13g2_decap_8 FILLER_153_1174 ();
 sg13g2_decap_4 FILLER_153_1181 ();
 sg13g2_fill_2 FILLER_153_1192 ();
 sg13g2_fill_1 FILLER_153_1194 ();
 sg13g2_decap_8 FILLER_153_1211 ();
 sg13g2_decap_4 FILLER_153_1218 ();
 sg13g2_fill_1 FILLER_153_1222 ();
 sg13g2_fill_2 FILLER_153_1235 ();
 sg13g2_decap_8 FILLER_153_1266 ();
 sg13g2_decap_8 FILLER_153_1273 ();
 sg13g2_decap_8 FILLER_153_1280 ();
 sg13g2_decap_8 FILLER_153_1317 ();
 sg13g2_decap_8 FILLER_153_1328 ();
 sg13g2_decap_8 FILLER_153_1335 ();
 sg13g2_decap_8 FILLER_153_1342 ();
 sg13g2_decap_8 FILLER_153_1349 ();
 sg13g2_decap_8 FILLER_153_1356 ();
 sg13g2_decap_8 FILLER_153_1363 ();
 sg13g2_decap_8 FILLER_153_1370 ();
 sg13g2_decap_8 FILLER_153_1377 ();
 sg13g2_decap_8 FILLER_153_1384 ();
 sg13g2_decap_8 FILLER_153_1391 ();
 sg13g2_decap_8 FILLER_153_1398 ();
 sg13g2_decap_8 FILLER_153_1405 ();
 sg13g2_decap_8 FILLER_153_1412 ();
 sg13g2_decap_8 FILLER_153_1419 ();
 sg13g2_decap_8 FILLER_153_1426 ();
 sg13g2_decap_8 FILLER_153_1433 ();
 sg13g2_decap_8 FILLER_153_1440 ();
 sg13g2_decap_8 FILLER_153_1447 ();
 sg13g2_decap_8 FILLER_153_1454 ();
 sg13g2_decap_8 FILLER_153_1461 ();
 sg13g2_decap_8 FILLER_153_1468 ();
 sg13g2_decap_8 FILLER_153_1475 ();
 sg13g2_decap_8 FILLER_153_1482 ();
 sg13g2_decap_8 FILLER_153_1489 ();
 sg13g2_decap_8 FILLER_153_1496 ();
 sg13g2_decap_8 FILLER_153_1503 ();
 sg13g2_decap_8 FILLER_153_1510 ();
 sg13g2_decap_8 FILLER_153_1517 ();
 sg13g2_decap_8 FILLER_153_1524 ();
 sg13g2_decap_8 FILLER_153_1531 ();
 sg13g2_decap_8 FILLER_153_1538 ();
 sg13g2_decap_8 FILLER_153_1545 ();
 sg13g2_decap_8 FILLER_153_1552 ();
 sg13g2_decap_8 FILLER_153_1559 ();
 sg13g2_decap_8 FILLER_153_1566 ();
 sg13g2_decap_8 FILLER_153_1573 ();
 sg13g2_decap_8 FILLER_153_1580 ();
 sg13g2_decap_8 FILLER_153_1587 ();
 sg13g2_decap_8 FILLER_153_1594 ();
 sg13g2_decap_8 FILLER_153_1601 ();
 sg13g2_decap_8 FILLER_153_1608 ();
 sg13g2_decap_8 FILLER_153_1615 ();
 sg13g2_fill_2 FILLER_153_1622 ();
 sg13g2_fill_1 FILLER_153_1624 ();
 sg13g2_decap_8 FILLER_154_0 ();
 sg13g2_decap_4 FILLER_154_7 ();
 sg13g2_fill_2 FILLER_154_11 ();
 sg13g2_decap_8 FILLER_154_17 ();
 sg13g2_decap_8 FILLER_154_24 ();
 sg13g2_fill_2 FILLER_154_31 ();
 sg13g2_fill_1 FILLER_154_33 ();
 sg13g2_decap_4 FILLER_154_39 ();
 sg13g2_decap_4 FILLER_154_47 ();
 sg13g2_decap_4 FILLER_154_91 ();
 sg13g2_fill_2 FILLER_154_95 ();
 sg13g2_fill_2 FILLER_154_112 ();
 sg13g2_decap_8 FILLER_154_127 ();
 sg13g2_decap_4 FILLER_154_134 ();
 sg13g2_decap_8 FILLER_154_143 ();
 sg13g2_fill_2 FILLER_154_150 ();
 sg13g2_decap_8 FILLER_154_156 ();
 sg13g2_decap_8 FILLER_154_250 ();
 sg13g2_decap_8 FILLER_154_257 ();
 sg13g2_decap_8 FILLER_154_264 ();
 sg13g2_fill_1 FILLER_154_271 ();
 sg13g2_decap_8 FILLER_154_276 ();
 sg13g2_decap_8 FILLER_154_283 ();
 sg13g2_fill_2 FILLER_154_290 ();
 sg13g2_fill_1 FILLER_154_292 ();
 sg13g2_decap_4 FILLER_154_323 ();
 sg13g2_decap_8 FILLER_154_336 ();
 sg13g2_fill_1 FILLER_154_369 ();
 sg13g2_fill_2 FILLER_154_373 ();
 sg13g2_decap_4 FILLER_154_380 ();
 sg13g2_fill_1 FILLER_154_384 ();
 sg13g2_fill_2 FILLER_154_394 ();
 sg13g2_decap_4 FILLER_154_400 ();
 sg13g2_decap_8 FILLER_154_408 ();
 sg13g2_decap_8 FILLER_154_415 ();
 sg13g2_decap_8 FILLER_154_422 ();
 sg13g2_decap_8 FILLER_154_429 ();
 sg13g2_fill_2 FILLER_154_436 ();
 sg13g2_fill_1 FILLER_154_438 ();
 sg13g2_decap_4 FILLER_154_477 ();
 sg13g2_decap_8 FILLER_154_485 ();
 sg13g2_decap_8 FILLER_154_492 ();
 sg13g2_decap_8 FILLER_154_499 ();
 sg13g2_fill_2 FILLER_154_506 ();
 sg13g2_decap_4 FILLER_154_512 ();
 sg13g2_fill_1 FILLER_154_516 ();
 sg13g2_decap_8 FILLER_154_522 ();
 sg13g2_fill_2 FILLER_154_529 ();
 sg13g2_fill_1 FILLER_154_531 ();
 sg13g2_decap_8 FILLER_154_538 ();
 sg13g2_decap_8 FILLER_154_545 ();
 sg13g2_decap_4 FILLER_154_557 ();
 sg13g2_fill_1 FILLER_154_561 ();
 sg13g2_fill_2 FILLER_154_581 ();
 sg13g2_decap_8 FILLER_154_592 ();
 sg13g2_fill_1 FILLER_154_599 ();
 sg13g2_decap_8 FILLER_154_604 ();
 sg13g2_decap_8 FILLER_154_611 ();
 sg13g2_decap_8 FILLER_154_618 ();
 sg13g2_fill_2 FILLER_154_625 ();
 sg13g2_fill_1 FILLER_154_627 ();
 sg13g2_decap_8 FILLER_154_632 ();
 sg13g2_decap_8 FILLER_154_639 ();
 sg13g2_decap_4 FILLER_154_646 ();
 sg13g2_fill_2 FILLER_154_650 ();
 sg13g2_fill_1 FILLER_154_662 ();
 sg13g2_decap_4 FILLER_154_707 ();
 sg13g2_fill_2 FILLER_154_711 ();
 sg13g2_decap_8 FILLER_154_747 ();
 sg13g2_decap_8 FILLER_154_754 ();
 sg13g2_decap_8 FILLER_154_761 ();
 sg13g2_fill_1 FILLER_154_768 ();
 sg13g2_fill_2 FILLER_154_804 ();
 sg13g2_decap_8 FILLER_154_810 ();
 sg13g2_decap_4 FILLER_154_817 ();
 sg13g2_fill_1 FILLER_154_821 ();
 sg13g2_decap_4 FILLER_154_847 ();
 sg13g2_fill_2 FILLER_154_851 ();
 sg13g2_decap_8 FILLER_154_858 ();
 sg13g2_decap_8 FILLER_154_865 ();
 sg13g2_decap_8 FILLER_154_872 ();
 sg13g2_decap_4 FILLER_154_879 ();
 sg13g2_fill_1 FILLER_154_883 ();
 sg13g2_decap_4 FILLER_154_890 ();
 sg13g2_fill_2 FILLER_154_894 ();
 sg13g2_fill_2 FILLER_154_905 ();
 sg13g2_fill_1 FILLER_154_907 ();
 sg13g2_decap_4 FILLER_154_934 ();
 sg13g2_fill_1 FILLER_154_938 ();
 sg13g2_decap_8 FILLER_154_943 ();
 sg13g2_decap_8 FILLER_154_950 ();
 sg13g2_decap_8 FILLER_154_957 ();
 sg13g2_decap_8 FILLER_154_964 ();
 sg13g2_fill_1 FILLER_154_971 ();
 sg13g2_decap_4 FILLER_154_977 ();
 sg13g2_fill_1 FILLER_154_981 ();
 sg13g2_decap_8 FILLER_154_986 ();
 sg13g2_decap_4 FILLER_154_993 ();
 sg13g2_fill_2 FILLER_154_997 ();
 sg13g2_decap_4 FILLER_154_1008 ();
 sg13g2_fill_1 FILLER_154_1012 ();
 sg13g2_fill_1 FILLER_154_1022 ();
 sg13g2_fill_2 FILLER_154_1033 ();
 sg13g2_fill_1 FILLER_154_1066 ();
 sg13g2_decap_8 FILLER_154_1077 ();
 sg13g2_fill_2 FILLER_154_1084 ();
 sg13g2_fill_1 FILLER_154_1086 ();
 sg13g2_decap_4 FILLER_154_1097 ();
 sg13g2_fill_2 FILLER_154_1101 ();
 sg13g2_decap_8 FILLER_154_1132 ();
 sg13g2_decap_8 FILLER_154_1139 ();
 sg13g2_decap_8 FILLER_154_1146 ();
 sg13g2_fill_1 FILLER_154_1183 ();
 sg13g2_decap_8 FILLER_154_1190 ();
 sg13g2_decap_8 FILLER_154_1197 ();
 sg13g2_decap_8 FILLER_154_1204 ();
 sg13g2_fill_2 FILLER_154_1211 ();
 sg13g2_decap_8 FILLER_154_1292 ();
 sg13g2_decap_8 FILLER_154_1299 ();
 sg13g2_fill_1 FILLER_154_1306 ();
 sg13g2_decap_4 FILLER_154_1311 ();
 sg13g2_decap_8 FILLER_154_1341 ();
 sg13g2_decap_8 FILLER_154_1348 ();
 sg13g2_decap_8 FILLER_154_1355 ();
 sg13g2_decap_8 FILLER_154_1362 ();
 sg13g2_decap_8 FILLER_154_1369 ();
 sg13g2_decap_8 FILLER_154_1376 ();
 sg13g2_decap_8 FILLER_154_1383 ();
 sg13g2_decap_8 FILLER_154_1390 ();
 sg13g2_decap_8 FILLER_154_1397 ();
 sg13g2_decap_8 FILLER_154_1404 ();
 sg13g2_decap_8 FILLER_154_1411 ();
 sg13g2_decap_8 FILLER_154_1418 ();
 sg13g2_decap_8 FILLER_154_1425 ();
 sg13g2_decap_8 FILLER_154_1432 ();
 sg13g2_decap_8 FILLER_154_1439 ();
 sg13g2_decap_8 FILLER_154_1446 ();
 sg13g2_decap_8 FILLER_154_1453 ();
 sg13g2_decap_8 FILLER_154_1460 ();
 sg13g2_decap_8 FILLER_154_1467 ();
 sg13g2_decap_8 FILLER_154_1474 ();
 sg13g2_decap_8 FILLER_154_1481 ();
 sg13g2_decap_8 FILLER_154_1488 ();
 sg13g2_decap_8 FILLER_154_1495 ();
 sg13g2_decap_8 FILLER_154_1502 ();
 sg13g2_decap_8 FILLER_154_1509 ();
 sg13g2_decap_8 FILLER_154_1516 ();
 sg13g2_decap_8 FILLER_154_1523 ();
 sg13g2_decap_8 FILLER_154_1530 ();
 sg13g2_decap_8 FILLER_154_1537 ();
 sg13g2_decap_8 FILLER_154_1544 ();
 sg13g2_decap_8 FILLER_154_1551 ();
 sg13g2_decap_8 FILLER_154_1558 ();
 sg13g2_decap_8 FILLER_154_1565 ();
 sg13g2_decap_8 FILLER_154_1572 ();
 sg13g2_decap_8 FILLER_154_1579 ();
 sg13g2_decap_8 FILLER_154_1586 ();
 sg13g2_decap_8 FILLER_154_1593 ();
 sg13g2_decap_8 FILLER_154_1600 ();
 sg13g2_decap_8 FILLER_154_1607 ();
 sg13g2_decap_8 FILLER_154_1614 ();
 sg13g2_decap_4 FILLER_154_1621 ();
 sg13g2_decap_8 FILLER_155_0 ();
 sg13g2_fill_2 FILLER_155_7 ();
 sg13g2_fill_2 FILLER_155_34 ();
 sg13g2_decap_4 FILLER_155_66 ();
 sg13g2_fill_2 FILLER_155_70 ();
 sg13g2_decap_8 FILLER_155_82 ();
 sg13g2_decap_8 FILLER_155_114 ();
 sg13g2_fill_2 FILLER_155_132 ();
 sg13g2_fill_1 FILLER_155_134 ();
 sg13g2_decap_8 FILLER_155_169 ();
 sg13g2_decap_4 FILLER_155_176 ();
 sg13g2_fill_1 FILLER_155_180 ();
 sg13g2_fill_1 FILLER_155_189 ();
 sg13g2_decap_4 FILLER_155_193 ();
 sg13g2_fill_2 FILLER_155_248 ();
 sg13g2_fill_1 FILLER_155_250 ();
 sg13g2_decap_8 FILLER_155_255 ();
 sg13g2_decap_8 FILLER_155_262 ();
 sg13g2_decap_8 FILLER_155_269 ();
 sg13g2_fill_1 FILLER_155_276 ();
 sg13g2_fill_1 FILLER_155_315 ();
 sg13g2_fill_2 FILLER_155_322 ();
 sg13g2_fill_1 FILLER_155_324 ();
 sg13g2_decap_8 FILLER_155_337 ();
 sg13g2_decap_8 FILLER_155_344 ();
 sg13g2_decap_8 FILLER_155_351 ();
 sg13g2_fill_2 FILLER_155_383 ();
 sg13g2_fill_1 FILLER_155_390 ();
 sg13g2_fill_1 FILLER_155_396 ();
 sg13g2_decap_8 FILLER_155_423 ();
 sg13g2_decap_4 FILLER_155_430 ();
 sg13g2_fill_2 FILLER_155_434 ();
 sg13g2_fill_2 FILLER_155_440 ();
 sg13g2_fill_1 FILLER_155_442 ();
 sg13g2_decap_8 FILLER_155_499 ();
 sg13g2_decap_4 FILLER_155_506 ();
 sg13g2_fill_2 FILLER_155_510 ();
 sg13g2_fill_2 FILLER_155_529 ();
 sg13g2_decap_4 FILLER_155_561 ();
 sg13g2_decap_4 FILLER_155_617 ();
 sg13g2_decap_8 FILLER_155_657 ();
 sg13g2_fill_2 FILLER_155_664 ();
 sg13g2_fill_1 FILLER_155_670 ();
 sg13g2_fill_2 FILLER_155_675 ();
 sg13g2_decap_8 FILLER_155_710 ();
 sg13g2_decap_4 FILLER_155_717 ();
 sg13g2_decap_8 FILLER_155_725 ();
 sg13g2_decap_8 FILLER_155_732 ();
 sg13g2_decap_8 FILLER_155_739 ();
 sg13g2_decap_8 FILLER_155_746 ();
 sg13g2_decap_8 FILLER_155_753 ();
 sg13g2_decap_8 FILLER_155_760 ();
 sg13g2_decap_8 FILLER_155_767 ();
 sg13g2_decap_8 FILLER_155_774 ();
 sg13g2_decap_8 FILLER_155_781 ();
 sg13g2_decap_4 FILLER_155_788 ();
 sg13g2_fill_1 FILLER_155_792 ();
 sg13g2_fill_2 FILLER_155_796 ();
 sg13g2_fill_1 FILLER_155_798 ();
 sg13g2_decap_8 FILLER_155_825 ();
 sg13g2_decap_8 FILLER_155_832 ();
 sg13g2_decap_8 FILLER_155_839 ();
 sg13g2_decap_8 FILLER_155_846 ();
 sg13g2_decap_8 FILLER_155_853 ();
 sg13g2_decap_8 FILLER_155_860 ();
 sg13g2_decap_8 FILLER_155_867 ();
 sg13g2_decap_4 FILLER_155_874 ();
 sg13g2_fill_1 FILLER_155_878 ();
 sg13g2_decap_4 FILLER_155_885 ();
 sg13g2_fill_2 FILLER_155_889 ();
 sg13g2_decap_4 FILLER_155_897 ();
 sg13g2_fill_1 FILLER_155_901 ();
 sg13g2_decap_8 FILLER_155_934 ();
 sg13g2_decap_4 FILLER_155_941 ();
 sg13g2_decap_8 FILLER_155_949 ();
 sg13g2_decap_8 FILLER_155_956 ();
 sg13g2_fill_2 FILLER_155_963 ();
 sg13g2_fill_1 FILLER_155_965 ();
 sg13g2_decap_4 FILLER_155_1000 ();
 sg13g2_decap_8 FILLER_155_1010 ();
 sg13g2_fill_2 FILLER_155_1017 ();
 sg13g2_fill_1 FILLER_155_1019 ();
 sg13g2_fill_1 FILLER_155_1025 ();
 sg13g2_decap_8 FILLER_155_1056 ();
 sg13g2_decap_8 FILLER_155_1101 ();
 sg13g2_decap_8 FILLER_155_1108 ();
 sg13g2_decap_4 FILLER_155_1115 ();
 sg13g2_fill_2 FILLER_155_1119 ();
 sg13g2_decap_8 FILLER_155_1150 ();
 sg13g2_decap_8 FILLER_155_1157 ();
 sg13g2_fill_2 FILLER_155_1164 ();
 sg13g2_decap_8 FILLER_155_1175 ();
 sg13g2_fill_2 FILLER_155_1182 ();
 sg13g2_fill_1 FILLER_155_1184 ();
 sg13g2_fill_2 FILLER_155_1193 ();
 sg13g2_decap_8 FILLER_155_1199 ();
 sg13g2_decap_4 FILLER_155_1206 ();
 sg13g2_fill_1 FILLER_155_1210 ();
 sg13g2_decap_8 FILLER_155_1214 ();
 sg13g2_decap_8 FILLER_155_1225 ();
 sg13g2_decap_4 FILLER_155_1232 ();
 sg13g2_fill_1 FILLER_155_1236 ();
 sg13g2_decap_8 FILLER_155_1240 ();
 sg13g2_decap_8 FILLER_155_1247 ();
 sg13g2_fill_1 FILLER_155_1254 ();
 sg13g2_decap_8 FILLER_155_1260 ();
 sg13g2_decap_4 FILLER_155_1267 ();
 sg13g2_fill_1 FILLER_155_1289 ();
 sg13g2_fill_1 FILLER_155_1299 ();
 sg13g2_fill_2 FILLER_155_1312 ();
 sg13g2_fill_1 FILLER_155_1314 ();
 sg13g2_decap_8 FILLER_155_1340 ();
 sg13g2_decap_8 FILLER_155_1347 ();
 sg13g2_decap_8 FILLER_155_1354 ();
 sg13g2_decap_8 FILLER_155_1361 ();
 sg13g2_decap_8 FILLER_155_1368 ();
 sg13g2_decap_8 FILLER_155_1375 ();
 sg13g2_decap_8 FILLER_155_1382 ();
 sg13g2_decap_8 FILLER_155_1389 ();
 sg13g2_decap_8 FILLER_155_1396 ();
 sg13g2_decap_8 FILLER_155_1403 ();
 sg13g2_decap_8 FILLER_155_1410 ();
 sg13g2_decap_8 FILLER_155_1417 ();
 sg13g2_decap_8 FILLER_155_1424 ();
 sg13g2_decap_8 FILLER_155_1431 ();
 sg13g2_decap_8 FILLER_155_1438 ();
 sg13g2_decap_8 FILLER_155_1445 ();
 sg13g2_decap_8 FILLER_155_1452 ();
 sg13g2_decap_8 FILLER_155_1459 ();
 sg13g2_decap_8 FILLER_155_1466 ();
 sg13g2_decap_8 FILLER_155_1473 ();
 sg13g2_decap_8 FILLER_155_1480 ();
 sg13g2_decap_8 FILLER_155_1487 ();
 sg13g2_decap_8 FILLER_155_1494 ();
 sg13g2_decap_8 FILLER_155_1501 ();
 sg13g2_decap_8 FILLER_155_1508 ();
 sg13g2_decap_8 FILLER_155_1515 ();
 sg13g2_decap_8 FILLER_155_1522 ();
 sg13g2_decap_8 FILLER_155_1529 ();
 sg13g2_decap_8 FILLER_155_1536 ();
 sg13g2_decap_8 FILLER_155_1543 ();
 sg13g2_decap_8 FILLER_155_1550 ();
 sg13g2_decap_8 FILLER_155_1557 ();
 sg13g2_decap_8 FILLER_155_1564 ();
 sg13g2_decap_8 FILLER_155_1571 ();
 sg13g2_decap_8 FILLER_155_1578 ();
 sg13g2_decap_8 FILLER_155_1585 ();
 sg13g2_decap_8 FILLER_155_1592 ();
 sg13g2_decap_8 FILLER_155_1599 ();
 sg13g2_decap_8 FILLER_155_1606 ();
 sg13g2_decap_8 FILLER_155_1613 ();
 sg13g2_decap_4 FILLER_155_1620 ();
 sg13g2_fill_1 FILLER_155_1624 ();
 sg13g2_decap_8 FILLER_156_0 ();
 sg13g2_decap_8 FILLER_156_43 ();
 sg13g2_decap_4 FILLER_156_50 ();
 sg13g2_fill_1 FILLER_156_54 ();
 sg13g2_decap_8 FILLER_156_60 ();
 sg13g2_decap_8 FILLER_156_72 ();
 sg13g2_fill_2 FILLER_156_79 ();
 sg13g2_fill_1 FILLER_156_112 ();
 sg13g2_decap_4 FILLER_156_117 ();
 sg13g2_fill_2 FILLER_156_121 ();
 sg13g2_fill_1 FILLER_156_128 ();
 sg13g2_fill_1 FILLER_156_144 ();
 sg13g2_decap_8 FILLER_156_200 ();
 sg13g2_fill_2 FILLER_156_207 ();
 sg13g2_fill_2 FILLER_156_297 ();
 sg13g2_decap_8 FILLER_156_329 ();
 sg13g2_decap_4 FILLER_156_336 ();
 sg13g2_fill_2 FILLER_156_340 ();
 sg13g2_decap_8 FILLER_156_346 ();
 sg13g2_decap_4 FILLER_156_353 ();
 sg13g2_fill_1 FILLER_156_357 ();
 sg13g2_fill_2 FILLER_156_361 ();
 sg13g2_fill_1 FILLER_156_363 ();
 sg13g2_fill_1 FILLER_156_367 ();
 sg13g2_decap_4 FILLER_156_416 ();
 sg13g2_fill_1 FILLER_156_420 ();
 sg13g2_decap_8 FILLER_156_455 ();
 sg13g2_decap_4 FILLER_156_462 ();
 sg13g2_fill_1 FILLER_156_466 ();
 sg13g2_fill_2 FILLER_156_483 ();
 sg13g2_fill_1 FILLER_156_485 ();
 sg13g2_decap_8 FILLER_156_496 ();
 sg13g2_decap_4 FILLER_156_503 ();
 sg13g2_fill_2 FILLER_156_541 ();
 sg13g2_fill_2 FILLER_156_547 ();
 sg13g2_fill_2 FILLER_156_558 ();
 sg13g2_fill_1 FILLER_156_560 ();
 sg13g2_decap_8 FILLER_156_565 ();
 sg13g2_decap_8 FILLER_156_572 ();
 sg13g2_decap_4 FILLER_156_579 ();
 sg13g2_decap_8 FILLER_156_612 ();
 sg13g2_decap_8 FILLER_156_619 ();
 sg13g2_decap_8 FILLER_156_626 ();
 sg13g2_fill_2 FILLER_156_637 ();
 sg13g2_fill_1 FILLER_156_639 ();
 sg13g2_decap_4 FILLER_156_645 ();
 sg13g2_fill_1 FILLER_156_649 ();
 sg13g2_fill_2 FILLER_156_660 ();
 sg13g2_fill_1 FILLER_156_662 ();
 sg13g2_fill_1 FILLER_156_693 ();
 sg13g2_decap_8 FILLER_156_699 ();
 sg13g2_fill_1 FILLER_156_706 ();
 sg13g2_fill_2 FILLER_156_711 ();
 sg13g2_fill_1 FILLER_156_713 ();
 sg13g2_decap_4 FILLER_156_740 ();
 sg13g2_fill_2 FILLER_156_744 ();
 sg13g2_decap_8 FILLER_156_750 ();
 sg13g2_decap_8 FILLER_156_757 ();
 sg13g2_decap_4 FILLER_156_764 ();
 sg13g2_decap_8 FILLER_156_782 ();
 sg13g2_decap_8 FILLER_156_818 ();
 sg13g2_decap_8 FILLER_156_825 ();
 sg13g2_decap_4 FILLER_156_832 ();
 sg13g2_fill_2 FILLER_156_836 ();
 sg13g2_decap_8 FILLER_156_857 ();
 sg13g2_fill_2 FILLER_156_882 ();
 sg13g2_fill_1 FILLER_156_893 ();
 sg13g2_fill_2 FILLER_156_936 ();
 sg13g2_decap_8 FILLER_156_964 ();
 sg13g2_decap_4 FILLER_156_971 ();
 sg13g2_fill_1 FILLER_156_975 ();
 sg13g2_decap_8 FILLER_156_981 ();
 sg13g2_decap_8 FILLER_156_988 ();
 sg13g2_decap_4 FILLER_156_995 ();
 sg13g2_fill_1 FILLER_156_999 ();
 sg13g2_fill_1 FILLER_156_1009 ();
 sg13g2_decap_8 FILLER_156_1025 ();
 sg13g2_fill_2 FILLER_156_1032 ();
 sg13g2_fill_1 FILLER_156_1034 ();
 sg13g2_fill_1 FILLER_156_1038 ();
 sg13g2_decap_8 FILLER_156_1046 ();
 sg13g2_decap_8 FILLER_156_1053 ();
 sg13g2_decap_8 FILLER_156_1060 ();
 sg13g2_decap_4 FILLER_156_1098 ();
 sg13g2_fill_2 FILLER_156_1102 ();
 sg13g2_decap_8 FILLER_156_1108 ();
 sg13g2_decap_4 FILLER_156_1127 ();
 sg13g2_fill_1 FILLER_156_1131 ();
 sg13g2_decap_4 FILLER_156_1183 ();
 sg13g2_fill_1 FILLER_156_1187 ();
 sg13g2_decap_8 FILLER_156_1227 ();
 sg13g2_decap_8 FILLER_156_1238 ();
 sg13g2_decap_8 FILLER_156_1245 ();
 sg13g2_decap_8 FILLER_156_1252 ();
 sg13g2_decap_4 FILLER_156_1259 ();
 sg13g2_fill_1 FILLER_156_1277 ();
 sg13g2_decap_8 FILLER_156_1282 ();
 sg13g2_decap_8 FILLER_156_1289 ();
 sg13g2_fill_2 FILLER_156_1296 ();
 sg13g2_fill_1 FILLER_156_1298 ();
 sg13g2_fill_1 FILLER_156_1307 ();
 sg13g2_decap_8 FILLER_156_1334 ();
 sg13g2_decap_8 FILLER_156_1341 ();
 sg13g2_decap_8 FILLER_156_1348 ();
 sg13g2_decap_8 FILLER_156_1355 ();
 sg13g2_decap_8 FILLER_156_1362 ();
 sg13g2_decap_8 FILLER_156_1369 ();
 sg13g2_decap_8 FILLER_156_1376 ();
 sg13g2_decap_8 FILLER_156_1383 ();
 sg13g2_decap_8 FILLER_156_1390 ();
 sg13g2_decap_8 FILLER_156_1397 ();
 sg13g2_decap_8 FILLER_156_1404 ();
 sg13g2_decap_8 FILLER_156_1411 ();
 sg13g2_decap_8 FILLER_156_1418 ();
 sg13g2_decap_8 FILLER_156_1425 ();
 sg13g2_decap_8 FILLER_156_1432 ();
 sg13g2_decap_8 FILLER_156_1439 ();
 sg13g2_decap_8 FILLER_156_1446 ();
 sg13g2_decap_8 FILLER_156_1453 ();
 sg13g2_decap_8 FILLER_156_1460 ();
 sg13g2_decap_8 FILLER_156_1467 ();
 sg13g2_decap_8 FILLER_156_1474 ();
 sg13g2_decap_8 FILLER_156_1481 ();
 sg13g2_decap_8 FILLER_156_1488 ();
 sg13g2_decap_8 FILLER_156_1495 ();
 sg13g2_decap_8 FILLER_156_1502 ();
 sg13g2_decap_8 FILLER_156_1509 ();
 sg13g2_decap_8 FILLER_156_1516 ();
 sg13g2_decap_8 FILLER_156_1523 ();
 sg13g2_decap_8 FILLER_156_1530 ();
 sg13g2_decap_8 FILLER_156_1537 ();
 sg13g2_decap_8 FILLER_156_1544 ();
 sg13g2_decap_8 FILLER_156_1551 ();
 sg13g2_decap_8 FILLER_156_1558 ();
 sg13g2_decap_8 FILLER_156_1565 ();
 sg13g2_decap_8 FILLER_156_1572 ();
 sg13g2_decap_8 FILLER_156_1579 ();
 sg13g2_decap_8 FILLER_156_1586 ();
 sg13g2_decap_8 FILLER_156_1593 ();
 sg13g2_decap_8 FILLER_156_1600 ();
 sg13g2_decap_8 FILLER_156_1607 ();
 sg13g2_decap_8 FILLER_156_1614 ();
 sg13g2_decap_4 FILLER_156_1621 ();
 sg13g2_decap_8 FILLER_157_0 ();
 sg13g2_decap_8 FILLER_157_7 ();
 sg13g2_decap_8 FILLER_157_14 ();
 sg13g2_decap_4 FILLER_157_26 ();
 sg13g2_fill_1 FILLER_157_30 ();
 sg13g2_decap_8 FILLER_157_35 ();
 sg13g2_decap_4 FILLER_157_42 ();
 sg13g2_decap_8 FILLER_157_49 ();
 sg13g2_decap_8 FILLER_157_56 ();
 sg13g2_decap_8 FILLER_157_63 ();
 sg13g2_decap_8 FILLER_157_70 ();
 sg13g2_decap_8 FILLER_157_77 ();
 sg13g2_decap_4 FILLER_157_84 ();
 sg13g2_fill_1 FILLER_157_88 ();
 sg13g2_decap_8 FILLER_157_93 ();
 sg13g2_decap_8 FILLER_157_100 ();
 sg13g2_decap_8 FILLER_157_107 ();
 sg13g2_fill_1 FILLER_157_114 ();
 sg13g2_fill_2 FILLER_157_120 ();
 sg13g2_fill_2 FILLER_157_127 ();
 sg13g2_fill_1 FILLER_157_129 ();
 sg13g2_fill_2 FILLER_157_134 ();
 sg13g2_fill_1 FILLER_157_151 ();
 sg13g2_decap_8 FILLER_157_178 ();
 sg13g2_decap_4 FILLER_157_185 ();
 sg13g2_fill_1 FILLER_157_189 ();
 sg13g2_fill_2 FILLER_157_215 ();
 sg13g2_decap_8 FILLER_157_221 ();
 sg13g2_fill_2 FILLER_157_238 ();
 sg13g2_fill_2 FILLER_157_245 ();
 sg13g2_fill_1 FILLER_157_247 ();
 sg13g2_decap_4 FILLER_157_280 ();
 sg13g2_fill_1 FILLER_157_284 ();
 sg13g2_decap_8 FILLER_157_289 ();
 sg13g2_decap_4 FILLER_157_296 ();
 sg13g2_fill_1 FILLER_157_300 ();
 sg13g2_decap_8 FILLER_157_306 ();
 sg13g2_decap_8 FILLER_157_313 ();
 sg13g2_fill_2 FILLER_157_320 ();
 sg13g2_fill_1 FILLER_157_322 ();
 sg13g2_fill_2 FILLER_157_326 ();
 sg13g2_fill_1 FILLER_157_328 ();
 sg13g2_fill_1 FILLER_157_333 ();
 sg13g2_fill_2 FILLER_157_360 ();
 sg13g2_decap_8 FILLER_157_437 ();
 sg13g2_decap_4 FILLER_157_444 ();
 sg13g2_fill_1 FILLER_157_448 ();
 sg13g2_decap_8 FILLER_157_492 ();
 sg13g2_decap_8 FILLER_157_503 ();
 sg13g2_decap_8 FILLER_157_536 ();
 sg13g2_fill_2 FILLER_157_586 ();
 sg13g2_fill_1 FILLER_157_588 ();
 sg13g2_decap_4 FILLER_157_620 ();
 sg13g2_fill_1 FILLER_157_624 ();
 sg13g2_decap_8 FILLER_157_653 ();
 sg13g2_fill_2 FILLER_157_686 ();
 sg13g2_fill_1 FILLER_157_688 ();
 sg13g2_decap_4 FILLER_157_695 ();
 sg13g2_fill_2 FILLER_157_735 ();
 sg13g2_fill_2 FILLER_157_767 ();
 sg13g2_fill_1 FILLER_157_795 ();
 sg13g2_fill_1 FILLER_157_822 ();
 sg13g2_fill_1 FILLER_157_828 ();
 sg13g2_fill_1 FILLER_157_833 ();
 sg13g2_fill_2 FILLER_157_840 ();
 sg13g2_decap_4 FILLER_157_865 ();
 sg13g2_fill_2 FILLER_157_869 ();
 sg13g2_decap_4 FILLER_157_876 ();
 sg13g2_fill_1 FILLER_157_880 ();
 sg13g2_decap_8 FILLER_157_894 ();
 sg13g2_decap_8 FILLER_157_901 ();
 sg13g2_decap_8 FILLER_157_908 ();
 sg13g2_decap_8 FILLER_157_915 ();
 sg13g2_decap_8 FILLER_157_922 ();
 sg13g2_fill_2 FILLER_157_929 ();
 sg13g2_decap_8 FILLER_157_939 ();
 sg13g2_fill_2 FILLER_157_983 ();
 sg13g2_fill_1 FILLER_157_985 ();
 sg13g2_decap_8 FILLER_157_990 ();
 sg13g2_decap_8 FILLER_157_997 ();
 sg13g2_decap_8 FILLER_157_1004 ();
 sg13g2_decap_8 FILLER_157_1011 ();
 sg13g2_fill_2 FILLER_157_1018 ();
 sg13g2_fill_1 FILLER_157_1020 ();
 sg13g2_decap_4 FILLER_157_1027 ();
 sg13g2_fill_2 FILLER_157_1031 ();
 sg13g2_decap_4 FILLER_157_1039 ();
 sg13g2_fill_1 FILLER_157_1043 ();
 sg13g2_decap_8 FILLER_157_1048 ();
 sg13g2_decap_8 FILLER_157_1067 ();
 sg13g2_decap_8 FILLER_157_1074 ();
 sg13g2_decap_8 FILLER_157_1081 ();
 sg13g2_fill_2 FILLER_157_1094 ();
 sg13g2_fill_2 FILLER_157_1127 ();
 sg13g2_fill_1 FILLER_157_1129 ();
 sg13g2_fill_1 FILLER_157_1156 ();
 sg13g2_decap_4 FILLER_157_1187 ();
 sg13g2_fill_2 FILLER_157_1191 ();
 sg13g2_decap_8 FILLER_157_1197 ();
 sg13g2_decap_8 FILLER_157_1204 ();
 sg13g2_fill_1 FILLER_157_1224 ();
 sg13g2_decap_8 FILLER_157_1251 ();
 sg13g2_decap_8 FILLER_157_1258 ();
 sg13g2_decap_4 FILLER_157_1265 ();
 sg13g2_decap_4 FILLER_157_1274 ();
 sg13g2_decap_8 FILLER_157_1282 ();
 sg13g2_decap_4 FILLER_157_1289 ();
 sg13g2_fill_2 FILLER_157_1305 ();
 sg13g2_decap_4 FILLER_157_1311 ();
 sg13g2_decap_8 FILLER_157_1319 ();
 sg13g2_decap_8 FILLER_157_1326 ();
 sg13g2_decap_8 FILLER_157_1333 ();
 sg13g2_decap_8 FILLER_157_1340 ();
 sg13g2_decap_8 FILLER_157_1347 ();
 sg13g2_decap_8 FILLER_157_1354 ();
 sg13g2_decap_8 FILLER_157_1361 ();
 sg13g2_decap_8 FILLER_157_1368 ();
 sg13g2_decap_8 FILLER_157_1375 ();
 sg13g2_decap_8 FILLER_157_1382 ();
 sg13g2_decap_8 FILLER_157_1389 ();
 sg13g2_decap_8 FILLER_157_1396 ();
 sg13g2_decap_8 FILLER_157_1403 ();
 sg13g2_decap_8 FILLER_157_1410 ();
 sg13g2_decap_8 FILLER_157_1417 ();
 sg13g2_decap_8 FILLER_157_1424 ();
 sg13g2_decap_8 FILLER_157_1431 ();
 sg13g2_decap_8 FILLER_157_1438 ();
 sg13g2_decap_8 FILLER_157_1445 ();
 sg13g2_decap_8 FILLER_157_1452 ();
 sg13g2_decap_8 FILLER_157_1459 ();
 sg13g2_decap_8 FILLER_157_1466 ();
 sg13g2_decap_8 FILLER_157_1473 ();
 sg13g2_decap_8 FILLER_157_1480 ();
 sg13g2_decap_8 FILLER_157_1487 ();
 sg13g2_decap_8 FILLER_157_1494 ();
 sg13g2_decap_8 FILLER_157_1501 ();
 sg13g2_decap_8 FILLER_157_1508 ();
 sg13g2_decap_8 FILLER_157_1515 ();
 sg13g2_decap_8 FILLER_157_1522 ();
 sg13g2_decap_8 FILLER_157_1529 ();
 sg13g2_decap_8 FILLER_157_1536 ();
 sg13g2_decap_8 FILLER_157_1543 ();
 sg13g2_decap_8 FILLER_157_1550 ();
 sg13g2_decap_8 FILLER_157_1557 ();
 sg13g2_decap_8 FILLER_157_1564 ();
 sg13g2_decap_8 FILLER_157_1571 ();
 sg13g2_decap_8 FILLER_157_1578 ();
 sg13g2_decap_8 FILLER_157_1585 ();
 sg13g2_decap_8 FILLER_157_1592 ();
 sg13g2_decap_8 FILLER_157_1599 ();
 sg13g2_decap_8 FILLER_157_1606 ();
 sg13g2_decap_8 FILLER_157_1613 ();
 sg13g2_decap_4 FILLER_157_1620 ();
 sg13g2_fill_1 FILLER_157_1624 ();
 sg13g2_decap_8 FILLER_158_0 ();
 sg13g2_decap_8 FILLER_158_7 ();
 sg13g2_decap_8 FILLER_158_14 ();
 sg13g2_decap_4 FILLER_158_55 ();
 sg13g2_fill_1 FILLER_158_59 ();
 sg13g2_decap_8 FILLER_158_65 ();
 sg13g2_decap_4 FILLER_158_86 ();
 sg13g2_fill_1 FILLER_158_90 ();
 sg13g2_decap_8 FILLER_158_95 ();
 sg13g2_decap_8 FILLER_158_102 ();
 sg13g2_decap_4 FILLER_158_119 ();
 sg13g2_fill_2 FILLER_158_136 ();
 sg13g2_fill_1 FILLER_158_138 ();
 sg13g2_decap_8 FILLER_158_165 ();
 sg13g2_decap_8 FILLER_158_172 ();
 sg13g2_decap_8 FILLER_158_179 ();
 sg13g2_decap_8 FILLER_158_186 ();
 sg13g2_decap_8 FILLER_158_193 ();
 sg13g2_decap_4 FILLER_158_200 ();
 sg13g2_fill_1 FILLER_158_204 ();
 sg13g2_decap_8 FILLER_158_219 ();
 sg13g2_fill_2 FILLER_158_226 ();
 sg13g2_fill_1 FILLER_158_228 ();
 sg13g2_decap_8 FILLER_158_234 ();
 sg13g2_decap_8 FILLER_158_241 ();
 sg13g2_decap_8 FILLER_158_248 ();
 sg13g2_fill_1 FILLER_158_255 ();
 sg13g2_decap_8 FILLER_158_282 ();
 sg13g2_decap_8 FILLER_158_289 ();
 sg13g2_fill_2 FILLER_158_296 ();
 sg13g2_fill_1 FILLER_158_298 ();
 sg13g2_decap_8 FILLER_158_348 ();
 sg13g2_decap_4 FILLER_158_355 ();
 sg13g2_fill_1 FILLER_158_359 ();
 sg13g2_fill_2 FILLER_158_374 ();
 sg13g2_fill_2 FILLER_158_433 ();
 sg13g2_fill_1 FILLER_158_435 ();
 sg13g2_fill_1 FILLER_158_502 ();
 sg13g2_fill_2 FILLER_158_513 ();
 sg13g2_fill_2 FILLER_158_519 ();
 sg13g2_fill_1 FILLER_158_521 ();
 sg13g2_fill_1 FILLER_158_526 ();
 sg13g2_fill_2 FILLER_158_532 ();
 sg13g2_decap_4 FILLER_158_540 ();
 sg13g2_decap_8 FILLER_158_574 ();
 sg13g2_fill_1 FILLER_158_581 ();
 sg13g2_decap_8 FILLER_158_614 ();
 sg13g2_decap_8 FILLER_158_651 ();
 sg13g2_decap_8 FILLER_158_658 ();
 sg13g2_decap_8 FILLER_158_665 ();
 sg13g2_decap_8 FILLER_158_672 ();
 sg13g2_fill_2 FILLER_158_679 ();
 sg13g2_fill_2 FILLER_158_718 ();
 sg13g2_decap_8 FILLER_158_780 ();
 sg13g2_fill_1 FILLER_158_812 ();
 sg13g2_decap_4 FILLER_158_842 ();
 sg13g2_fill_1 FILLER_158_846 ();
 sg13g2_decap_8 FILLER_158_880 ();
 sg13g2_decap_8 FILLER_158_887 ();
 sg13g2_decap_4 FILLER_158_894 ();
 sg13g2_fill_1 FILLER_158_898 ();
 sg13g2_fill_2 FILLER_158_939 ();
 sg13g2_fill_1 FILLER_158_941 ();
 sg13g2_fill_1 FILLER_158_947 ();
 sg13g2_decap_4 FILLER_158_974 ();
 sg13g2_fill_1 FILLER_158_1004 ();
 sg13g2_decap_4 FILLER_158_1016 ();
 sg13g2_fill_1 FILLER_158_1020 ();
 sg13g2_decap_8 FILLER_158_1025 ();
 sg13g2_decap_4 FILLER_158_1062 ();
 sg13g2_fill_1 FILLER_158_1066 ();
 sg13g2_fill_2 FILLER_158_1072 ();
 sg13g2_fill_1 FILLER_158_1074 ();
 sg13g2_decap_8 FILLER_158_1079 ();
 sg13g2_decap_8 FILLER_158_1092 ();
 sg13g2_decap_8 FILLER_158_1099 ();
 sg13g2_fill_2 FILLER_158_1106 ();
 sg13g2_decap_8 FILLER_158_1154 ();
 sg13g2_decap_8 FILLER_158_1161 ();
 sg13g2_decap_4 FILLER_158_1168 ();
 sg13g2_decap_8 FILLER_158_1180 ();
 sg13g2_decap_8 FILLER_158_1205 ();
 sg13g2_decap_8 FILLER_158_1217 ();
 sg13g2_decap_8 FILLER_158_1224 ();
 sg13g2_decap_4 FILLER_158_1231 ();
 sg13g2_fill_1 FILLER_158_1235 ();
 sg13g2_fill_2 FILLER_158_1249 ();
 sg13g2_fill_1 FILLER_158_1251 ();
 sg13g2_fill_1 FILLER_158_1266 ();
 sg13g2_decap_8 FILLER_158_1271 ();
 sg13g2_decap_4 FILLER_158_1278 ();
 sg13g2_decap_8 FILLER_158_1298 ();
 sg13g2_fill_1 FILLER_158_1305 ();
 sg13g2_decap_8 FILLER_158_1332 ();
 sg13g2_decap_8 FILLER_158_1339 ();
 sg13g2_decap_8 FILLER_158_1346 ();
 sg13g2_decap_8 FILLER_158_1353 ();
 sg13g2_decap_8 FILLER_158_1360 ();
 sg13g2_decap_8 FILLER_158_1367 ();
 sg13g2_decap_8 FILLER_158_1374 ();
 sg13g2_decap_8 FILLER_158_1381 ();
 sg13g2_decap_8 FILLER_158_1388 ();
 sg13g2_decap_8 FILLER_158_1395 ();
 sg13g2_decap_8 FILLER_158_1402 ();
 sg13g2_decap_8 FILLER_158_1409 ();
 sg13g2_decap_8 FILLER_158_1416 ();
 sg13g2_decap_8 FILLER_158_1423 ();
 sg13g2_decap_8 FILLER_158_1430 ();
 sg13g2_decap_8 FILLER_158_1437 ();
 sg13g2_decap_8 FILLER_158_1444 ();
 sg13g2_decap_8 FILLER_158_1451 ();
 sg13g2_decap_8 FILLER_158_1458 ();
 sg13g2_decap_8 FILLER_158_1465 ();
 sg13g2_decap_8 FILLER_158_1472 ();
 sg13g2_decap_8 FILLER_158_1479 ();
 sg13g2_decap_8 FILLER_158_1486 ();
 sg13g2_decap_8 FILLER_158_1493 ();
 sg13g2_decap_8 FILLER_158_1500 ();
 sg13g2_decap_8 FILLER_158_1507 ();
 sg13g2_decap_8 FILLER_158_1514 ();
 sg13g2_decap_8 FILLER_158_1521 ();
 sg13g2_decap_8 FILLER_158_1528 ();
 sg13g2_decap_8 FILLER_158_1535 ();
 sg13g2_decap_8 FILLER_158_1542 ();
 sg13g2_decap_8 FILLER_158_1549 ();
 sg13g2_decap_8 FILLER_158_1556 ();
 sg13g2_decap_8 FILLER_158_1563 ();
 sg13g2_decap_8 FILLER_158_1570 ();
 sg13g2_decap_8 FILLER_158_1577 ();
 sg13g2_decap_8 FILLER_158_1584 ();
 sg13g2_decap_8 FILLER_158_1591 ();
 sg13g2_decap_8 FILLER_158_1598 ();
 sg13g2_decap_8 FILLER_158_1605 ();
 sg13g2_decap_8 FILLER_158_1612 ();
 sg13g2_decap_4 FILLER_158_1619 ();
 sg13g2_fill_2 FILLER_158_1623 ();
 sg13g2_decap_8 FILLER_159_0 ();
 sg13g2_decap_8 FILLER_159_7 ();
 sg13g2_decap_8 FILLER_159_14 ();
 sg13g2_decap_8 FILLER_159_21 ();
 sg13g2_decap_4 FILLER_159_28 ();
 sg13g2_fill_2 FILLER_159_32 ();
 sg13g2_decap_4 FILLER_159_70 ();
 sg13g2_fill_1 FILLER_159_74 ();
 sg13g2_decap_8 FILLER_159_127 ();
 sg13g2_decap_8 FILLER_159_134 ();
 sg13g2_fill_1 FILLER_159_141 ();
 sg13g2_decap_8 FILLER_159_146 ();
 sg13g2_decap_8 FILLER_159_153 ();
 sg13g2_decap_8 FILLER_159_160 ();
 sg13g2_decap_8 FILLER_159_167 ();
 sg13g2_decap_8 FILLER_159_174 ();
 sg13g2_decap_8 FILLER_159_181 ();
 sg13g2_decap_8 FILLER_159_188 ();
 sg13g2_decap_8 FILLER_159_195 ();
 sg13g2_decap_8 FILLER_159_202 ();
 sg13g2_decap_8 FILLER_159_209 ();
 sg13g2_decap_8 FILLER_159_216 ();
 sg13g2_decap_8 FILLER_159_223 ();
 sg13g2_decap_8 FILLER_159_256 ();
 sg13g2_decap_8 FILLER_159_263 ();
 sg13g2_decap_8 FILLER_159_270 ();
 sg13g2_fill_2 FILLER_159_277 ();
 sg13g2_fill_1 FILLER_159_279 ();
 sg13g2_decap_8 FILLER_159_284 ();
 sg13g2_decap_8 FILLER_159_291 ();
 sg13g2_fill_1 FILLER_159_298 ();
 sg13g2_fill_1 FILLER_159_305 ();
 sg13g2_decap_8 FILLER_159_312 ();
 sg13g2_fill_2 FILLER_159_324 ();
 sg13g2_fill_1 FILLER_159_326 ();
 sg13g2_fill_2 FILLER_159_336 ();
 sg13g2_fill_1 FILLER_159_338 ();
 sg13g2_decap_8 FILLER_159_343 ();
 sg13g2_decap_8 FILLER_159_350 ();
 sg13g2_decap_4 FILLER_159_357 ();
 sg13g2_fill_1 FILLER_159_489 ();
 sg13g2_fill_2 FILLER_159_516 ();
 sg13g2_decap_4 FILLER_159_532 ();
 sg13g2_decap_8 FILLER_159_546 ();
 sg13g2_decap_4 FILLER_159_565 ();
 sg13g2_fill_2 FILLER_159_605 ();
 sg13g2_decap_8 FILLER_159_613 ();
 sg13g2_decap_8 FILLER_159_620 ();
 sg13g2_fill_2 FILLER_159_627 ();
 sg13g2_decap_4 FILLER_159_640 ();
 sg13g2_fill_1 FILLER_159_644 ();
 sg13g2_fill_2 FILLER_159_655 ();
 sg13g2_fill_1 FILLER_159_657 ();
 sg13g2_fill_2 FILLER_159_662 ();
 sg13g2_fill_1 FILLER_159_664 ();
 sg13g2_fill_1 FILLER_159_676 ();
 sg13g2_fill_1 FILLER_159_714 ();
 sg13g2_fill_2 FILLER_159_725 ();
 sg13g2_fill_2 FILLER_159_778 ();
 sg13g2_fill_1 FILLER_159_780 ();
 sg13g2_decap_4 FILLER_159_785 ();
 sg13g2_fill_2 FILLER_159_789 ();
 sg13g2_fill_2 FILLER_159_801 ();
 sg13g2_decap_8 FILLER_159_807 ();
 sg13g2_decap_4 FILLER_159_814 ();
 sg13g2_fill_2 FILLER_159_818 ();
 sg13g2_decap_8 FILLER_159_844 ();
 sg13g2_decap_8 FILLER_159_851 ();
 sg13g2_decap_8 FILLER_159_858 ();
 sg13g2_decap_8 FILLER_159_865 ();
 sg13g2_decap_8 FILLER_159_872 ();
 sg13g2_decap_4 FILLER_159_879 ();
 sg13g2_fill_2 FILLER_159_883 ();
 sg13g2_decap_4 FILLER_159_894 ();
 sg13g2_fill_1 FILLER_159_898 ();
 sg13g2_fill_1 FILLER_159_904 ();
 sg13g2_fill_2 FILLER_159_909 ();
 sg13g2_fill_1 FILLER_159_911 ();
 sg13g2_fill_1 FILLER_159_937 ();
 sg13g2_decap_4 FILLER_159_955 ();
 sg13g2_fill_2 FILLER_159_959 ();
 sg13g2_decap_4 FILLER_159_969 ();
 sg13g2_decap_4 FILLER_159_977 ();
 sg13g2_fill_1 FILLER_159_981 ();
 sg13g2_decap_8 FILLER_159_988 ();
 sg13g2_decap_4 FILLER_159_995 ();
 sg13g2_fill_1 FILLER_159_999 ();
 sg13g2_decap_4 FILLER_159_1004 ();
 sg13g2_fill_1 FILLER_159_1008 ();
 sg13g2_decap_8 FILLER_159_1014 ();
 sg13g2_decap_4 FILLER_159_1027 ();
 sg13g2_fill_2 FILLER_159_1031 ();
 sg13g2_decap_8 FILLER_159_1039 ();
 sg13g2_decap_8 FILLER_159_1046 ();
 sg13g2_decap_8 FILLER_159_1053 ();
 sg13g2_fill_2 FILLER_159_1086 ();
 sg13g2_fill_1 FILLER_159_1088 ();
 sg13g2_decap_4 FILLER_159_1093 ();
 sg13g2_fill_1 FILLER_159_1097 ();
 sg13g2_decap_8 FILLER_159_1102 ();
 sg13g2_fill_1 FILLER_159_1109 ();
 sg13g2_decap_4 FILLER_159_1115 ();
 sg13g2_fill_1 FILLER_159_1145 ();
 sg13g2_decap_4 FILLER_159_1150 ();
 sg13g2_fill_2 FILLER_159_1158 ();
 sg13g2_fill_2 FILLER_159_1177 ();
 sg13g2_decap_4 FILLER_159_1192 ();
 sg13g2_fill_2 FILLER_159_1196 ();
 sg13g2_decap_4 FILLER_159_1207 ();
 sg13g2_fill_2 FILLER_159_1211 ();
 sg13g2_fill_1 FILLER_159_1218 ();
 sg13g2_decap_8 FILLER_159_1227 ();
 sg13g2_fill_2 FILLER_159_1259 ();
 sg13g2_fill_1 FILLER_159_1261 ();
 sg13g2_decap_4 FILLER_159_1270 ();
 sg13g2_fill_1 FILLER_159_1274 ();
 sg13g2_decap_8 FILLER_159_1279 ();
 sg13g2_decap_8 FILLER_159_1286 ();
 sg13g2_decap_8 FILLER_159_1293 ();
 sg13g2_decap_8 FILLER_159_1300 ();
 sg13g2_decap_8 FILLER_159_1307 ();
 sg13g2_decap_8 FILLER_159_1318 ();
 sg13g2_decap_8 FILLER_159_1325 ();
 sg13g2_decap_8 FILLER_159_1332 ();
 sg13g2_decap_8 FILLER_159_1339 ();
 sg13g2_decap_8 FILLER_159_1346 ();
 sg13g2_decap_8 FILLER_159_1353 ();
 sg13g2_decap_8 FILLER_159_1360 ();
 sg13g2_decap_8 FILLER_159_1367 ();
 sg13g2_decap_8 FILLER_159_1374 ();
 sg13g2_decap_8 FILLER_159_1381 ();
 sg13g2_decap_8 FILLER_159_1388 ();
 sg13g2_decap_8 FILLER_159_1395 ();
 sg13g2_decap_8 FILLER_159_1402 ();
 sg13g2_decap_8 FILLER_159_1409 ();
 sg13g2_decap_8 FILLER_159_1416 ();
 sg13g2_decap_8 FILLER_159_1423 ();
 sg13g2_decap_8 FILLER_159_1430 ();
 sg13g2_decap_8 FILLER_159_1437 ();
 sg13g2_decap_8 FILLER_159_1444 ();
 sg13g2_decap_8 FILLER_159_1451 ();
 sg13g2_decap_8 FILLER_159_1458 ();
 sg13g2_decap_8 FILLER_159_1465 ();
 sg13g2_decap_8 FILLER_159_1472 ();
 sg13g2_decap_8 FILLER_159_1479 ();
 sg13g2_decap_8 FILLER_159_1486 ();
 sg13g2_decap_8 FILLER_159_1493 ();
 sg13g2_decap_8 FILLER_159_1500 ();
 sg13g2_decap_8 FILLER_159_1507 ();
 sg13g2_decap_8 FILLER_159_1514 ();
 sg13g2_decap_8 FILLER_159_1521 ();
 sg13g2_decap_8 FILLER_159_1528 ();
 sg13g2_decap_8 FILLER_159_1535 ();
 sg13g2_decap_8 FILLER_159_1542 ();
 sg13g2_decap_8 FILLER_159_1549 ();
 sg13g2_decap_8 FILLER_159_1556 ();
 sg13g2_decap_8 FILLER_159_1563 ();
 sg13g2_decap_8 FILLER_159_1570 ();
 sg13g2_decap_8 FILLER_159_1577 ();
 sg13g2_decap_8 FILLER_159_1584 ();
 sg13g2_decap_8 FILLER_159_1591 ();
 sg13g2_decap_8 FILLER_159_1598 ();
 sg13g2_decap_8 FILLER_159_1605 ();
 sg13g2_decap_8 FILLER_159_1612 ();
 sg13g2_decap_4 FILLER_159_1619 ();
 sg13g2_fill_2 FILLER_159_1623 ();
 sg13g2_decap_8 FILLER_160_0 ();
 sg13g2_decap_8 FILLER_160_7 ();
 sg13g2_decap_8 FILLER_160_14 ();
 sg13g2_decap_8 FILLER_160_21 ();
 sg13g2_decap_8 FILLER_160_28 ();
 sg13g2_fill_2 FILLER_160_35 ();
 sg13g2_fill_1 FILLER_160_37 ();
 sg13g2_decap_8 FILLER_160_77 ();
 sg13g2_decap_8 FILLER_160_84 ();
 sg13g2_fill_2 FILLER_160_91 ();
 sg13g2_decap_8 FILLER_160_118 ();
 sg13g2_decap_8 FILLER_160_125 ();
 sg13g2_decap_8 FILLER_160_132 ();
 sg13g2_decap_8 FILLER_160_139 ();
 sg13g2_decap_8 FILLER_160_146 ();
 sg13g2_decap_8 FILLER_160_153 ();
 sg13g2_decap_8 FILLER_160_160 ();
 sg13g2_decap_8 FILLER_160_167 ();
 sg13g2_decap_8 FILLER_160_174 ();
 sg13g2_decap_8 FILLER_160_181 ();
 sg13g2_decap_8 FILLER_160_188 ();
 sg13g2_decap_8 FILLER_160_195 ();
 sg13g2_decap_8 FILLER_160_202 ();
 sg13g2_decap_8 FILLER_160_209 ();
 sg13g2_decap_8 FILLER_160_216 ();
 sg13g2_decap_8 FILLER_160_223 ();
 sg13g2_decap_8 FILLER_160_230 ();
 sg13g2_decap_8 FILLER_160_241 ();
 sg13g2_decap_8 FILLER_160_248 ();
 sg13g2_decap_8 FILLER_160_255 ();
 sg13g2_decap_8 FILLER_160_262 ();
 sg13g2_decap_4 FILLER_160_269 ();
 sg13g2_decap_8 FILLER_160_299 ();
 sg13g2_decap_4 FILLER_160_306 ();
 sg13g2_fill_2 FILLER_160_310 ();
 sg13g2_decap_4 FILLER_160_316 ();
 sg13g2_fill_1 FILLER_160_320 ();
 sg13g2_decap_4 FILLER_160_324 ();
 sg13g2_fill_2 FILLER_160_463 ();
 sg13g2_fill_1 FILLER_160_465 ();
 sg13g2_fill_2 FILLER_160_475 ();
 sg13g2_decap_8 FILLER_160_509 ();
 sg13g2_decap_8 FILLER_160_516 ();
 sg13g2_decap_4 FILLER_160_523 ();
 sg13g2_decap_8 FILLER_160_532 ();
 sg13g2_fill_1 FILLER_160_539 ();
 sg13g2_fill_2 FILLER_160_578 ();
 sg13g2_fill_2 FILLER_160_595 ();
 sg13g2_decap_8 FILLER_160_601 ();
 sg13g2_fill_2 FILLER_160_613 ();
 sg13g2_fill_1 FILLER_160_615 ();
 sg13g2_fill_2 FILLER_160_626 ();
 sg13g2_fill_1 FILLER_160_628 ();
 sg13g2_decap_8 FILLER_160_637 ();
 sg13g2_fill_1 FILLER_160_644 ();
 sg13g2_fill_2 FILLER_160_679 ();
 sg13g2_decap_8 FILLER_160_691 ();
 sg13g2_decap_4 FILLER_160_698 ();
 sg13g2_fill_2 FILLER_160_702 ();
 sg13g2_decap_8 FILLER_160_719 ();
 sg13g2_decap_8 FILLER_160_726 ();
 sg13g2_fill_2 FILLER_160_733 ();
 sg13g2_fill_1 FILLER_160_749 ();
 sg13g2_fill_2 FILLER_160_759 ();
 sg13g2_fill_1 FILLER_160_761 ();
 sg13g2_fill_2 FILLER_160_808 ();
 sg13g2_fill_2 FILLER_160_839 ();
 sg13g2_fill_1 FILLER_160_841 ();
 sg13g2_decap_4 FILLER_160_854 ();
 sg13g2_fill_2 FILLER_160_858 ();
 sg13g2_fill_2 FILLER_160_870 ();
 sg13g2_decap_8 FILLER_160_876 ();
 sg13g2_fill_1 FILLER_160_883 ();
 sg13g2_fill_2 FILLER_160_895 ();
 sg13g2_fill_1 FILLER_160_964 ();
 sg13g2_fill_2 FILLER_160_991 ();
 sg13g2_decap_8 FILLER_160_1019 ();
 sg13g2_decap_4 FILLER_160_1026 ();
 sg13g2_decap_8 FILLER_160_1034 ();
 sg13g2_fill_2 FILLER_160_1041 ();
 sg13g2_fill_1 FILLER_160_1043 ();
 sg13g2_decap_8 FILLER_160_1048 ();
 sg13g2_decap_8 FILLER_160_1055 ();
 sg13g2_decap_4 FILLER_160_1062 ();
 sg13g2_fill_1 FILLER_160_1066 ();
 sg13g2_decap_8 FILLER_160_1071 ();
 sg13g2_decap_8 FILLER_160_1078 ();
 sg13g2_decap_8 FILLER_160_1085 ();
 sg13g2_decap_4 FILLER_160_1118 ();
 sg13g2_fill_2 FILLER_160_1126 ();
 sg13g2_fill_1 FILLER_160_1128 ();
 sg13g2_decap_8 FILLER_160_1132 ();
 sg13g2_decap_8 FILLER_160_1139 ();
 sg13g2_fill_1 FILLER_160_1146 ();
 sg13g2_fill_2 FILLER_160_1173 ();
 sg13g2_fill_1 FILLER_160_1179 ();
 sg13g2_fill_1 FILLER_160_1184 ();
 sg13g2_decap_8 FILLER_160_1194 ();
 sg13g2_decap_8 FILLER_160_1201 ();
 sg13g2_fill_1 FILLER_160_1208 ();
 sg13g2_decap_4 FILLER_160_1226 ();
 sg13g2_fill_2 FILLER_160_1230 ();
 sg13g2_decap_4 FILLER_160_1292 ();
 sg13g2_fill_2 FILLER_160_1296 ();
 sg13g2_decap_8 FILLER_160_1302 ();
 sg13g2_fill_1 FILLER_160_1309 ();
 sg13g2_decap_8 FILLER_160_1314 ();
 sg13g2_decap_8 FILLER_160_1321 ();
 sg13g2_decap_8 FILLER_160_1328 ();
 sg13g2_decap_8 FILLER_160_1335 ();
 sg13g2_decap_8 FILLER_160_1342 ();
 sg13g2_decap_8 FILLER_160_1349 ();
 sg13g2_decap_8 FILLER_160_1356 ();
 sg13g2_decap_8 FILLER_160_1363 ();
 sg13g2_decap_8 FILLER_160_1370 ();
 sg13g2_decap_8 FILLER_160_1377 ();
 sg13g2_decap_8 FILLER_160_1384 ();
 sg13g2_decap_8 FILLER_160_1391 ();
 sg13g2_decap_8 FILLER_160_1398 ();
 sg13g2_decap_8 FILLER_160_1405 ();
 sg13g2_decap_8 FILLER_160_1412 ();
 sg13g2_decap_8 FILLER_160_1419 ();
 sg13g2_decap_8 FILLER_160_1426 ();
 sg13g2_decap_8 FILLER_160_1433 ();
 sg13g2_decap_8 FILLER_160_1440 ();
 sg13g2_decap_8 FILLER_160_1447 ();
 sg13g2_decap_8 FILLER_160_1454 ();
 sg13g2_decap_8 FILLER_160_1461 ();
 sg13g2_decap_8 FILLER_160_1468 ();
 sg13g2_decap_8 FILLER_160_1475 ();
 sg13g2_decap_8 FILLER_160_1482 ();
 sg13g2_decap_8 FILLER_160_1489 ();
 sg13g2_decap_8 FILLER_160_1496 ();
 sg13g2_decap_8 FILLER_160_1503 ();
 sg13g2_decap_8 FILLER_160_1510 ();
 sg13g2_decap_8 FILLER_160_1517 ();
 sg13g2_decap_8 FILLER_160_1524 ();
 sg13g2_decap_8 FILLER_160_1531 ();
 sg13g2_decap_8 FILLER_160_1538 ();
 sg13g2_decap_8 FILLER_160_1545 ();
 sg13g2_decap_8 FILLER_160_1552 ();
 sg13g2_decap_8 FILLER_160_1559 ();
 sg13g2_decap_8 FILLER_160_1566 ();
 sg13g2_decap_8 FILLER_160_1573 ();
 sg13g2_decap_8 FILLER_160_1580 ();
 sg13g2_decap_8 FILLER_160_1587 ();
 sg13g2_decap_8 FILLER_160_1594 ();
 sg13g2_decap_8 FILLER_160_1601 ();
 sg13g2_decap_8 FILLER_160_1608 ();
 sg13g2_decap_8 FILLER_160_1615 ();
 sg13g2_fill_2 FILLER_160_1622 ();
 sg13g2_fill_1 FILLER_160_1624 ();
 sg13g2_decap_8 FILLER_161_0 ();
 sg13g2_decap_8 FILLER_161_7 ();
 sg13g2_decap_4 FILLER_161_44 ();
 sg13g2_decap_8 FILLER_161_77 ();
 sg13g2_decap_8 FILLER_161_84 ();
 sg13g2_decap_8 FILLER_161_91 ();
 sg13g2_decap_8 FILLER_161_98 ();
 sg13g2_fill_2 FILLER_161_105 ();
 sg13g2_fill_1 FILLER_161_107 ();
 sg13g2_decap_8 FILLER_161_112 ();
 sg13g2_decap_8 FILLER_161_119 ();
 sg13g2_decap_8 FILLER_161_126 ();
 sg13g2_decap_8 FILLER_161_133 ();
 sg13g2_decap_8 FILLER_161_140 ();
 sg13g2_decap_8 FILLER_161_147 ();
 sg13g2_decap_8 FILLER_161_154 ();
 sg13g2_decap_8 FILLER_161_161 ();
 sg13g2_decap_8 FILLER_161_168 ();
 sg13g2_decap_8 FILLER_161_175 ();
 sg13g2_decap_8 FILLER_161_182 ();
 sg13g2_decap_8 FILLER_161_189 ();
 sg13g2_decap_8 FILLER_161_196 ();
 sg13g2_decap_8 FILLER_161_203 ();
 sg13g2_decap_8 FILLER_161_210 ();
 sg13g2_decap_8 FILLER_161_217 ();
 sg13g2_decap_8 FILLER_161_224 ();
 sg13g2_decap_8 FILLER_161_231 ();
 sg13g2_fill_2 FILLER_161_238 ();
 sg13g2_decap_8 FILLER_161_244 ();
 sg13g2_decap_8 FILLER_161_251 ();
 sg13g2_decap_4 FILLER_161_258 ();
 sg13g2_decap_8 FILLER_161_266 ();
 sg13g2_decap_8 FILLER_161_273 ();
 sg13g2_fill_2 FILLER_161_280 ();
 sg13g2_fill_1 FILLER_161_286 ();
 sg13g2_fill_1 FILLER_161_299 ();
 sg13g2_decap_4 FILLER_161_334 ();
 sg13g2_fill_2 FILLER_161_338 ();
 sg13g2_fill_2 FILLER_161_382 ();
 sg13g2_fill_2 FILLER_161_410 ();
 sg13g2_fill_1 FILLER_161_412 ();
 sg13g2_fill_1 FILLER_161_439 ();
 sg13g2_fill_2 FILLER_161_450 ();
 sg13g2_decap_8 FILLER_161_487 ();
 sg13g2_decap_4 FILLER_161_494 ();
 sg13g2_fill_1 FILLER_161_498 ();
 sg13g2_fill_2 FILLER_161_503 ();
 sg13g2_fill_1 FILLER_161_505 ();
 sg13g2_decap_4 FILLER_161_510 ();
 sg13g2_fill_2 FILLER_161_518 ();
 sg13g2_fill_1 FILLER_161_520 ();
 sg13g2_decap_8 FILLER_161_525 ();
 sg13g2_decap_8 FILLER_161_532 ();
 sg13g2_decap_4 FILLER_161_539 ();
 sg13g2_fill_2 FILLER_161_543 ();
 sg13g2_decap_4 FILLER_161_584 ();
 sg13g2_decap_8 FILLER_161_640 ();
 sg13g2_fill_2 FILLER_161_688 ();
 sg13g2_fill_2 FILLER_161_696 ();
 sg13g2_decap_4 FILLER_161_702 ();
 sg13g2_fill_1 FILLER_161_706 ();
 sg13g2_fill_1 FILLER_161_712 ();
 sg13g2_decap_8 FILLER_161_717 ();
 sg13g2_decap_8 FILLER_161_724 ();
 sg13g2_decap_8 FILLER_161_731 ();
 sg13g2_fill_2 FILLER_161_777 ();
 sg13g2_decap_8 FILLER_161_782 ();
 sg13g2_decap_8 FILLER_161_789 ();
 sg13g2_decap_8 FILLER_161_796 ();
 sg13g2_fill_2 FILLER_161_803 ();
 sg13g2_fill_2 FILLER_161_831 ();
 sg13g2_fill_2 FILLER_161_896 ();
 sg13g2_fill_1 FILLER_161_898 ();
 sg13g2_fill_1 FILLER_161_937 ();
 sg13g2_decap_4 FILLER_161_974 ();
 sg13g2_fill_2 FILLER_161_978 ();
 sg13g2_decap_8 FILLER_161_1061 ();
 sg13g2_fill_1 FILLER_161_1068 ();
 sg13g2_decap_8 FILLER_161_1073 ();
 sg13g2_decap_8 FILLER_161_1084 ();
 sg13g2_decap_8 FILLER_161_1091 ();
 sg13g2_decap_8 FILLER_161_1098 ();
 sg13g2_decap_8 FILLER_161_1133 ();
 sg13g2_decap_8 FILLER_161_1140 ();
 sg13g2_decap_4 FILLER_161_1147 ();
 sg13g2_fill_1 FILLER_161_1151 ();
 sg13g2_fill_2 FILLER_161_1157 ();
 sg13g2_fill_1 FILLER_161_1159 ();
 sg13g2_decap_8 FILLER_161_1164 ();
 sg13g2_decap_8 FILLER_161_1176 ();
 sg13g2_fill_1 FILLER_161_1183 ();
 sg13g2_decap_8 FILLER_161_1194 ();
 sg13g2_fill_2 FILLER_161_1201 ();
 sg13g2_fill_1 FILLER_161_1203 ();
 sg13g2_fill_2 FILLER_161_1219 ();
 sg13g2_decap_8 FILLER_161_1251 ();
 sg13g2_fill_2 FILLER_161_1258 ();
 sg13g2_decap_8 FILLER_161_1267 ();
 sg13g2_decap_8 FILLER_161_1274 ();
 sg13g2_decap_4 FILLER_161_1281 ();
 sg13g2_fill_2 FILLER_161_1285 ();
 sg13g2_fill_2 FILLER_161_1299 ();
 sg13g2_decap_8 FILLER_161_1327 ();
 sg13g2_decap_8 FILLER_161_1334 ();
 sg13g2_decap_8 FILLER_161_1341 ();
 sg13g2_decap_8 FILLER_161_1348 ();
 sg13g2_decap_8 FILLER_161_1355 ();
 sg13g2_decap_8 FILLER_161_1362 ();
 sg13g2_decap_8 FILLER_161_1369 ();
 sg13g2_decap_8 FILLER_161_1376 ();
 sg13g2_decap_8 FILLER_161_1383 ();
 sg13g2_decap_8 FILLER_161_1390 ();
 sg13g2_decap_8 FILLER_161_1397 ();
 sg13g2_decap_8 FILLER_161_1404 ();
 sg13g2_decap_8 FILLER_161_1411 ();
 sg13g2_decap_8 FILLER_161_1418 ();
 sg13g2_decap_8 FILLER_161_1425 ();
 sg13g2_decap_8 FILLER_161_1432 ();
 sg13g2_decap_8 FILLER_161_1439 ();
 sg13g2_decap_8 FILLER_161_1446 ();
 sg13g2_decap_8 FILLER_161_1453 ();
 sg13g2_decap_8 FILLER_161_1460 ();
 sg13g2_decap_8 FILLER_161_1467 ();
 sg13g2_decap_8 FILLER_161_1474 ();
 sg13g2_decap_8 FILLER_161_1481 ();
 sg13g2_decap_8 FILLER_161_1488 ();
 sg13g2_decap_8 FILLER_161_1495 ();
 sg13g2_decap_8 FILLER_161_1502 ();
 sg13g2_decap_8 FILLER_161_1509 ();
 sg13g2_decap_8 FILLER_161_1516 ();
 sg13g2_decap_8 FILLER_161_1523 ();
 sg13g2_decap_8 FILLER_161_1530 ();
 sg13g2_decap_8 FILLER_161_1537 ();
 sg13g2_decap_8 FILLER_161_1544 ();
 sg13g2_decap_8 FILLER_161_1551 ();
 sg13g2_decap_8 FILLER_161_1558 ();
 sg13g2_decap_8 FILLER_161_1565 ();
 sg13g2_decap_8 FILLER_161_1572 ();
 sg13g2_decap_8 FILLER_161_1579 ();
 sg13g2_decap_8 FILLER_161_1586 ();
 sg13g2_decap_8 FILLER_161_1593 ();
 sg13g2_decap_8 FILLER_161_1600 ();
 sg13g2_decap_8 FILLER_161_1607 ();
 sg13g2_decap_8 FILLER_161_1614 ();
 sg13g2_decap_4 FILLER_161_1621 ();
 sg13g2_decap_8 FILLER_162_0 ();
 sg13g2_decap_8 FILLER_162_7 ();
 sg13g2_decap_8 FILLER_162_14 ();
 sg13g2_fill_2 FILLER_162_21 ();
 sg13g2_decap_8 FILLER_162_27 ();
 sg13g2_decap_8 FILLER_162_34 ();
 sg13g2_decap_8 FILLER_162_41 ();
 sg13g2_fill_1 FILLER_162_48 ();
 sg13g2_decap_8 FILLER_162_75 ();
 sg13g2_decap_8 FILLER_162_82 ();
 sg13g2_decap_8 FILLER_162_89 ();
 sg13g2_decap_8 FILLER_162_96 ();
 sg13g2_decap_8 FILLER_162_103 ();
 sg13g2_decap_8 FILLER_162_110 ();
 sg13g2_decap_8 FILLER_162_117 ();
 sg13g2_decap_8 FILLER_162_124 ();
 sg13g2_decap_8 FILLER_162_131 ();
 sg13g2_decap_8 FILLER_162_138 ();
 sg13g2_decap_8 FILLER_162_145 ();
 sg13g2_decap_8 FILLER_162_152 ();
 sg13g2_decap_8 FILLER_162_159 ();
 sg13g2_decap_8 FILLER_162_166 ();
 sg13g2_decap_8 FILLER_162_173 ();
 sg13g2_decap_8 FILLER_162_180 ();
 sg13g2_decap_8 FILLER_162_187 ();
 sg13g2_decap_8 FILLER_162_194 ();
 sg13g2_decap_4 FILLER_162_201 ();
 sg13g2_decap_8 FILLER_162_209 ();
 sg13g2_decap_8 FILLER_162_216 ();
 sg13g2_decap_8 FILLER_162_223 ();
 sg13g2_fill_1 FILLER_162_230 ();
 sg13g2_fill_1 FILLER_162_286 ();
 sg13g2_decap_8 FILLER_162_310 ();
 sg13g2_decap_4 FILLER_162_317 ();
 sg13g2_fill_1 FILLER_162_336 ();
 sg13g2_fill_2 FILLER_162_363 ();
 sg13g2_fill_1 FILLER_162_365 ();
 sg13g2_decap_8 FILLER_162_370 ();
 sg13g2_fill_2 FILLER_162_377 ();
 sg13g2_decap_8 FILLER_162_383 ();
 sg13g2_fill_1 FILLER_162_390 ();
 sg13g2_fill_1 FILLER_162_425 ();
 sg13g2_decap_8 FILLER_162_459 ();
 sg13g2_decap_4 FILLER_162_466 ();
 sg13g2_fill_1 FILLER_162_470 ();
 sg13g2_fill_2 FILLER_162_500 ();
 sg13g2_fill_1 FILLER_162_502 ();
 sg13g2_fill_2 FILLER_162_513 ();
 sg13g2_decap_8 FILLER_162_519 ();
 sg13g2_decap_4 FILLER_162_526 ();
 sg13g2_fill_2 FILLER_162_530 ();
 sg13g2_decap_8 FILLER_162_568 ();
 sg13g2_decap_8 FILLER_162_575 ();
 sg13g2_decap_8 FILLER_162_582 ();
 sg13g2_decap_8 FILLER_162_589 ();
 sg13g2_decap_8 FILLER_162_596 ();
 sg13g2_decap_4 FILLER_162_603 ();
 sg13g2_fill_2 FILLER_162_607 ();
 sg13g2_fill_2 FILLER_162_638 ();
 sg13g2_decap_8 FILLER_162_693 ();
 sg13g2_fill_1 FILLER_162_700 ();
 sg13g2_fill_2 FILLER_162_727 ();
 sg13g2_fill_2 FILLER_162_755 ();
 sg13g2_fill_1 FILLER_162_757 ();
 sg13g2_decap_4 FILLER_162_813 ();
 sg13g2_fill_2 FILLER_162_817 ();
 sg13g2_decap_8 FILLER_162_849 ();
 sg13g2_decap_8 FILLER_162_856 ();
 sg13g2_decap_8 FILLER_162_863 ();
 sg13g2_fill_1 FILLER_162_870 ();
 sg13g2_decap_8 FILLER_162_875 ();
 sg13g2_decap_8 FILLER_162_882 ();
 sg13g2_decap_8 FILLER_162_889 ();
 sg13g2_decap_8 FILLER_162_896 ();
 sg13g2_decap_8 FILLER_162_903 ();
 sg13g2_fill_2 FILLER_162_952 ();
 sg13g2_fill_1 FILLER_162_954 ();
 sg13g2_fill_1 FILLER_162_995 ();
 sg13g2_decap_8 FILLER_162_1029 ();
 sg13g2_decap_8 FILLER_162_1036 ();
 sg13g2_decap_8 FILLER_162_1043 ();
 sg13g2_decap_8 FILLER_162_1050 ();
 sg13g2_fill_1 FILLER_162_1057 ();
 sg13g2_fill_1 FILLER_162_1063 ();
 sg13g2_fill_1 FILLER_162_1072 ();
 sg13g2_decap_8 FILLER_162_1104 ();
 sg13g2_decap_4 FILLER_162_1111 ();
 sg13g2_decap_4 FILLER_162_1141 ();
 sg13g2_fill_2 FILLER_162_1145 ();
 sg13g2_fill_1 FILLER_162_1179 ();
 sg13g2_decap_8 FILLER_162_1185 ();
 sg13g2_decap_4 FILLER_162_1192 ();
 sg13g2_fill_1 FILLER_162_1196 ();
 sg13g2_decap_8 FILLER_162_1211 ();
 sg13g2_decap_8 FILLER_162_1218 ();
 sg13g2_decap_8 FILLER_162_1225 ();
 sg13g2_fill_2 FILLER_162_1232 ();
 sg13g2_decap_8 FILLER_162_1238 ();
 sg13g2_decap_8 FILLER_162_1245 ();
 sg13g2_fill_2 FILLER_162_1252 ();
 sg13g2_fill_2 FILLER_162_1260 ();
 sg13g2_decap_4 FILLER_162_1270 ();
 sg13g2_fill_2 FILLER_162_1274 ();
 sg13g2_decap_8 FILLER_162_1280 ();
 sg13g2_decap_4 FILLER_162_1287 ();
 sg13g2_fill_1 FILLER_162_1291 ();
 sg13g2_fill_2 FILLER_162_1300 ();
 sg13g2_decap_8 FILLER_162_1331 ();
 sg13g2_decap_8 FILLER_162_1338 ();
 sg13g2_decap_8 FILLER_162_1345 ();
 sg13g2_decap_8 FILLER_162_1352 ();
 sg13g2_decap_8 FILLER_162_1359 ();
 sg13g2_decap_8 FILLER_162_1366 ();
 sg13g2_decap_8 FILLER_162_1373 ();
 sg13g2_decap_8 FILLER_162_1380 ();
 sg13g2_decap_8 FILLER_162_1387 ();
 sg13g2_decap_8 FILLER_162_1394 ();
 sg13g2_decap_8 FILLER_162_1401 ();
 sg13g2_decap_8 FILLER_162_1408 ();
 sg13g2_decap_8 FILLER_162_1415 ();
 sg13g2_decap_8 FILLER_162_1422 ();
 sg13g2_decap_8 FILLER_162_1429 ();
 sg13g2_decap_8 FILLER_162_1436 ();
 sg13g2_decap_8 FILLER_162_1443 ();
 sg13g2_decap_8 FILLER_162_1450 ();
 sg13g2_decap_8 FILLER_162_1457 ();
 sg13g2_decap_8 FILLER_162_1464 ();
 sg13g2_decap_8 FILLER_162_1471 ();
 sg13g2_decap_8 FILLER_162_1478 ();
 sg13g2_decap_8 FILLER_162_1485 ();
 sg13g2_decap_8 FILLER_162_1492 ();
 sg13g2_decap_8 FILLER_162_1499 ();
 sg13g2_decap_8 FILLER_162_1506 ();
 sg13g2_decap_8 FILLER_162_1513 ();
 sg13g2_decap_8 FILLER_162_1520 ();
 sg13g2_decap_8 FILLER_162_1527 ();
 sg13g2_decap_8 FILLER_162_1534 ();
 sg13g2_decap_8 FILLER_162_1541 ();
 sg13g2_decap_8 FILLER_162_1548 ();
 sg13g2_decap_8 FILLER_162_1555 ();
 sg13g2_decap_8 FILLER_162_1562 ();
 sg13g2_decap_8 FILLER_162_1569 ();
 sg13g2_decap_8 FILLER_162_1576 ();
 sg13g2_decap_8 FILLER_162_1583 ();
 sg13g2_decap_8 FILLER_162_1590 ();
 sg13g2_decap_8 FILLER_162_1597 ();
 sg13g2_decap_8 FILLER_162_1604 ();
 sg13g2_decap_8 FILLER_162_1611 ();
 sg13g2_decap_8 FILLER_162_1618 ();
 sg13g2_decap_8 FILLER_163_0 ();
 sg13g2_decap_8 FILLER_163_7 ();
 sg13g2_decap_8 FILLER_163_14 ();
 sg13g2_decap_8 FILLER_163_21 ();
 sg13g2_decap_8 FILLER_163_28 ();
 sg13g2_decap_8 FILLER_163_35 ();
 sg13g2_decap_8 FILLER_163_42 ();
 sg13g2_decap_8 FILLER_163_49 ();
 sg13g2_decap_8 FILLER_163_56 ();
 sg13g2_decap_8 FILLER_163_63 ();
 sg13g2_decap_8 FILLER_163_70 ();
 sg13g2_decap_8 FILLER_163_77 ();
 sg13g2_decap_8 FILLER_163_84 ();
 sg13g2_decap_8 FILLER_163_91 ();
 sg13g2_decap_8 FILLER_163_98 ();
 sg13g2_decap_8 FILLER_163_105 ();
 sg13g2_decap_8 FILLER_163_112 ();
 sg13g2_decap_8 FILLER_163_119 ();
 sg13g2_decap_8 FILLER_163_126 ();
 sg13g2_decap_8 FILLER_163_133 ();
 sg13g2_decap_8 FILLER_163_140 ();
 sg13g2_decap_8 FILLER_163_147 ();
 sg13g2_decap_8 FILLER_163_154 ();
 sg13g2_decap_8 FILLER_163_161 ();
 sg13g2_decap_8 FILLER_163_168 ();
 sg13g2_decap_8 FILLER_163_175 ();
 sg13g2_decap_8 FILLER_163_182 ();
 sg13g2_decap_4 FILLER_163_189 ();
 sg13g2_fill_2 FILLER_163_193 ();
 sg13g2_fill_2 FILLER_163_225 ();
 sg13g2_fill_1 FILLER_163_231 ();
 sg13g2_fill_2 FILLER_163_268 ();
 sg13g2_fill_1 FILLER_163_279 ();
 sg13g2_fill_1 FILLER_163_314 ();
 sg13g2_fill_2 FILLER_163_319 ();
 sg13g2_decap_8 FILLER_163_346 ();
 sg13g2_decap_4 FILLER_163_353 ();
 sg13g2_decap_4 FILLER_163_371 ();
 sg13g2_fill_1 FILLER_163_375 ();
 sg13g2_fill_2 FILLER_163_381 ();
 sg13g2_fill_2 FILLER_163_412 ();
 sg13g2_fill_1 FILLER_163_414 ();
 sg13g2_fill_1 FILLER_163_435 ();
 sg13g2_decap_4 FILLER_163_441 ();
 sg13g2_fill_2 FILLER_163_454 ();
 sg13g2_fill_1 FILLER_163_456 ();
 sg13g2_decap_4 FILLER_163_463 ();
 sg13g2_fill_1 FILLER_163_471 ();
 sg13g2_decap_8 FILLER_163_534 ();
 sg13g2_decap_8 FILLER_163_541 ();
 sg13g2_fill_2 FILLER_163_548 ();
 sg13g2_fill_1 FILLER_163_550 ();
 sg13g2_fill_2 FILLER_163_561 ();
 sg13g2_fill_1 FILLER_163_563 ();
 sg13g2_decap_8 FILLER_163_574 ();
 sg13g2_fill_2 FILLER_163_581 ();
 sg13g2_decap_4 FILLER_163_615 ();
 sg13g2_fill_1 FILLER_163_619 ();
 sg13g2_decap_8 FILLER_163_649 ();
 sg13g2_decap_8 FILLER_163_656 ();
 sg13g2_decap_8 FILLER_163_663 ();
 sg13g2_decap_8 FILLER_163_670 ();
 sg13g2_decap_8 FILLER_163_677 ();
 sg13g2_decap_8 FILLER_163_684 ();
 sg13g2_decap_8 FILLER_163_691 ();
 sg13g2_fill_2 FILLER_163_698 ();
 sg13g2_fill_1 FILLER_163_700 ();
 sg13g2_decap_8 FILLER_163_706 ();
 sg13g2_decap_8 FILLER_163_713 ();
 sg13g2_decap_8 FILLER_163_720 ();
 sg13g2_decap_8 FILLER_163_727 ();
 sg13g2_fill_2 FILLER_163_734 ();
 sg13g2_fill_1 FILLER_163_736 ();
 sg13g2_decap_8 FILLER_163_741 ();
 sg13g2_fill_2 FILLER_163_748 ();
 sg13g2_fill_2 FILLER_163_760 ();
 sg13g2_fill_1 FILLER_163_767 ();
 sg13g2_decap_8 FILLER_163_777 ();
 sg13g2_fill_2 FILLER_163_784 ();
 sg13g2_decap_8 FILLER_163_790 ();
 sg13g2_decap_4 FILLER_163_797 ();
 sg13g2_decap_8 FILLER_163_831 ();
 sg13g2_decap_8 FILLER_163_838 ();
 sg13g2_fill_2 FILLER_163_845 ();
 sg13g2_fill_1 FILLER_163_847 ();
 sg13g2_decap_8 FILLER_163_898 ();
 sg13g2_fill_2 FILLER_163_905 ();
 sg13g2_decap_4 FILLER_163_941 ();
 sg13g2_fill_1 FILLER_163_945 ();
 sg13g2_fill_2 FILLER_163_976 ();
 sg13g2_fill_2 FILLER_163_986 ();
 sg13g2_fill_1 FILLER_163_988 ();
 sg13g2_fill_2 FILLER_163_1023 ();
 sg13g2_fill_1 FILLER_163_1025 ();
 sg13g2_fill_1 FILLER_163_1072 ();
 sg13g2_decap_8 FILLER_163_1098 ();
 sg13g2_fill_2 FILLER_163_1105 ();
 sg13g2_fill_2 FILLER_163_1128 ();
 sg13g2_decap_8 FILLER_163_1147 ();
 sg13g2_fill_1 FILLER_163_1180 ();
 sg13g2_fill_1 FILLER_163_1185 ();
 sg13g2_fill_1 FILLER_163_1191 ();
 sg13g2_decap_8 FILLER_163_1195 ();
 sg13g2_decap_4 FILLER_163_1202 ();
 sg13g2_decap_8 FILLER_163_1217 ();
 sg13g2_decap_4 FILLER_163_1224 ();
 sg13g2_fill_2 FILLER_163_1228 ();
 sg13g2_decap_8 FILLER_163_1234 ();
 sg13g2_decap_8 FILLER_163_1241 ();
 sg13g2_fill_2 FILLER_163_1248 ();
 sg13g2_fill_1 FILLER_163_1250 ();
 sg13g2_fill_2 FILLER_163_1266 ();
 sg13g2_fill_2 FILLER_163_1299 ();
 sg13g2_decap_8 FILLER_163_1327 ();
 sg13g2_decap_8 FILLER_163_1334 ();
 sg13g2_decap_8 FILLER_163_1341 ();
 sg13g2_decap_8 FILLER_163_1348 ();
 sg13g2_decap_8 FILLER_163_1355 ();
 sg13g2_decap_8 FILLER_163_1362 ();
 sg13g2_decap_8 FILLER_163_1369 ();
 sg13g2_decap_8 FILLER_163_1376 ();
 sg13g2_decap_8 FILLER_163_1383 ();
 sg13g2_decap_8 FILLER_163_1390 ();
 sg13g2_decap_8 FILLER_163_1397 ();
 sg13g2_decap_8 FILLER_163_1404 ();
 sg13g2_decap_8 FILLER_163_1411 ();
 sg13g2_decap_8 FILLER_163_1418 ();
 sg13g2_decap_8 FILLER_163_1425 ();
 sg13g2_decap_8 FILLER_163_1432 ();
 sg13g2_decap_8 FILLER_163_1439 ();
 sg13g2_decap_8 FILLER_163_1446 ();
 sg13g2_decap_8 FILLER_163_1453 ();
 sg13g2_decap_8 FILLER_163_1460 ();
 sg13g2_decap_8 FILLER_163_1467 ();
 sg13g2_decap_8 FILLER_163_1474 ();
 sg13g2_decap_8 FILLER_163_1481 ();
 sg13g2_decap_8 FILLER_163_1488 ();
 sg13g2_decap_8 FILLER_163_1495 ();
 sg13g2_decap_8 FILLER_163_1502 ();
 sg13g2_decap_8 FILLER_163_1509 ();
 sg13g2_decap_8 FILLER_163_1516 ();
 sg13g2_decap_8 FILLER_163_1523 ();
 sg13g2_decap_8 FILLER_163_1530 ();
 sg13g2_decap_8 FILLER_163_1537 ();
 sg13g2_decap_8 FILLER_163_1544 ();
 sg13g2_decap_8 FILLER_163_1551 ();
 sg13g2_decap_8 FILLER_163_1558 ();
 sg13g2_decap_8 FILLER_163_1565 ();
 sg13g2_decap_8 FILLER_163_1572 ();
 sg13g2_decap_8 FILLER_163_1579 ();
 sg13g2_decap_8 FILLER_163_1586 ();
 sg13g2_decap_8 FILLER_163_1593 ();
 sg13g2_decap_8 FILLER_163_1600 ();
 sg13g2_decap_8 FILLER_163_1607 ();
 sg13g2_decap_8 FILLER_163_1614 ();
 sg13g2_decap_4 FILLER_163_1621 ();
 sg13g2_decap_8 FILLER_164_0 ();
 sg13g2_decap_8 FILLER_164_7 ();
 sg13g2_decap_8 FILLER_164_14 ();
 sg13g2_decap_8 FILLER_164_21 ();
 sg13g2_decap_8 FILLER_164_28 ();
 sg13g2_decap_8 FILLER_164_35 ();
 sg13g2_decap_8 FILLER_164_42 ();
 sg13g2_decap_8 FILLER_164_49 ();
 sg13g2_decap_8 FILLER_164_56 ();
 sg13g2_decap_8 FILLER_164_63 ();
 sg13g2_decap_8 FILLER_164_70 ();
 sg13g2_decap_8 FILLER_164_77 ();
 sg13g2_decap_8 FILLER_164_84 ();
 sg13g2_decap_8 FILLER_164_91 ();
 sg13g2_decap_8 FILLER_164_98 ();
 sg13g2_decap_8 FILLER_164_105 ();
 sg13g2_decap_8 FILLER_164_112 ();
 sg13g2_decap_8 FILLER_164_119 ();
 sg13g2_decap_8 FILLER_164_126 ();
 sg13g2_decap_8 FILLER_164_133 ();
 sg13g2_decap_8 FILLER_164_140 ();
 sg13g2_decap_8 FILLER_164_147 ();
 sg13g2_decap_8 FILLER_164_154 ();
 sg13g2_decap_8 FILLER_164_161 ();
 sg13g2_decap_8 FILLER_164_168 ();
 sg13g2_decap_8 FILLER_164_175 ();
 sg13g2_decap_8 FILLER_164_182 ();
 sg13g2_decap_4 FILLER_164_189 ();
 sg13g2_decap_8 FILLER_164_201 ();
 sg13g2_fill_2 FILLER_164_208 ();
 sg13g2_decap_4 FILLER_164_221 ();
 sg13g2_decap_4 FILLER_164_237 ();
 sg13g2_fill_2 FILLER_164_241 ();
 sg13g2_fill_1 FILLER_164_275 ();
 sg13g2_fill_1 FILLER_164_282 ();
 sg13g2_decap_8 FILLER_164_340 ();
 sg13g2_fill_2 FILLER_164_347 ();
 sg13g2_decap_8 FILLER_164_353 ();
 sg13g2_decap_8 FILLER_164_365 ();
 sg13g2_decap_4 FILLER_164_372 ();
 sg13g2_fill_1 FILLER_164_376 ();
 sg13g2_fill_2 FILLER_164_438 ();
 sg13g2_fill_1 FILLER_164_440 ();
 sg13g2_decap_4 FILLER_164_445 ();
 sg13g2_fill_2 FILLER_164_449 ();
 sg13g2_decap_8 FILLER_164_490 ();
 sg13g2_decap_8 FILLER_164_497 ();
 sg13g2_decap_8 FILLER_164_504 ();
 sg13g2_decap_8 FILLER_164_511 ();
 sg13g2_decap_8 FILLER_164_518 ();
 sg13g2_decap_8 FILLER_164_525 ();
 sg13g2_decap_8 FILLER_164_536 ();
 sg13g2_decap_4 FILLER_164_543 ();
 sg13g2_fill_2 FILLER_164_547 ();
 sg13g2_fill_1 FILLER_164_600 ();
 sg13g2_fill_2 FILLER_164_627 ();
 sg13g2_fill_1 FILLER_164_629 ();
 sg13g2_fill_2 FILLER_164_661 ();
 sg13g2_fill_1 FILLER_164_663 ();
 sg13g2_decap_8 FILLER_164_668 ();
 sg13g2_decap_8 FILLER_164_685 ();
 sg13g2_fill_1 FILLER_164_692 ();
 sg13g2_decap_8 FILLER_164_697 ();
 sg13g2_decap_4 FILLER_164_704 ();
 sg13g2_decap_4 FILLER_164_716 ();
 sg13g2_fill_1 FILLER_164_720 ();
 sg13g2_decap_4 FILLER_164_734 ();
 sg13g2_decap_8 FILLER_164_741 ();
 sg13g2_decap_8 FILLER_164_748 ();
 sg13g2_decap_8 FILLER_164_755 ();
 sg13g2_decap_4 FILLER_164_762 ();
 sg13g2_decap_8 FILLER_164_807 ();
 sg13g2_decap_8 FILLER_164_814 ();
 sg13g2_decap_8 FILLER_164_821 ();
 sg13g2_decap_8 FILLER_164_828 ();
 sg13g2_decap_8 FILLER_164_835 ();
 sg13g2_decap_8 FILLER_164_842 ();
 sg13g2_decap_8 FILLER_164_849 ();
 sg13g2_decap_8 FILLER_164_860 ();
 sg13g2_decap_4 FILLER_164_867 ();
 sg13g2_fill_2 FILLER_164_901 ();
 sg13g2_fill_1 FILLER_164_911 ();
 sg13g2_decap_8 FILLER_164_1007 ();
 sg13g2_decap_4 FILLER_164_1014 ();
 sg13g2_fill_1 FILLER_164_1018 ();
 sg13g2_fill_2 FILLER_164_1058 ();
 sg13g2_decap_4 FILLER_164_1115 ();
 sg13g2_decap_8 FILLER_164_1123 ();
 sg13g2_fill_2 FILLER_164_1130 ();
 sg13g2_decap_8 FILLER_164_1136 ();
 sg13g2_fill_1 FILLER_164_1143 ();
 sg13g2_fill_2 FILLER_164_1148 ();
 sg13g2_decap_8 FILLER_164_1154 ();
 sg13g2_decap_8 FILLER_164_1161 ();
 sg13g2_fill_2 FILLER_164_1168 ();
 sg13g2_fill_1 FILLER_164_1175 ();
 sg13g2_fill_1 FILLER_164_1198 ();
 sg13g2_decap_8 FILLER_164_1204 ();
 sg13g2_decap_8 FILLER_164_1211 ();
 sg13g2_decap_8 FILLER_164_1249 ();
 sg13g2_decap_8 FILLER_164_1256 ();
 sg13g2_fill_2 FILLER_164_1263 ();
 sg13g2_decap_8 FILLER_164_1273 ();
 sg13g2_decap_8 FILLER_164_1280 ();
 sg13g2_decap_8 FILLER_164_1287 ();
 sg13g2_decap_4 FILLER_164_1294 ();
 sg13g2_decap_4 FILLER_164_1309 ();
 sg13g2_fill_2 FILLER_164_1313 ();
 sg13g2_decap_8 FILLER_164_1341 ();
 sg13g2_decap_8 FILLER_164_1348 ();
 sg13g2_decap_8 FILLER_164_1355 ();
 sg13g2_decap_8 FILLER_164_1362 ();
 sg13g2_decap_8 FILLER_164_1369 ();
 sg13g2_decap_8 FILLER_164_1376 ();
 sg13g2_decap_8 FILLER_164_1383 ();
 sg13g2_decap_8 FILLER_164_1390 ();
 sg13g2_decap_8 FILLER_164_1397 ();
 sg13g2_decap_8 FILLER_164_1404 ();
 sg13g2_decap_8 FILLER_164_1411 ();
 sg13g2_decap_8 FILLER_164_1418 ();
 sg13g2_decap_8 FILLER_164_1425 ();
 sg13g2_decap_8 FILLER_164_1432 ();
 sg13g2_decap_8 FILLER_164_1439 ();
 sg13g2_decap_8 FILLER_164_1446 ();
 sg13g2_decap_8 FILLER_164_1453 ();
 sg13g2_decap_8 FILLER_164_1460 ();
 sg13g2_decap_8 FILLER_164_1467 ();
 sg13g2_decap_8 FILLER_164_1474 ();
 sg13g2_decap_8 FILLER_164_1481 ();
 sg13g2_decap_8 FILLER_164_1488 ();
 sg13g2_decap_8 FILLER_164_1495 ();
 sg13g2_decap_8 FILLER_164_1502 ();
 sg13g2_decap_8 FILLER_164_1509 ();
 sg13g2_decap_8 FILLER_164_1516 ();
 sg13g2_decap_8 FILLER_164_1523 ();
 sg13g2_decap_8 FILLER_164_1530 ();
 sg13g2_decap_8 FILLER_164_1537 ();
 sg13g2_decap_8 FILLER_164_1544 ();
 sg13g2_decap_8 FILLER_164_1551 ();
 sg13g2_decap_8 FILLER_164_1558 ();
 sg13g2_decap_8 FILLER_164_1565 ();
 sg13g2_decap_8 FILLER_164_1572 ();
 sg13g2_decap_8 FILLER_164_1579 ();
 sg13g2_decap_8 FILLER_164_1586 ();
 sg13g2_decap_8 FILLER_164_1593 ();
 sg13g2_decap_8 FILLER_164_1600 ();
 sg13g2_decap_8 FILLER_164_1607 ();
 sg13g2_decap_8 FILLER_164_1614 ();
 sg13g2_decap_4 FILLER_164_1621 ();
 sg13g2_decap_8 FILLER_165_0 ();
 sg13g2_decap_8 FILLER_165_7 ();
 sg13g2_decap_8 FILLER_165_14 ();
 sg13g2_decap_8 FILLER_165_21 ();
 sg13g2_decap_8 FILLER_165_28 ();
 sg13g2_decap_8 FILLER_165_35 ();
 sg13g2_decap_8 FILLER_165_42 ();
 sg13g2_decap_8 FILLER_165_49 ();
 sg13g2_decap_8 FILLER_165_56 ();
 sg13g2_decap_8 FILLER_165_63 ();
 sg13g2_decap_8 FILLER_165_70 ();
 sg13g2_decap_8 FILLER_165_77 ();
 sg13g2_decap_8 FILLER_165_84 ();
 sg13g2_decap_8 FILLER_165_91 ();
 sg13g2_decap_8 FILLER_165_98 ();
 sg13g2_decap_8 FILLER_165_105 ();
 sg13g2_decap_8 FILLER_165_112 ();
 sg13g2_decap_8 FILLER_165_119 ();
 sg13g2_decap_8 FILLER_165_126 ();
 sg13g2_decap_8 FILLER_165_133 ();
 sg13g2_decap_8 FILLER_165_140 ();
 sg13g2_decap_8 FILLER_165_147 ();
 sg13g2_decap_8 FILLER_165_154 ();
 sg13g2_decap_8 FILLER_165_161 ();
 sg13g2_fill_2 FILLER_165_168 ();
 sg13g2_decap_8 FILLER_165_174 ();
 sg13g2_decap_8 FILLER_165_181 ();
 sg13g2_decap_4 FILLER_165_218 ();
 sg13g2_decap_8 FILLER_165_227 ();
 sg13g2_decap_4 FILLER_165_234 ();
 sg13g2_fill_1 FILLER_165_238 ();
 sg13g2_decap_4 FILLER_165_255 ();
 sg13g2_fill_1 FILLER_165_259 ();
 sg13g2_decap_4 FILLER_165_265 ();
 sg13g2_fill_1 FILLER_165_269 ();
 sg13g2_fill_2 FILLER_165_280 ();
 sg13g2_fill_1 FILLER_165_282 ();
 sg13g2_fill_2 FILLER_165_287 ();
 sg13g2_fill_1 FILLER_165_289 ();
 sg13g2_decap_8 FILLER_165_313 ();
 sg13g2_decap_8 FILLER_165_320 ();
 sg13g2_fill_2 FILLER_165_327 ();
 sg13g2_fill_2 FILLER_165_368 ();
 sg13g2_fill_1 FILLER_165_370 ();
 sg13g2_fill_2 FILLER_165_375 ();
 sg13g2_decap_4 FILLER_165_382 ();
 sg13g2_fill_1 FILLER_165_386 ();
 sg13g2_decap_8 FILLER_165_391 ();
 sg13g2_decap_8 FILLER_165_398 ();
 sg13g2_decap_4 FILLER_165_405 ();
 sg13g2_fill_2 FILLER_165_409 ();
 sg13g2_decap_8 FILLER_165_415 ();
 sg13g2_fill_2 FILLER_165_422 ();
 sg13g2_decap_8 FILLER_165_460 ();
 sg13g2_decap_8 FILLER_165_467 ();
 sg13g2_fill_2 FILLER_165_479 ();
 sg13g2_decap_4 FILLER_165_493 ();
 sg13g2_fill_2 FILLER_165_497 ();
 sg13g2_fill_2 FILLER_165_505 ();
 sg13g2_decap_4 FILLER_165_549 ();
 sg13g2_fill_1 FILLER_165_553 ();
 sg13g2_fill_1 FILLER_165_580 ();
 sg13g2_decap_8 FILLER_165_585 ();
 sg13g2_decap_8 FILLER_165_592 ();
 sg13g2_decap_8 FILLER_165_599 ();
 sg13g2_decap_8 FILLER_165_606 ();
 sg13g2_decap_8 FILLER_165_613 ();
 sg13g2_decap_8 FILLER_165_620 ();
 sg13g2_decap_8 FILLER_165_627 ();
 sg13g2_fill_2 FILLER_165_634 ();
 sg13g2_fill_1 FILLER_165_636 ();
 sg13g2_decap_4 FILLER_165_642 ();
 sg13g2_fill_1 FILLER_165_646 ();
 sg13g2_fill_2 FILLER_165_683 ();
 sg13g2_fill_1 FILLER_165_711 ();
 sg13g2_fill_2 FILLER_165_717 ();
 sg13g2_fill_1 FILLER_165_719 ();
 sg13g2_decap_4 FILLER_165_728 ();
 sg13g2_fill_2 FILLER_165_732 ();
 sg13g2_decap_4 FILLER_165_750 ();
 sg13g2_decap_8 FILLER_165_759 ();
 sg13g2_decap_8 FILLER_165_766 ();
 sg13g2_decap_8 FILLER_165_773 ();
 sg13g2_decap_8 FILLER_165_780 ();
 sg13g2_decap_8 FILLER_165_787 ();
 sg13g2_decap_4 FILLER_165_794 ();
 sg13g2_fill_1 FILLER_165_798 ();
 sg13g2_fill_1 FILLER_165_805 ();
 sg13g2_decap_8 FILLER_165_810 ();
 sg13g2_decap_8 FILLER_165_817 ();
 sg13g2_decap_8 FILLER_165_824 ();
 sg13g2_fill_1 FILLER_165_831 ();
 sg13g2_fill_1 FILLER_165_836 ();
 sg13g2_decap_8 FILLER_165_842 ();
 sg13g2_decap_8 FILLER_165_875 ();
 sg13g2_decap_8 FILLER_165_882 ();
 sg13g2_decap_8 FILLER_165_925 ();
 sg13g2_decap_8 FILLER_165_932 ();
 sg13g2_fill_1 FILLER_165_939 ();
 sg13g2_decap_8 FILLER_165_970 ();
 sg13g2_fill_2 FILLER_165_977 ();
 sg13g2_decap_4 FILLER_165_984 ();
 sg13g2_fill_1 FILLER_165_988 ();
 sg13g2_decap_8 FILLER_165_997 ();
 sg13g2_fill_2 FILLER_165_1004 ();
 sg13g2_fill_1 FILLER_165_1006 ();
 sg13g2_decap_8 FILLER_165_1011 ();
 sg13g2_decap_8 FILLER_165_1018 ();
 sg13g2_decap_8 FILLER_165_1025 ();
 sg13g2_decap_8 FILLER_165_1032 ();
 sg13g2_decap_8 FILLER_165_1039 ();
 sg13g2_decap_8 FILLER_165_1046 ();
 sg13g2_decap_8 FILLER_165_1053 ();
 sg13g2_decap_8 FILLER_165_1060 ();
 sg13g2_decap_8 FILLER_165_1067 ();
 sg13g2_fill_1 FILLER_165_1078 ();
 sg13g2_fill_2 FILLER_165_1083 ();
 sg13g2_decap_8 FILLER_165_1102 ();
 sg13g2_decap_4 FILLER_165_1109 ();
 sg13g2_fill_1 FILLER_165_1113 ();
 sg13g2_decap_8 FILLER_165_1126 ();
 sg13g2_decap_8 FILLER_165_1133 ();
 sg13g2_decap_8 FILLER_165_1140 ();
 sg13g2_fill_2 FILLER_165_1185 ();
 sg13g2_fill_2 FILLER_165_1205 ();
 sg13g2_fill_2 FILLER_165_1211 ();
 sg13g2_decap_4 FILLER_165_1242 ();
 sg13g2_fill_1 FILLER_165_1246 ();
 sg13g2_fill_2 FILLER_165_1259 ();
 sg13g2_fill_1 FILLER_165_1261 ();
 sg13g2_fill_2 FILLER_165_1268 ();
 sg13g2_fill_1 FILLER_165_1270 ();
 sg13g2_decap_4 FILLER_165_1277 ();
 sg13g2_fill_2 FILLER_165_1281 ();
 sg13g2_fill_2 FILLER_165_1290 ();
 sg13g2_fill_1 FILLER_165_1292 ();
 sg13g2_fill_1 FILLER_165_1306 ();
 sg13g2_decap_8 FILLER_165_1343 ();
 sg13g2_decap_8 FILLER_165_1350 ();
 sg13g2_decap_8 FILLER_165_1357 ();
 sg13g2_decap_8 FILLER_165_1364 ();
 sg13g2_decap_8 FILLER_165_1371 ();
 sg13g2_decap_8 FILLER_165_1378 ();
 sg13g2_decap_8 FILLER_165_1385 ();
 sg13g2_decap_8 FILLER_165_1392 ();
 sg13g2_decap_8 FILLER_165_1399 ();
 sg13g2_decap_8 FILLER_165_1406 ();
 sg13g2_decap_8 FILLER_165_1413 ();
 sg13g2_decap_8 FILLER_165_1420 ();
 sg13g2_decap_8 FILLER_165_1427 ();
 sg13g2_decap_8 FILLER_165_1434 ();
 sg13g2_decap_8 FILLER_165_1441 ();
 sg13g2_decap_8 FILLER_165_1448 ();
 sg13g2_decap_8 FILLER_165_1455 ();
 sg13g2_decap_8 FILLER_165_1462 ();
 sg13g2_decap_8 FILLER_165_1469 ();
 sg13g2_decap_8 FILLER_165_1476 ();
 sg13g2_decap_8 FILLER_165_1483 ();
 sg13g2_decap_8 FILLER_165_1490 ();
 sg13g2_decap_8 FILLER_165_1497 ();
 sg13g2_decap_8 FILLER_165_1504 ();
 sg13g2_decap_8 FILLER_165_1511 ();
 sg13g2_decap_8 FILLER_165_1518 ();
 sg13g2_decap_8 FILLER_165_1525 ();
 sg13g2_decap_8 FILLER_165_1532 ();
 sg13g2_decap_8 FILLER_165_1539 ();
 sg13g2_decap_8 FILLER_165_1546 ();
 sg13g2_decap_8 FILLER_165_1553 ();
 sg13g2_decap_8 FILLER_165_1560 ();
 sg13g2_decap_8 FILLER_165_1567 ();
 sg13g2_decap_8 FILLER_165_1574 ();
 sg13g2_decap_8 FILLER_165_1581 ();
 sg13g2_decap_8 FILLER_165_1588 ();
 sg13g2_decap_8 FILLER_165_1595 ();
 sg13g2_decap_8 FILLER_165_1602 ();
 sg13g2_decap_8 FILLER_165_1609 ();
 sg13g2_decap_8 FILLER_165_1616 ();
 sg13g2_fill_2 FILLER_165_1623 ();
 sg13g2_decap_8 FILLER_166_0 ();
 sg13g2_decap_8 FILLER_166_7 ();
 sg13g2_decap_8 FILLER_166_14 ();
 sg13g2_decap_8 FILLER_166_21 ();
 sg13g2_decap_8 FILLER_166_28 ();
 sg13g2_decap_8 FILLER_166_35 ();
 sg13g2_decap_8 FILLER_166_42 ();
 sg13g2_decap_8 FILLER_166_49 ();
 sg13g2_decap_8 FILLER_166_56 ();
 sg13g2_decap_8 FILLER_166_63 ();
 sg13g2_decap_8 FILLER_166_70 ();
 sg13g2_decap_8 FILLER_166_77 ();
 sg13g2_decap_8 FILLER_166_84 ();
 sg13g2_decap_8 FILLER_166_91 ();
 sg13g2_decap_8 FILLER_166_98 ();
 sg13g2_decap_8 FILLER_166_105 ();
 sg13g2_decap_8 FILLER_166_112 ();
 sg13g2_decap_8 FILLER_166_119 ();
 sg13g2_decap_8 FILLER_166_126 ();
 sg13g2_decap_8 FILLER_166_133 ();
 sg13g2_decap_8 FILLER_166_140 ();
 sg13g2_decap_8 FILLER_166_147 ();
 sg13g2_decap_8 FILLER_166_154 ();
 sg13g2_fill_2 FILLER_166_161 ();
 sg13g2_fill_1 FILLER_166_163 ();
 sg13g2_decap_4 FILLER_166_215 ();
 sg13g2_fill_2 FILLER_166_219 ();
 sg13g2_fill_2 FILLER_166_229 ();
 sg13g2_fill_2 FILLER_166_244 ();
 sg13g2_decap_8 FILLER_166_262 ();
 sg13g2_decap_8 FILLER_166_269 ();
 sg13g2_fill_2 FILLER_166_276 ();
 sg13g2_decap_8 FILLER_166_329 ();
 sg13g2_fill_2 FILLER_166_336 ();
 sg13g2_decap_8 FILLER_166_343 ();
 sg13g2_fill_2 FILLER_166_350 ();
 sg13g2_fill_1 FILLER_166_374 ();
 sg13g2_decap_8 FILLER_166_406 ();
 sg13g2_decap_8 FILLER_166_413 ();
 sg13g2_decap_4 FILLER_166_420 ();
 sg13g2_fill_1 FILLER_166_424 ();
 sg13g2_decap_8 FILLER_166_450 ();
 sg13g2_decap_4 FILLER_166_457 ();
 sg13g2_fill_2 FILLER_166_461 ();
 sg13g2_decap_8 FILLER_166_467 ();
 sg13g2_decap_8 FILLER_166_474 ();
 sg13g2_fill_2 FILLER_166_491 ();
 sg13g2_fill_2 FILLER_166_497 ();
 sg13g2_decap_4 FILLER_166_505 ();
 sg13g2_fill_1 FILLER_166_509 ();
 sg13g2_decap_8 FILLER_166_553 ();
 sg13g2_decap_8 FILLER_166_564 ();
 sg13g2_decap_4 FILLER_166_571 ();
 sg13g2_fill_1 FILLER_166_575 ();
 sg13g2_decap_8 FILLER_166_580 ();
 sg13g2_decap_4 FILLER_166_587 ();
 sg13g2_fill_1 FILLER_166_591 ();
 sg13g2_decap_4 FILLER_166_606 ();
 sg13g2_fill_1 FILLER_166_610 ();
 sg13g2_fill_2 FILLER_166_626 ();
 sg13g2_decap_4 FILLER_166_632 ();
 sg13g2_fill_2 FILLER_166_636 ();
 sg13g2_decap_8 FILLER_166_668 ();
 sg13g2_decap_8 FILLER_166_675 ();
 sg13g2_decap_4 FILLER_166_682 ();
 sg13g2_fill_1 FILLER_166_686 ();
 sg13g2_fill_2 FILLER_166_697 ();
 sg13g2_decap_8 FILLER_166_708 ();
 sg13g2_decap_8 FILLER_166_715 ();
 sg13g2_decap_8 FILLER_166_722 ();
 sg13g2_decap_4 FILLER_166_729 ();
 sg13g2_fill_2 FILLER_166_733 ();
 sg13g2_fill_1 FILLER_166_746 ();
 sg13g2_fill_2 FILLER_166_755 ();
 sg13g2_decap_4 FILLER_166_762 ();
 sg13g2_decap_4 FILLER_166_772 ();
 sg13g2_fill_1 FILLER_166_776 ();
 sg13g2_decap_8 FILLER_166_781 ();
 sg13g2_decap_4 FILLER_166_850 ();
 sg13g2_fill_2 FILLER_166_858 ();
 sg13g2_decap_4 FILLER_166_868 ();
 sg13g2_fill_1 FILLER_166_872 ();
 sg13g2_fill_2 FILLER_166_885 ();
 sg13g2_fill_1 FILLER_166_887 ();
 sg13g2_decap_4 FILLER_166_904 ();
 sg13g2_fill_1 FILLER_166_908 ();
 sg13g2_decap_8 FILLER_166_916 ();
 sg13g2_decap_8 FILLER_166_923 ();
 sg13g2_decap_4 FILLER_166_930 ();
 sg13g2_fill_2 FILLER_166_934 ();
 sg13g2_fill_2 FILLER_166_948 ();
 sg13g2_fill_1 FILLER_166_954 ();
 sg13g2_fill_1 FILLER_166_960 ();
 sg13g2_fill_2 FILLER_166_966 ();
 sg13g2_fill_1 FILLER_166_980 ();
 sg13g2_fill_2 FILLER_166_991 ();
 sg13g2_fill_2 FILLER_166_997 ();
 sg13g2_decap_8 FILLER_166_1025 ();
 sg13g2_decap_8 FILLER_166_1032 ();
 sg13g2_decap_4 FILLER_166_1039 ();
 sg13g2_fill_1 FILLER_166_1043 ();
 sg13g2_decap_8 FILLER_166_1048 ();
 sg13g2_decap_8 FILLER_166_1055 ();
 sg13g2_decap_4 FILLER_166_1062 ();
 sg13g2_fill_2 FILLER_166_1066 ();
 sg13g2_decap_8 FILLER_166_1094 ();
 sg13g2_decap_8 FILLER_166_1101 ();
 sg13g2_fill_2 FILLER_166_1108 ();
 sg13g2_decap_8 FILLER_166_1144 ();
 sg13g2_decap_8 FILLER_166_1261 ();
 sg13g2_decap_8 FILLER_166_1268 ();
 sg13g2_decap_8 FILLER_166_1275 ();
 sg13g2_decap_8 FILLER_166_1282 ();
 sg13g2_fill_1 FILLER_166_1289 ();
 sg13g2_fill_1 FILLER_166_1302 ();
 sg13g2_decap_4 FILLER_166_1307 ();
 sg13g2_decap_8 FILLER_166_1337 ();
 sg13g2_decap_8 FILLER_166_1344 ();
 sg13g2_decap_8 FILLER_166_1351 ();
 sg13g2_decap_8 FILLER_166_1358 ();
 sg13g2_decap_8 FILLER_166_1365 ();
 sg13g2_decap_8 FILLER_166_1372 ();
 sg13g2_decap_8 FILLER_166_1379 ();
 sg13g2_decap_8 FILLER_166_1386 ();
 sg13g2_decap_8 FILLER_166_1393 ();
 sg13g2_decap_8 FILLER_166_1400 ();
 sg13g2_decap_8 FILLER_166_1407 ();
 sg13g2_decap_8 FILLER_166_1414 ();
 sg13g2_decap_8 FILLER_166_1421 ();
 sg13g2_decap_8 FILLER_166_1428 ();
 sg13g2_decap_8 FILLER_166_1435 ();
 sg13g2_decap_8 FILLER_166_1442 ();
 sg13g2_decap_8 FILLER_166_1449 ();
 sg13g2_decap_8 FILLER_166_1456 ();
 sg13g2_decap_8 FILLER_166_1463 ();
 sg13g2_decap_8 FILLER_166_1470 ();
 sg13g2_decap_8 FILLER_166_1477 ();
 sg13g2_decap_8 FILLER_166_1484 ();
 sg13g2_decap_8 FILLER_166_1491 ();
 sg13g2_decap_8 FILLER_166_1498 ();
 sg13g2_decap_8 FILLER_166_1505 ();
 sg13g2_decap_8 FILLER_166_1512 ();
 sg13g2_decap_8 FILLER_166_1519 ();
 sg13g2_decap_8 FILLER_166_1526 ();
 sg13g2_decap_8 FILLER_166_1533 ();
 sg13g2_decap_8 FILLER_166_1540 ();
 sg13g2_decap_8 FILLER_166_1547 ();
 sg13g2_decap_8 FILLER_166_1554 ();
 sg13g2_decap_8 FILLER_166_1561 ();
 sg13g2_decap_8 FILLER_166_1568 ();
 sg13g2_decap_8 FILLER_166_1575 ();
 sg13g2_decap_8 FILLER_166_1582 ();
 sg13g2_decap_8 FILLER_166_1589 ();
 sg13g2_decap_8 FILLER_166_1596 ();
 sg13g2_decap_8 FILLER_166_1603 ();
 sg13g2_decap_8 FILLER_166_1610 ();
 sg13g2_decap_8 FILLER_166_1617 ();
 sg13g2_fill_1 FILLER_166_1624 ();
 sg13g2_decap_8 FILLER_167_0 ();
 sg13g2_decap_8 FILLER_167_7 ();
 sg13g2_decap_8 FILLER_167_14 ();
 sg13g2_decap_8 FILLER_167_21 ();
 sg13g2_decap_8 FILLER_167_28 ();
 sg13g2_decap_8 FILLER_167_35 ();
 sg13g2_decap_8 FILLER_167_42 ();
 sg13g2_decap_8 FILLER_167_49 ();
 sg13g2_decap_8 FILLER_167_56 ();
 sg13g2_decap_8 FILLER_167_63 ();
 sg13g2_decap_8 FILLER_167_70 ();
 sg13g2_decap_8 FILLER_167_77 ();
 sg13g2_decap_8 FILLER_167_84 ();
 sg13g2_decap_8 FILLER_167_91 ();
 sg13g2_decap_8 FILLER_167_98 ();
 sg13g2_decap_8 FILLER_167_105 ();
 sg13g2_decap_8 FILLER_167_112 ();
 sg13g2_decap_8 FILLER_167_119 ();
 sg13g2_decap_8 FILLER_167_126 ();
 sg13g2_decap_8 FILLER_167_133 ();
 sg13g2_decap_8 FILLER_167_140 ();
 sg13g2_decap_8 FILLER_167_147 ();
 sg13g2_decap_8 FILLER_167_154 ();
 sg13g2_fill_2 FILLER_167_161 ();
 sg13g2_decap_8 FILLER_167_172 ();
 sg13g2_decap_8 FILLER_167_179 ();
 sg13g2_decap_4 FILLER_167_186 ();
 sg13g2_decap_8 FILLER_167_224 ();
 sg13g2_decap_8 FILLER_167_231 ();
 sg13g2_decap_4 FILLER_167_238 ();
 sg13g2_decap_8 FILLER_167_268 ();
 sg13g2_decap_8 FILLER_167_275 ();
 sg13g2_decap_4 FILLER_167_299 ();
 sg13g2_fill_1 FILLER_167_303 ();
 sg13g2_fill_2 FILLER_167_315 ();
 sg13g2_decap_8 FILLER_167_321 ();
 sg13g2_fill_2 FILLER_167_333 ();
 sg13g2_fill_1 FILLER_167_335 ();
 sg13g2_fill_2 FILLER_167_340 ();
 sg13g2_fill_1 FILLER_167_342 ();
 sg13g2_decap_8 FILLER_167_373 ();
 sg13g2_decap_4 FILLER_167_380 ();
 sg13g2_fill_1 FILLER_167_384 ();
 sg13g2_decap_4 FILLER_167_419 ();
 sg13g2_decap_4 FILLER_167_428 ();
 sg13g2_fill_1 FILLER_167_432 ();
 sg13g2_decap_4 FILLER_167_437 ();
 sg13g2_fill_1 FILLER_167_441 ();
 sg13g2_decap_4 FILLER_167_481 ();
 sg13g2_fill_1 FILLER_167_485 ();
 sg13g2_decap_8 FILLER_167_512 ();
 sg13g2_decap_8 FILLER_167_519 ();
 sg13g2_decap_8 FILLER_167_526 ();
 sg13g2_decap_8 FILLER_167_533 ();
 sg13g2_decap_4 FILLER_167_540 ();
 sg13g2_decap_8 FILLER_167_558 ();
 sg13g2_fill_2 FILLER_167_565 ();
 sg13g2_fill_1 FILLER_167_567 ();
 sg13g2_fill_1 FILLER_167_594 ();
 sg13g2_decap_4 FILLER_167_651 ();
 sg13g2_decap_8 FILLER_167_660 ();
 sg13g2_fill_1 FILLER_167_667 ();
 sg13g2_decap_8 FILLER_167_723 ();
 sg13g2_decap_4 FILLER_167_730 ();
 sg13g2_fill_2 FILLER_167_734 ();
 sg13g2_decap_8 FILLER_167_749 ();
 sg13g2_fill_1 FILLER_167_756 ();
 sg13g2_decap_8 FILLER_167_845 ();
 sg13g2_decap_8 FILLER_167_852 ();
 sg13g2_fill_2 FILLER_167_859 ();
 sg13g2_fill_2 FILLER_167_865 ();
 sg13g2_fill_1 FILLER_167_867 ();
 sg13g2_decap_8 FILLER_167_878 ();
 sg13g2_decap_8 FILLER_167_885 ();
 sg13g2_fill_2 FILLER_167_892 ();
 sg13g2_decap_8 FILLER_167_898 ();
 sg13g2_fill_2 FILLER_167_905 ();
 sg13g2_fill_1 FILLER_167_907 ();
 sg13g2_decap_4 FILLER_167_919 ();
 sg13g2_decap_4 FILLER_167_930 ();
 sg13g2_decap_8 FILLER_167_988 ();
 sg13g2_decap_8 FILLER_167_995 ();
 sg13g2_decap_8 FILLER_167_1002 ();
 sg13g2_decap_8 FILLER_167_1009 ();
 sg13g2_fill_2 FILLER_167_1016 ();
 sg13g2_decap_8 FILLER_167_1022 ();
 sg13g2_fill_1 FILLER_167_1032 ();
 sg13g2_decap_8 FILLER_167_1063 ();
 sg13g2_decap_8 FILLER_167_1070 ();
 sg13g2_fill_2 FILLER_167_1077 ();
 sg13g2_fill_1 FILLER_167_1079 ();
 sg13g2_decap_4 FILLER_167_1088 ();
 sg13g2_fill_2 FILLER_167_1092 ();
 sg13g2_fill_1 FILLER_167_1194 ();
 sg13g2_fill_2 FILLER_167_1249 ();
 sg13g2_fill_1 FILLER_167_1251 ();
 sg13g2_decap_8 FILLER_167_1258 ();
 sg13g2_decap_4 FILLER_167_1277 ();
 sg13g2_decap_8 FILLER_167_1286 ();
 sg13g2_decap_8 FILLER_167_1297 ();
 sg13g2_fill_1 FILLER_167_1304 ();
 sg13g2_decap_8 FILLER_167_1309 ();
 sg13g2_decap_8 FILLER_167_1316 ();
 sg13g2_decap_8 FILLER_167_1323 ();
 sg13g2_decap_8 FILLER_167_1330 ();
 sg13g2_decap_8 FILLER_167_1337 ();
 sg13g2_decap_8 FILLER_167_1344 ();
 sg13g2_decap_8 FILLER_167_1351 ();
 sg13g2_decap_8 FILLER_167_1358 ();
 sg13g2_decap_8 FILLER_167_1365 ();
 sg13g2_decap_8 FILLER_167_1372 ();
 sg13g2_decap_8 FILLER_167_1379 ();
 sg13g2_decap_8 FILLER_167_1386 ();
 sg13g2_decap_8 FILLER_167_1393 ();
 sg13g2_decap_8 FILLER_167_1400 ();
 sg13g2_decap_8 FILLER_167_1407 ();
 sg13g2_decap_8 FILLER_167_1414 ();
 sg13g2_decap_8 FILLER_167_1421 ();
 sg13g2_decap_8 FILLER_167_1428 ();
 sg13g2_decap_8 FILLER_167_1435 ();
 sg13g2_decap_8 FILLER_167_1442 ();
 sg13g2_decap_8 FILLER_167_1449 ();
 sg13g2_decap_8 FILLER_167_1456 ();
 sg13g2_decap_8 FILLER_167_1463 ();
 sg13g2_decap_8 FILLER_167_1470 ();
 sg13g2_decap_8 FILLER_167_1477 ();
 sg13g2_decap_8 FILLER_167_1484 ();
 sg13g2_decap_8 FILLER_167_1491 ();
 sg13g2_decap_8 FILLER_167_1498 ();
 sg13g2_decap_8 FILLER_167_1505 ();
 sg13g2_decap_8 FILLER_167_1512 ();
 sg13g2_decap_8 FILLER_167_1519 ();
 sg13g2_decap_8 FILLER_167_1526 ();
 sg13g2_decap_8 FILLER_167_1533 ();
 sg13g2_decap_8 FILLER_167_1540 ();
 sg13g2_decap_8 FILLER_167_1547 ();
 sg13g2_decap_8 FILLER_167_1554 ();
 sg13g2_decap_8 FILLER_167_1561 ();
 sg13g2_decap_8 FILLER_167_1568 ();
 sg13g2_decap_8 FILLER_167_1575 ();
 sg13g2_decap_8 FILLER_167_1582 ();
 sg13g2_decap_8 FILLER_167_1589 ();
 sg13g2_decap_8 FILLER_167_1596 ();
 sg13g2_decap_8 FILLER_167_1603 ();
 sg13g2_decap_8 FILLER_167_1610 ();
 sg13g2_decap_8 FILLER_167_1617 ();
 sg13g2_fill_1 FILLER_167_1624 ();
 sg13g2_decap_8 FILLER_168_0 ();
 sg13g2_decap_8 FILLER_168_7 ();
 sg13g2_decap_8 FILLER_168_14 ();
 sg13g2_decap_8 FILLER_168_21 ();
 sg13g2_decap_8 FILLER_168_28 ();
 sg13g2_decap_8 FILLER_168_35 ();
 sg13g2_decap_8 FILLER_168_42 ();
 sg13g2_decap_8 FILLER_168_49 ();
 sg13g2_decap_8 FILLER_168_56 ();
 sg13g2_decap_8 FILLER_168_63 ();
 sg13g2_decap_8 FILLER_168_70 ();
 sg13g2_decap_8 FILLER_168_77 ();
 sg13g2_decap_8 FILLER_168_84 ();
 sg13g2_decap_8 FILLER_168_91 ();
 sg13g2_decap_8 FILLER_168_98 ();
 sg13g2_decap_8 FILLER_168_105 ();
 sg13g2_decap_8 FILLER_168_112 ();
 sg13g2_decap_8 FILLER_168_119 ();
 sg13g2_fill_1 FILLER_168_126 ();
 sg13g2_decap_8 FILLER_168_131 ();
 sg13g2_decap_8 FILLER_168_138 ();
 sg13g2_decap_8 FILLER_168_145 ();
 sg13g2_decap_4 FILLER_168_152 ();
 sg13g2_decap_4 FILLER_168_169 ();
 sg13g2_fill_1 FILLER_168_173 ();
 sg13g2_fill_1 FILLER_168_192 ();
 sg13g2_decap_8 FILLER_168_202 ();
 sg13g2_decap_4 FILLER_168_209 ();
 sg13g2_decap_4 FILLER_168_243 ();
 sg13g2_decap_8 FILLER_168_258 ();
 sg13g2_fill_2 FILLER_168_265 ();
 sg13g2_fill_1 FILLER_168_267 ();
 sg13g2_fill_1 FILLER_168_280 ();
 sg13g2_fill_1 FILLER_168_335 ();
 sg13g2_decap_8 FILLER_168_371 ();
 sg13g2_decap_8 FILLER_168_378 ();
 sg13g2_decap_8 FILLER_168_385 ();
 sg13g2_fill_2 FILLER_168_392 ();
 sg13g2_decap_8 FILLER_168_476 ();
 sg13g2_decap_8 FILLER_168_483 ();
 sg13g2_decap_8 FILLER_168_490 ();
 sg13g2_decap_8 FILLER_168_497 ();
 sg13g2_decap_8 FILLER_168_504 ();
 sg13g2_decap_8 FILLER_168_583 ();
 sg13g2_fill_1 FILLER_168_590 ();
 sg13g2_decap_8 FILLER_168_619 ();
 sg13g2_fill_1 FILLER_168_626 ();
 sg13g2_decap_8 FILLER_168_693 ();
 sg13g2_fill_2 FILLER_168_700 ();
 sg13g2_fill_1 FILLER_168_702 ();
 sg13g2_fill_2 FILLER_168_708 ();
 sg13g2_fill_2 FILLER_168_715 ();
 sg13g2_decap_4 FILLER_168_725 ();
 sg13g2_fill_2 FILLER_168_734 ();
 sg13g2_fill_2 FILLER_168_741 ();
 sg13g2_fill_1 FILLER_168_743 ();
 sg13g2_decap_8 FILLER_168_752 ();
 sg13g2_decap_8 FILLER_168_759 ();
 sg13g2_decap_4 FILLER_168_766 ();
 sg13g2_fill_2 FILLER_168_774 ();
 sg13g2_decap_8 FILLER_168_782 ();
 sg13g2_decap_8 FILLER_168_789 ();
 sg13g2_decap_4 FILLER_168_796 ();
 sg13g2_fill_2 FILLER_168_800 ();
 sg13g2_fill_1 FILLER_168_806 ();
 sg13g2_decap_8 FILLER_168_833 ();
 sg13g2_fill_2 FILLER_168_844 ();
 sg13g2_fill_2 FILLER_168_850 ();
 sg13g2_fill_1 FILLER_168_852 ();
 sg13g2_fill_2 FILLER_168_861 ();
 sg13g2_fill_2 FILLER_168_882 ();
 sg13g2_decap_8 FILLER_168_926 ();
 sg13g2_decap_4 FILLER_168_933 ();
 sg13g2_decap_4 FILLER_168_968 ();
 sg13g2_fill_2 FILLER_168_976 ();
 sg13g2_decap_4 FILLER_168_982 ();
 sg13g2_decap_8 FILLER_168_990 ();
 sg13g2_decap_8 FILLER_168_997 ();
 sg13g2_decap_8 FILLER_168_1004 ();
 sg13g2_fill_1 FILLER_168_1011 ();
 sg13g2_fill_2 FILLER_168_1055 ();
 sg13g2_fill_1 FILLER_168_1057 ();
 sg13g2_fill_2 FILLER_168_1063 ();
 sg13g2_fill_1 FILLER_168_1065 ();
 sg13g2_decap_4 FILLER_168_1073 ();
 sg13g2_fill_2 FILLER_168_1077 ();
 sg13g2_fill_1 FILLER_168_1109 ();
 sg13g2_fill_2 FILLER_168_1157 ();
 sg13g2_decap_4 FILLER_168_1163 ();
 sg13g2_fill_2 FILLER_168_1196 ();
 sg13g2_fill_1 FILLER_168_1198 ();
 sg13g2_decap_4 FILLER_168_1242 ();
 sg13g2_fill_1 FILLER_168_1246 ();
 sg13g2_fill_2 FILLER_168_1253 ();
 sg13g2_fill_1 FILLER_168_1255 ();
 sg13g2_fill_2 FILLER_168_1268 ();
 sg13g2_fill_1 FILLER_168_1270 ();
 sg13g2_decap_8 FILLER_168_1277 ();
 sg13g2_fill_1 FILLER_168_1296 ();
 sg13g2_decap_8 FILLER_168_1323 ();
 sg13g2_decap_8 FILLER_168_1330 ();
 sg13g2_decap_8 FILLER_168_1337 ();
 sg13g2_decap_8 FILLER_168_1344 ();
 sg13g2_decap_8 FILLER_168_1351 ();
 sg13g2_decap_8 FILLER_168_1358 ();
 sg13g2_decap_8 FILLER_168_1365 ();
 sg13g2_decap_8 FILLER_168_1372 ();
 sg13g2_decap_8 FILLER_168_1379 ();
 sg13g2_decap_8 FILLER_168_1386 ();
 sg13g2_decap_8 FILLER_168_1393 ();
 sg13g2_decap_8 FILLER_168_1400 ();
 sg13g2_decap_8 FILLER_168_1407 ();
 sg13g2_decap_8 FILLER_168_1414 ();
 sg13g2_decap_8 FILLER_168_1421 ();
 sg13g2_decap_8 FILLER_168_1428 ();
 sg13g2_decap_8 FILLER_168_1435 ();
 sg13g2_decap_8 FILLER_168_1442 ();
 sg13g2_decap_8 FILLER_168_1449 ();
 sg13g2_decap_8 FILLER_168_1456 ();
 sg13g2_decap_8 FILLER_168_1463 ();
 sg13g2_decap_8 FILLER_168_1470 ();
 sg13g2_decap_8 FILLER_168_1477 ();
 sg13g2_decap_8 FILLER_168_1484 ();
 sg13g2_decap_8 FILLER_168_1491 ();
 sg13g2_decap_8 FILLER_168_1498 ();
 sg13g2_decap_8 FILLER_168_1505 ();
 sg13g2_decap_8 FILLER_168_1512 ();
 sg13g2_decap_8 FILLER_168_1519 ();
 sg13g2_decap_8 FILLER_168_1526 ();
 sg13g2_decap_8 FILLER_168_1533 ();
 sg13g2_decap_8 FILLER_168_1540 ();
 sg13g2_decap_8 FILLER_168_1547 ();
 sg13g2_decap_8 FILLER_168_1554 ();
 sg13g2_decap_8 FILLER_168_1561 ();
 sg13g2_decap_8 FILLER_168_1568 ();
 sg13g2_decap_8 FILLER_168_1575 ();
 sg13g2_decap_8 FILLER_168_1582 ();
 sg13g2_decap_8 FILLER_168_1589 ();
 sg13g2_decap_8 FILLER_168_1596 ();
 sg13g2_decap_8 FILLER_168_1603 ();
 sg13g2_decap_8 FILLER_168_1610 ();
 sg13g2_decap_8 FILLER_168_1617 ();
 sg13g2_fill_1 FILLER_168_1624 ();
 sg13g2_decap_8 FILLER_169_0 ();
 sg13g2_decap_8 FILLER_169_7 ();
 sg13g2_decap_8 FILLER_169_14 ();
 sg13g2_decap_8 FILLER_169_21 ();
 sg13g2_decap_8 FILLER_169_28 ();
 sg13g2_decap_8 FILLER_169_35 ();
 sg13g2_decap_8 FILLER_169_42 ();
 sg13g2_decap_8 FILLER_169_49 ();
 sg13g2_decap_8 FILLER_169_56 ();
 sg13g2_decap_8 FILLER_169_63 ();
 sg13g2_decap_8 FILLER_169_70 ();
 sg13g2_decap_8 FILLER_169_77 ();
 sg13g2_decap_8 FILLER_169_84 ();
 sg13g2_decap_8 FILLER_169_91 ();
 sg13g2_decap_8 FILLER_169_98 ();
 sg13g2_decap_8 FILLER_169_105 ();
 sg13g2_fill_2 FILLER_169_112 ();
 sg13g2_fill_2 FILLER_169_119 ();
 sg13g2_decap_4 FILLER_169_147 ();
 sg13g2_fill_2 FILLER_169_151 ();
 sg13g2_decap_8 FILLER_169_158 ();
 sg13g2_decap_8 FILLER_169_165 ();
 sg13g2_decap_4 FILLER_169_172 ();
 sg13g2_fill_2 FILLER_169_176 ();
 sg13g2_fill_2 FILLER_169_191 ();
 sg13g2_fill_2 FILLER_169_293 ();
 sg13g2_fill_1 FILLER_169_295 ();
 sg13g2_fill_2 FILLER_169_300 ();
 sg13g2_fill_1 FILLER_169_312 ();
 sg13g2_decap_8 FILLER_169_317 ();
 sg13g2_decap_4 FILLER_169_334 ();
 sg13g2_decap_8 FILLER_169_343 ();
 sg13g2_decap_8 FILLER_169_350 ();
 sg13g2_decap_8 FILLER_169_357 ();
 sg13g2_fill_2 FILLER_169_364 ();
 sg13g2_fill_1 FILLER_169_366 ();
 sg13g2_decap_8 FILLER_169_373 ();
 sg13g2_decap_8 FILLER_169_380 ();
 sg13g2_decap_4 FILLER_169_387 ();
 sg13g2_decap_4 FILLER_169_397 ();
 sg13g2_fill_1 FILLER_169_401 ();
 sg13g2_fill_2 FILLER_169_431 ();
 sg13g2_fill_1 FILLER_169_433 ();
 sg13g2_fill_1 FILLER_169_458 ();
 sg13g2_decap_8 FILLER_169_465 ();
 sg13g2_decap_8 FILLER_169_472 ();
 sg13g2_fill_2 FILLER_169_479 ();
 sg13g2_fill_1 FILLER_169_481 ();
 sg13g2_fill_1 FILLER_169_486 ();
 sg13g2_decap_8 FILLER_169_491 ();
 sg13g2_decap_8 FILLER_169_498 ();
 sg13g2_decap_8 FILLER_169_505 ();
 sg13g2_decap_8 FILLER_169_512 ();
 sg13g2_decap_8 FILLER_169_519 ();
 sg13g2_fill_2 FILLER_169_526 ();
 sg13g2_fill_1 FILLER_169_528 ();
 sg13g2_fill_1 FILLER_169_533 ();
 sg13g2_decap_8 FILLER_169_541 ();
 sg13g2_decap_8 FILLER_169_548 ();
 sg13g2_decap_8 FILLER_169_555 ();
 sg13g2_decap_8 FILLER_169_562 ();
 sg13g2_decap_8 FILLER_169_569 ();
 sg13g2_decap_8 FILLER_169_576 ();
 sg13g2_fill_2 FILLER_169_583 ();
 sg13g2_fill_1 FILLER_169_585 ();
 sg13g2_decap_8 FILLER_169_590 ();
 sg13g2_fill_2 FILLER_169_597 ();
 sg13g2_fill_1 FILLER_169_599 ();
 sg13g2_fill_1 FILLER_169_613 ();
 sg13g2_decap_8 FILLER_169_618 ();
 sg13g2_decap_4 FILLER_169_625 ();
 sg13g2_decap_8 FILLER_169_665 ();
 sg13g2_decap_8 FILLER_169_672 ();
 sg13g2_decap_8 FILLER_169_679 ();
 sg13g2_decap_8 FILLER_169_686 ();
 sg13g2_decap_8 FILLER_169_693 ();
 sg13g2_decap_8 FILLER_169_700 ();
 sg13g2_fill_1 FILLER_169_707 ();
 sg13g2_fill_1 FILLER_169_733 ();
 sg13g2_fill_1 FILLER_169_743 ();
 sg13g2_fill_2 FILLER_169_754 ();
 sg13g2_fill_1 FILLER_169_783 ();
 sg13g2_decap_8 FILLER_169_788 ();
 sg13g2_fill_2 FILLER_169_795 ();
 sg13g2_decap_8 FILLER_169_809 ();
 sg13g2_fill_1 FILLER_169_820 ();
 sg13g2_decap_8 FILLER_169_825 ();
 sg13g2_fill_1 FILLER_169_832 ();
 sg13g2_fill_2 FILLER_169_859 ();
 sg13g2_fill_1 FILLER_169_869 ();
 sg13g2_decap_8 FILLER_169_875 ();
 sg13g2_fill_2 FILLER_169_882 ();
 sg13g2_decap_8 FILLER_169_925 ();
 sg13g2_decap_8 FILLER_169_932 ();
 sg13g2_decap_8 FILLER_169_939 ();
 sg13g2_decap_8 FILLER_169_946 ();
 sg13g2_decap_8 FILLER_169_953 ();
 sg13g2_decap_8 FILLER_169_960 ();
 sg13g2_decap_8 FILLER_169_967 ();
 sg13g2_decap_4 FILLER_169_1009 ();
 sg13g2_fill_1 FILLER_169_1013 ();
 sg13g2_fill_2 FILLER_169_1026 ();
 sg13g2_fill_1 FILLER_169_1028 ();
 sg13g2_decap_4 FILLER_169_1054 ();
 sg13g2_fill_2 FILLER_169_1058 ();
 sg13g2_fill_1 FILLER_169_1064 ();
 sg13g2_decap_8 FILLER_169_1071 ();
 sg13g2_decap_8 FILLER_169_1078 ();
 sg13g2_decap_4 FILLER_169_1085 ();
 sg13g2_fill_1 FILLER_169_1089 ();
 sg13g2_fill_2 FILLER_169_1094 ();
 sg13g2_fill_1 FILLER_169_1104 ();
 sg13g2_fill_2 FILLER_169_1156 ();
 sg13g2_fill_1 FILLER_169_1158 ();
 sg13g2_decap_8 FILLER_169_1163 ();
 sg13g2_fill_2 FILLER_169_1170 ();
 sg13g2_fill_1 FILLER_169_1172 ();
 sg13g2_fill_1 FILLER_169_1209 ();
 sg13g2_decap_4 FILLER_169_1244 ();
 sg13g2_decap_4 FILLER_169_1252 ();
 sg13g2_decap_4 FILLER_169_1264 ();
 sg13g2_fill_2 FILLER_169_1280 ();
 sg13g2_decap_8 FILLER_169_1324 ();
 sg13g2_decap_8 FILLER_169_1331 ();
 sg13g2_decap_8 FILLER_169_1338 ();
 sg13g2_decap_8 FILLER_169_1345 ();
 sg13g2_decap_8 FILLER_169_1352 ();
 sg13g2_decap_8 FILLER_169_1359 ();
 sg13g2_decap_8 FILLER_169_1366 ();
 sg13g2_decap_8 FILLER_169_1373 ();
 sg13g2_decap_8 FILLER_169_1380 ();
 sg13g2_decap_8 FILLER_169_1387 ();
 sg13g2_decap_8 FILLER_169_1394 ();
 sg13g2_decap_8 FILLER_169_1401 ();
 sg13g2_decap_8 FILLER_169_1408 ();
 sg13g2_decap_8 FILLER_169_1415 ();
 sg13g2_decap_8 FILLER_169_1422 ();
 sg13g2_decap_8 FILLER_169_1429 ();
 sg13g2_decap_8 FILLER_169_1436 ();
 sg13g2_decap_8 FILLER_169_1443 ();
 sg13g2_decap_8 FILLER_169_1450 ();
 sg13g2_decap_8 FILLER_169_1457 ();
 sg13g2_decap_8 FILLER_169_1464 ();
 sg13g2_decap_8 FILLER_169_1471 ();
 sg13g2_decap_8 FILLER_169_1478 ();
 sg13g2_decap_8 FILLER_169_1485 ();
 sg13g2_decap_8 FILLER_169_1492 ();
 sg13g2_decap_8 FILLER_169_1499 ();
 sg13g2_decap_8 FILLER_169_1506 ();
 sg13g2_decap_8 FILLER_169_1513 ();
 sg13g2_decap_8 FILLER_169_1520 ();
 sg13g2_decap_8 FILLER_169_1527 ();
 sg13g2_decap_8 FILLER_169_1534 ();
 sg13g2_decap_8 FILLER_169_1541 ();
 sg13g2_decap_8 FILLER_169_1548 ();
 sg13g2_decap_8 FILLER_169_1555 ();
 sg13g2_decap_8 FILLER_169_1562 ();
 sg13g2_decap_8 FILLER_169_1569 ();
 sg13g2_decap_8 FILLER_169_1576 ();
 sg13g2_decap_8 FILLER_169_1583 ();
 sg13g2_decap_8 FILLER_169_1590 ();
 sg13g2_decap_8 FILLER_169_1597 ();
 sg13g2_decap_8 FILLER_169_1604 ();
 sg13g2_decap_8 FILLER_169_1611 ();
 sg13g2_decap_8 FILLER_169_1618 ();
 sg13g2_decap_8 FILLER_170_0 ();
 sg13g2_decap_8 FILLER_170_7 ();
 sg13g2_decap_8 FILLER_170_14 ();
 sg13g2_decap_8 FILLER_170_21 ();
 sg13g2_decap_8 FILLER_170_28 ();
 sg13g2_decap_8 FILLER_170_35 ();
 sg13g2_decap_8 FILLER_170_42 ();
 sg13g2_decap_8 FILLER_170_49 ();
 sg13g2_decap_8 FILLER_170_56 ();
 sg13g2_decap_8 FILLER_170_63 ();
 sg13g2_decap_8 FILLER_170_70 ();
 sg13g2_decap_8 FILLER_170_77 ();
 sg13g2_decap_8 FILLER_170_84 ();
 sg13g2_decap_8 FILLER_170_91 ();
 sg13g2_decap_8 FILLER_170_98 ();
 sg13g2_decap_8 FILLER_170_105 ();
 sg13g2_fill_1 FILLER_170_112 ();
 sg13g2_decap_8 FILLER_170_167 ();
 sg13g2_fill_1 FILLER_170_174 ();
 sg13g2_decap_4 FILLER_170_188 ();
 sg13g2_decap_4 FILLER_170_222 ();
 sg13g2_fill_1 FILLER_170_252 ();
 sg13g2_decap_4 FILLER_170_301 ();
 sg13g2_fill_2 FILLER_170_305 ();
 sg13g2_fill_1 FILLER_170_356 ();
 sg13g2_decap_4 FILLER_170_368 ();
 sg13g2_fill_1 FILLER_170_372 ();
 sg13g2_decap_8 FILLER_170_381 ();
 sg13g2_fill_1 FILLER_170_388 ();
 sg13g2_fill_2 FILLER_170_400 ();
 sg13g2_decap_8 FILLER_170_406 ();
 sg13g2_decap_4 FILLER_170_413 ();
 sg13g2_fill_1 FILLER_170_417 ();
 sg13g2_fill_2 FILLER_170_426 ();
 sg13g2_fill_1 FILLER_170_428 ();
 sg13g2_fill_2 FILLER_170_433 ();
 sg13g2_decap_8 FILLER_170_444 ();
 sg13g2_decap_8 FILLER_170_451 ();
 sg13g2_decap_8 FILLER_170_458 ();
 sg13g2_decap_4 FILLER_170_465 ();
 sg13g2_fill_2 FILLER_170_469 ();
 sg13g2_decap_4 FILLER_170_507 ();
 sg13g2_decap_8 FILLER_170_515 ();
 sg13g2_fill_2 FILLER_170_522 ();
 sg13g2_fill_1 FILLER_170_524 ();
 sg13g2_fill_1 FILLER_170_535 ();
 sg13g2_fill_1 FILLER_170_546 ();
 sg13g2_fill_1 FILLER_170_557 ();
 sg13g2_decap_4 FILLER_170_562 ();
 sg13g2_fill_2 FILLER_170_566 ();
 sg13g2_fill_2 FILLER_170_604 ();
 sg13g2_fill_1 FILLER_170_642 ();
 sg13g2_decap_8 FILLER_170_647 ();
 sg13g2_decap_8 FILLER_170_654 ();
 sg13g2_fill_2 FILLER_170_661 ();
 sg13g2_fill_2 FILLER_170_673 ();
 sg13g2_decap_8 FILLER_170_679 ();
 sg13g2_decap_8 FILLER_170_686 ();
 sg13g2_fill_2 FILLER_170_693 ();
 sg13g2_fill_1 FILLER_170_705 ();
 sg13g2_decap_4 FILLER_170_736 ();
 sg13g2_decap_8 FILLER_170_754 ();
 sg13g2_decap_8 FILLER_170_761 ();
 sg13g2_decap_8 FILLER_170_768 ();
 sg13g2_fill_1 FILLER_170_775 ();
 sg13g2_fill_2 FILLER_170_838 ();
 sg13g2_decap_8 FILLER_170_870 ();
 sg13g2_decap_8 FILLER_170_877 ();
 sg13g2_decap_4 FILLER_170_884 ();
 sg13g2_decap_4 FILLER_170_929 ();
 sg13g2_fill_1 FILLER_170_933 ();
 sg13g2_decap_8 FILLER_170_938 ();
 sg13g2_decap_8 FILLER_170_945 ();
 sg13g2_fill_2 FILLER_170_952 ();
 sg13g2_decap_8 FILLER_170_971 ();
 sg13g2_decap_8 FILLER_170_978 ();
 sg13g2_decap_4 FILLER_170_985 ();
 sg13g2_fill_2 FILLER_170_1017 ();
 sg13g2_fill_2 FILLER_170_1033 ();
 sg13g2_decap_4 FILLER_170_1040 ();
 sg13g2_fill_2 FILLER_170_1044 ();
 sg13g2_fill_2 FILLER_170_1052 ();
 sg13g2_fill_1 FILLER_170_1063 ();
 sg13g2_decap_8 FILLER_170_1073 ();
 sg13g2_decap_8 FILLER_170_1080 ();
 sg13g2_fill_1 FILLER_170_1138 ();
 sg13g2_fill_2 FILLER_170_1185 ();
 sg13g2_decap_8 FILLER_170_1196 ();
 sg13g2_decap_4 FILLER_170_1203 ();
 sg13g2_fill_2 FILLER_170_1207 ();
 sg13g2_decap_8 FILLER_170_1213 ();
 sg13g2_decap_8 FILLER_170_1220 ();
 sg13g2_decap_4 FILLER_170_1227 ();
 sg13g2_fill_2 FILLER_170_1231 ();
 sg13g2_decap_4 FILLER_170_1267 ();
 sg13g2_decap_8 FILLER_170_1279 ();
 sg13g2_fill_2 FILLER_170_1286 ();
 sg13g2_fill_1 FILLER_170_1288 ();
 sg13g2_decap_4 FILLER_170_1293 ();
 sg13g2_fill_1 FILLER_170_1297 ();
 sg13g2_decap_8 FILLER_170_1323 ();
 sg13g2_decap_8 FILLER_170_1330 ();
 sg13g2_decap_8 FILLER_170_1337 ();
 sg13g2_decap_8 FILLER_170_1344 ();
 sg13g2_decap_8 FILLER_170_1351 ();
 sg13g2_decap_8 FILLER_170_1358 ();
 sg13g2_decap_8 FILLER_170_1365 ();
 sg13g2_decap_8 FILLER_170_1372 ();
 sg13g2_decap_8 FILLER_170_1379 ();
 sg13g2_decap_8 FILLER_170_1386 ();
 sg13g2_decap_8 FILLER_170_1393 ();
 sg13g2_decap_8 FILLER_170_1400 ();
 sg13g2_decap_8 FILLER_170_1407 ();
 sg13g2_decap_8 FILLER_170_1414 ();
 sg13g2_decap_8 FILLER_170_1421 ();
 sg13g2_decap_8 FILLER_170_1428 ();
 sg13g2_decap_8 FILLER_170_1435 ();
 sg13g2_decap_8 FILLER_170_1442 ();
 sg13g2_decap_8 FILLER_170_1449 ();
 sg13g2_decap_8 FILLER_170_1456 ();
 sg13g2_decap_8 FILLER_170_1463 ();
 sg13g2_decap_8 FILLER_170_1470 ();
 sg13g2_decap_8 FILLER_170_1477 ();
 sg13g2_decap_8 FILLER_170_1484 ();
 sg13g2_decap_8 FILLER_170_1491 ();
 sg13g2_decap_8 FILLER_170_1498 ();
 sg13g2_decap_8 FILLER_170_1505 ();
 sg13g2_decap_8 FILLER_170_1512 ();
 sg13g2_decap_8 FILLER_170_1519 ();
 sg13g2_decap_8 FILLER_170_1526 ();
 sg13g2_decap_8 FILLER_170_1533 ();
 sg13g2_decap_8 FILLER_170_1540 ();
 sg13g2_decap_8 FILLER_170_1547 ();
 sg13g2_decap_8 FILLER_170_1554 ();
 sg13g2_decap_8 FILLER_170_1561 ();
 sg13g2_decap_8 FILLER_170_1568 ();
 sg13g2_decap_8 FILLER_170_1575 ();
 sg13g2_decap_8 FILLER_170_1582 ();
 sg13g2_decap_8 FILLER_170_1589 ();
 sg13g2_decap_8 FILLER_170_1596 ();
 sg13g2_decap_8 FILLER_170_1603 ();
 sg13g2_decap_8 FILLER_170_1610 ();
 sg13g2_decap_8 FILLER_170_1617 ();
 sg13g2_fill_1 FILLER_170_1624 ();
 sg13g2_decap_8 FILLER_171_0 ();
 sg13g2_decap_8 FILLER_171_7 ();
 sg13g2_decap_8 FILLER_171_14 ();
 sg13g2_decap_8 FILLER_171_21 ();
 sg13g2_decap_8 FILLER_171_28 ();
 sg13g2_decap_8 FILLER_171_35 ();
 sg13g2_decap_8 FILLER_171_42 ();
 sg13g2_decap_8 FILLER_171_49 ();
 sg13g2_decap_8 FILLER_171_56 ();
 sg13g2_decap_8 FILLER_171_63 ();
 sg13g2_decap_8 FILLER_171_70 ();
 sg13g2_decap_8 FILLER_171_77 ();
 sg13g2_decap_8 FILLER_171_84 ();
 sg13g2_decap_8 FILLER_171_91 ();
 sg13g2_decap_8 FILLER_171_98 ();
 sg13g2_decap_8 FILLER_171_105 ();
 sg13g2_decap_8 FILLER_171_112 ();
 sg13g2_decap_8 FILLER_171_119 ();
 sg13g2_fill_2 FILLER_171_126 ();
 sg13g2_fill_1 FILLER_171_128 ();
 sg13g2_fill_2 FILLER_171_139 ();
 sg13g2_fill_1 FILLER_171_141 ();
 sg13g2_decap_8 FILLER_171_172 ();
 sg13g2_decap_4 FILLER_171_179 ();
 sg13g2_fill_2 FILLER_171_183 ();
 sg13g2_decap_4 FILLER_171_190 ();
 sg13g2_fill_2 FILLER_171_194 ();
 sg13g2_decap_4 FILLER_171_200 ();
 sg13g2_fill_1 FILLER_171_204 ();
 sg13g2_decap_8 FILLER_171_209 ();
 sg13g2_fill_1 FILLER_171_216 ();
 sg13g2_decap_8 FILLER_171_270 ();
 sg13g2_decap_4 FILLER_171_277 ();
 sg13g2_fill_2 FILLER_171_281 ();
 sg13g2_decap_8 FILLER_171_292 ();
 sg13g2_decap_4 FILLER_171_299 ();
 sg13g2_fill_1 FILLER_171_368 ();
 sg13g2_fill_1 FILLER_171_421 ();
 sg13g2_decap_4 FILLER_171_448 ();
 sg13g2_decap_8 FILLER_171_456 ();
 sg13g2_decap_4 FILLER_171_463 ();
 sg13g2_fill_1 FILLER_171_467 ();
 sg13g2_fill_1 FILLER_171_473 ();
 sg13g2_decap_4 FILLER_171_499 ();
 sg13g2_fill_1 FILLER_171_594 ();
 sg13g2_fill_1 FILLER_171_634 ();
 sg13g2_decap_8 FILLER_171_661 ();
 sg13g2_fill_1 FILLER_171_694 ();
 sg13g2_decap_8 FILLER_171_710 ();
 sg13g2_decap_8 FILLER_171_717 ();
 sg13g2_decap_4 FILLER_171_724 ();
 sg13g2_decap_4 FILLER_171_764 ();
 sg13g2_fill_2 FILLER_171_768 ();
 sg13g2_decap_8 FILLER_171_780 ();
 sg13g2_decap_8 FILLER_171_787 ();
 sg13g2_decap_4 FILLER_171_794 ();
 sg13g2_decap_8 FILLER_171_802 ();
 sg13g2_fill_2 FILLER_171_809 ();
 sg13g2_decap_8 FILLER_171_836 ();
 sg13g2_fill_1 FILLER_171_843 ();
 sg13g2_decap_8 FILLER_171_879 ();
 sg13g2_fill_2 FILLER_171_886 ();
 sg13g2_decap_8 FILLER_171_892 ();
 sg13g2_decap_8 FILLER_171_899 ();
 sg13g2_decap_8 FILLER_171_906 ();
 sg13g2_decap_8 FILLER_171_913 ();
 sg13g2_decap_4 FILLER_171_920 ();
 sg13g2_fill_1 FILLER_171_962 ();
 sg13g2_fill_2 FILLER_171_993 ();
 sg13g2_fill_2 FILLER_171_1039 ();
 sg13g2_decap_8 FILLER_171_1046 ();
 sg13g2_decap_4 FILLER_171_1057 ();
 sg13g2_fill_1 FILLER_171_1061 ();
 sg13g2_decap_4 FILLER_171_1067 ();
 sg13g2_fill_1 FILLER_171_1071 ();
 sg13g2_decap_8 FILLER_171_1083 ();
 sg13g2_fill_2 FILLER_171_1116 ();
 sg13g2_fill_1 FILLER_171_1118 ();
 sg13g2_decap_4 FILLER_171_1140 ();
 sg13g2_fill_1 FILLER_171_1144 ();
 sg13g2_decap_8 FILLER_171_1149 ();
 sg13g2_decap_8 FILLER_171_1156 ();
 sg13g2_decap_8 FILLER_171_1163 ();
 sg13g2_decap_8 FILLER_171_1170 ();
 sg13g2_decap_8 FILLER_171_1177 ();
 sg13g2_decap_8 FILLER_171_1184 ();
 sg13g2_decap_4 FILLER_171_1191 ();
 sg13g2_fill_2 FILLER_171_1195 ();
 sg13g2_decap_8 FILLER_171_1205 ();
 sg13g2_fill_2 FILLER_171_1212 ();
 sg13g2_fill_1 FILLER_171_1214 ();
 sg13g2_fill_2 FILLER_171_1219 ();
 sg13g2_decap_8 FILLER_171_1255 ();
 sg13g2_decap_8 FILLER_171_1262 ();
 sg13g2_decap_8 FILLER_171_1269 ();
 sg13g2_fill_2 FILLER_171_1280 ();
 sg13g2_decap_8 FILLER_171_1312 ();
 sg13g2_decap_8 FILLER_171_1319 ();
 sg13g2_decap_8 FILLER_171_1326 ();
 sg13g2_decap_8 FILLER_171_1333 ();
 sg13g2_decap_8 FILLER_171_1340 ();
 sg13g2_decap_8 FILLER_171_1347 ();
 sg13g2_decap_8 FILLER_171_1354 ();
 sg13g2_decap_8 FILLER_171_1361 ();
 sg13g2_decap_8 FILLER_171_1368 ();
 sg13g2_decap_8 FILLER_171_1375 ();
 sg13g2_decap_8 FILLER_171_1382 ();
 sg13g2_decap_8 FILLER_171_1389 ();
 sg13g2_decap_8 FILLER_171_1396 ();
 sg13g2_decap_8 FILLER_171_1403 ();
 sg13g2_decap_8 FILLER_171_1410 ();
 sg13g2_decap_8 FILLER_171_1417 ();
 sg13g2_decap_8 FILLER_171_1424 ();
 sg13g2_decap_8 FILLER_171_1431 ();
 sg13g2_decap_8 FILLER_171_1438 ();
 sg13g2_decap_8 FILLER_171_1445 ();
 sg13g2_decap_8 FILLER_171_1452 ();
 sg13g2_decap_8 FILLER_171_1459 ();
 sg13g2_decap_8 FILLER_171_1466 ();
 sg13g2_decap_8 FILLER_171_1473 ();
 sg13g2_decap_8 FILLER_171_1480 ();
 sg13g2_decap_8 FILLER_171_1487 ();
 sg13g2_decap_8 FILLER_171_1494 ();
 sg13g2_decap_8 FILLER_171_1501 ();
 sg13g2_decap_8 FILLER_171_1508 ();
 sg13g2_decap_8 FILLER_171_1515 ();
 sg13g2_decap_8 FILLER_171_1522 ();
 sg13g2_decap_8 FILLER_171_1529 ();
 sg13g2_decap_8 FILLER_171_1536 ();
 sg13g2_decap_8 FILLER_171_1543 ();
 sg13g2_decap_8 FILLER_171_1550 ();
 sg13g2_decap_8 FILLER_171_1557 ();
 sg13g2_decap_8 FILLER_171_1564 ();
 sg13g2_decap_8 FILLER_171_1571 ();
 sg13g2_decap_8 FILLER_171_1578 ();
 sg13g2_decap_8 FILLER_171_1585 ();
 sg13g2_decap_8 FILLER_171_1592 ();
 sg13g2_decap_8 FILLER_171_1599 ();
 sg13g2_decap_8 FILLER_171_1606 ();
 sg13g2_decap_8 FILLER_171_1613 ();
 sg13g2_decap_4 FILLER_171_1620 ();
 sg13g2_fill_1 FILLER_171_1624 ();
 sg13g2_decap_8 FILLER_172_0 ();
 sg13g2_decap_8 FILLER_172_7 ();
 sg13g2_decap_8 FILLER_172_14 ();
 sg13g2_decap_8 FILLER_172_21 ();
 sg13g2_decap_8 FILLER_172_28 ();
 sg13g2_decap_8 FILLER_172_35 ();
 sg13g2_decap_8 FILLER_172_42 ();
 sg13g2_decap_8 FILLER_172_49 ();
 sg13g2_decap_8 FILLER_172_56 ();
 sg13g2_decap_8 FILLER_172_63 ();
 sg13g2_decap_8 FILLER_172_70 ();
 sg13g2_decap_8 FILLER_172_77 ();
 sg13g2_decap_8 FILLER_172_84 ();
 sg13g2_decap_8 FILLER_172_91 ();
 sg13g2_decap_8 FILLER_172_98 ();
 sg13g2_decap_8 FILLER_172_105 ();
 sg13g2_decap_8 FILLER_172_112 ();
 sg13g2_decap_8 FILLER_172_119 ();
 sg13g2_decap_8 FILLER_172_126 ();
 sg13g2_decap_8 FILLER_172_133 ();
 sg13g2_decap_8 FILLER_172_140 ();
 sg13g2_decap_8 FILLER_172_147 ();
 sg13g2_decap_8 FILLER_172_154 ();
 sg13g2_decap_8 FILLER_172_161 ();
 sg13g2_decap_8 FILLER_172_168 ();
 sg13g2_decap_8 FILLER_172_175 ();
 sg13g2_decap_8 FILLER_172_182 ();
 sg13g2_decap_4 FILLER_172_189 ();
 sg13g2_decap_8 FILLER_172_197 ();
 sg13g2_decap_8 FILLER_172_204 ();
 sg13g2_decap_8 FILLER_172_211 ();
 sg13g2_decap_8 FILLER_172_218 ();
 sg13g2_decap_8 FILLER_172_225 ();
 sg13g2_decap_8 FILLER_172_232 ();
 sg13g2_fill_2 FILLER_172_239 ();
 sg13g2_fill_1 FILLER_172_266 ();
 sg13g2_decap_8 FILLER_172_282 ();
 sg13g2_decap_8 FILLER_172_299 ();
 sg13g2_fill_1 FILLER_172_306 ();
 sg13g2_fill_2 FILLER_172_311 ();
 sg13g2_decap_8 FILLER_172_318 ();
 sg13g2_fill_2 FILLER_172_325 ();
 sg13g2_decap_8 FILLER_172_331 ();
 sg13g2_decap_8 FILLER_172_338 ();
 sg13g2_decap_8 FILLER_172_345 ();
 sg13g2_decap_8 FILLER_172_352 ();
 sg13g2_decap_4 FILLER_172_359 ();
 sg13g2_decap_8 FILLER_172_367 ();
 sg13g2_decap_8 FILLER_172_374 ();
 sg13g2_fill_1 FILLER_172_386 ();
 sg13g2_fill_2 FILLER_172_412 ();
 sg13g2_fill_1 FILLER_172_414 ();
 sg13g2_fill_1 FILLER_172_510 ();
 sg13g2_decap_8 FILLER_172_561 ();
 sg13g2_fill_2 FILLER_172_568 ();
 sg13g2_fill_1 FILLER_172_570 ();
 sg13g2_decap_4 FILLER_172_600 ();
 sg13g2_decap_8 FILLER_172_654 ();
 sg13g2_decap_8 FILLER_172_661 ();
 sg13g2_decap_4 FILLER_172_668 ();
 sg13g2_decap_8 FILLER_172_701 ();
 sg13g2_fill_2 FILLER_172_708 ();
 sg13g2_decap_4 FILLER_172_746 ();
 sg13g2_fill_2 FILLER_172_750 ();
 sg13g2_decap_8 FILLER_172_778 ();
 sg13g2_fill_2 FILLER_172_785 ();
 sg13g2_decap_8 FILLER_172_791 ();
 sg13g2_fill_2 FILLER_172_798 ();
 sg13g2_decap_8 FILLER_172_826 ();
 sg13g2_decap_8 FILLER_172_833 ();
 sg13g2_decap_8 FILLER_172_840 ();
 sg13g2_decap_8 FILLER_172_847 ();
 sg13g2_decap_8 FILLER_172_858 ();
 sg13g2_decap_8 FILLER_172_865 ();
 sg13g2_decap_4 FILLER_172_872 ();
 sg13g2_fill_1 FILLER_172_876 ();
 sg13g2_decap_4 FILLER_172_907 ();
 sg13g2_decap_8 FILLER_172_920 ();
 sg13g2_fill_1 FILLER_172_927 ();
 sg13g2_fill_2 FILLER_172_961 ();
 sg13g2_fill_1 FILLER_172_963 ();
 sg13g2_decap_8 FILLER_172_1000 ();
 sg13g2_decap_8 FILLER_172_1007 ();
 sg13g2_decap_8 FILLER_172_1014 ();
 sg13g2_fill_2 FILLER_172_1021 ();
 sg13g2_fill_1 FILLER_172_1023 ();
 sg13g2_fill_1 FILLER_172_1032 ();
 sg13g2_decap_8 FILLER_172_1038 ();
 sg13g2_decap_4 FILLER_172_1045 ();
 sg13g2_fill_2 FILLER_172_1049 ();
 sg13g2_decap_4 FILLER_172_1055 ();
 sg13g2_decap_4 FILLER_172_1101 ();
 sg13g2_fill_1 FILLER_172_1168 ();
 sg13g2_decap_4 FILLER_172_1173 ();
 sg13g2_fill_1 FILLER_172_1177 ();
 sg13g2_fill_1 FILLER_172_1191 ();
 sg13g2_decap_8 FILLER_172_1196 ();
 sg13g2_fill_2 FILLER_172_1233 ();
 sg13g2_decap_8 FILLER_172_1261 ();
 sg13g2_decap_8 FILLER_172_1268 ();
 sg13g2_fill_2 FILLER_172_1275 ();
 sg13g2_fill_1 FILLER_172_1277 ();
 sg13g2_decap_8 FILLER_172_1282 ();
 sg13g2_fill_1 FILLER_172_1289 ();
 sg13g2_decap_8 FILLER_172_1320 ();
 sg13g2_decap_8 FILLER_172_1327 ();
 sg13g2_decap_8 FILLER_172_1334 ();
 sg13g2_decap_8 FILLER_172_1341 ();
 sg13g2_decap_8 FILLER_172_1348 ();
 sg13g2_decap_8 FILLER_172_1355 ();
 sg13g2_decap_8 FILLER_172_1362 ();
 sg13g2_decap_8 FILLER_172_1369 ();
 sg13g2_decap_8 FILLER_172_1376 ();
 sg13g2_decap_8 FILLER_172_1383 ();
 sg13g2_decap_8 FILLER_172_1390 ();
 sg13g2_decap_8 FILLER_172_1397 ();
 sg13g2_decap_8 FILLER_172_1404 ();
 sg13g2_decap_8 FILLER_172_1411 ();
 sg13g2_decap_8 FILLER_172_1418 ();
 sg13g2_decap_8 FILLER_172_1425 ();
 sg13g2_decap_8 FILLER_172_1432 ();
 sg13g2_decap_8 FILLER_172_1439 ();
 sg13g2_decap_8 FILLER_172_1446 ();
 sg13g2_decap_8 FILLER_172_1453 ();
 sg13g2_decap_8 FILLER_172_1460 ();
 sg13g2_decap_8 FILLER_172_1467 ();
 sg13g2_decap_8 FILLER_172_1474 ();
 sg13g2_decap_8 FILLER_172_1481 ();
 sg13g2_decap_8 FILLER_172_1488 ();
 sg13g2_decap_8 FILLER_172_1495 ();
 sg13g2_decap_8 FILLER_172_1502 ();
 sg13g2_decap_8 FILLER_172_1509 ();
 sg13g2_decap_8 FILLER_172_1516 ();
 sg13g2_decap_8 FILLER_172_1523 ();
 sg13g2_decap_8 FILLER_172_1530 ();
 sg13g2_decap_8 FILLER_172_1537 ();
 sg13g2_decap_8 FILLER_172_1544 ();
 sg13g2_decap_8 FILLER_172_1551 ();
 sg13g2_decap_8 FILLER_172_1558 ();
 sg13g2_decap_8 FILLER_172_1565 ();
 sg13g2_decap_8 FILLER_172_1572 ();
 sg13g2_decap_8 FILLER_172_1579 ();
 sg13g2_decap_8 FILLER_172_1586 ();
 sg13g2_decap_8 FILLER_172_1593 ();
 sg13g2_decap_8 FILLER_172_1600 ();
 sg13g2_decap_8 FILLER_172_1607 ();
 sg13g2_decap_8 FILLER_172_1614 ();
 sg13g2_decap_4 FILLER_172_1621 ();
 sg13g2_decap_8 FILLER_173_0 ();
 sg13g2_decap_8 FILLER_173_7 ();
 sg13g2_decap_8 FILLER_173_14 ();
 sg13g2_decap_8 FILLER_173_21 ();
 sg13g2_decap_8 FILLER_173_28 ();
 sg13g2_decap_8 FILLER_173_35 ();
 sg13g2_decap_8 FILLER_173_42 ();
 sg13g2_decap_8 FILLER_173_49 ();
 sg13g2_decap_8 FILLER_173_56 ();
 sg13g2_decap_8 FILLER_173_63 ();
 sg13g2_decap_8 FILLER_173_70 ();
 sg13g2_decap_8 FILLER_173_77 ();
 sg13g2_decap_8 FILLER_173_84 ();
 sg13g2_decap_8 FILLER_173_91 ();
 sg13g2_decap_8 FILLER_173_98 ();
 sg13g2_decap_8 FILLER_173_105 ();
 sg13g2_decap_8 FILLER_173_112 ();
 sg13g2_decap_8 FILLER_173_119 ();
 sg13g2_decap_8 FILLER_173_126 ();
 sg13g2_decap_8 FILLER_173_133 ();
 sg13g2_decap_8 FILLER_173_140 ();
 sg13g2_decap_8 FILLER_173_147 ();
 sg13g2_decap_8 FILLER_173_154 ();
 sg13g2_decap_8 FILLER_173_161 ();
 sg13g2_decap_8 FILLER_173_168 ();
 sg13g2_decap_8 FILLER_173_175 ();
 sg13g2_decap_4 FILLER_173_182 ();
 sg13g2_decap_8 FILLER_173_212 ();
 sg13g2_fill_2 FILLER_173_219 ();
 sg13g2_fill_1 FILLER_173_221 ();
 sg13g2_fill_2 FILLER_173_226 ();
 sg13g2_fill_1 FILLER_173_228 ();
 sg13g2_decap_8 FILLER_173_237 ();
 sg13g2_fill_2 FILLER_173_244 ();
 sg13g2_fill_1 FILLER_173_246 ();
 sg13g2_decap_4 FILLER_173_273 ();
 sg13g2_fill_1 FILLER_173_294 ();
 sg13g2_fill_2 FILLER_173_305 ();
 sg13g2_fill_1 FILLER_173_307 ();
 sg13g2_decap_8 FILLER_173_312 ();
 sg13g2_fill_1 FILLER_173_319 ();
 sg13g2_decap_8 FILLER_173_324 ();
 sg13g2_decap_8 FILLER_173_331 ();
 sg13g2_fill_2 FILLER_173_338 ();
 sg13g2_decap_8 FILLER_173_345 ();
 sg13g2_fill_2 FILLER_173_352 ();
 sg13g2_decap_8 FILLER_173_358 ();
 sg13g2_decap_4 FILLER_173_365 ();
 sg13g2_decap_8 FILLER_173_373 ();
 sg13g2_decap_4 FILLER_173_380 ();
 sg13g2_fill_1 FILLER_173_384 ();
 sg13g2_decap_8 FILLER_173_453 ();
 sg13g2_decap_4 FILLER_173_460 ();
 sg13g2_fill_2 FILLER_173_474 ();
 sg13g2_fill_1 FILLER_173_476 ();
 sg13g2_fill_2 FILLER_173_512 ();
 sg13g2_fill_2 FILLER_173_518 ();
 sg13g2_fill_1 FILLER_173_520 ();
 sg13g2_fill_1 FILLER_173_524 ();
 sg13g2_fill_1 FILLER_173_554 ();
 sg13g2_fill_2 FILLER_173_564 ();
 sg13g2_fill_2 FILLER_173_570 ();
 sg13g2_decap_4 FILLER_173_581 ();
 sg13g2_fill_1 FILLER_173_585 ();
 sg13g2_fill_1 FILLER_173_612 ();
 sg13g2_decap_8 FILLER_173_642 ();
 sg13g2_decap_4 FILLER_173_649 ();
 sg13g2_fill_2 FILLER_173_653 ();
 sg13g2_decap_8 FILLER_173_701 ();
 sg13g2_decap_8 FILLER_173_708 ();
 sg13g2_fill_2 FILLER_173_715 ();
 sg13g2_fill_1 FILLER_173_717 ();
 sg13g2_decap_8 FILLER_173_722 ();
 sg13g2_decap_4 FILLER_173_754 ();
 sg13g2_fill_2 FILLER_173_758 ();
 sg13g2_decap_8 FILLER_173_764 ();
 sg13g2_decap_8 FILLER_173_771 ();
 sg13g2_fill_1 FILLER_173_778 ();
 sg13g2_fill_2 FILLER_173_805 ();
 sg13g2_fill_1 FILLER_173_807 ();
 sg13g2_decap_8 FILLER_173_812 ();
 sg13g2_decap_8 FILLER_173_819 ();
 sg13g2_decap_8 FILLER_173_826 ();
 sg13g2_decap_8 FILLER_173_833 ();
 sg13g2_fill_2 FILLER_173_840 ();
 sg13g2_decap_8 FILLER_173_847 ();
 sg13g2_fill_2 FILLER_173_854 ();
 sg13g2_decap_8 FILLER_173_865 ();
 sg13g2_fill_1 FILLER_173_872 ();
 sg13g2_decap_8 FILLER_173_881 ();
 sg13g2_decap_8 FILLER_173_900 ();
 sg13g2_decap_8 FILLER_173_907 ();
 sg13g2_fill_2 FILLER_173_914 ();
 sg13g2_fill_1 FILLER_173_920 ();
 sg13g2_decap_8 FILLER_173_926 ();
 sg13g2_fill_1 FILLER_173_933 ();
 sg13g2_decap_8 FILLER_173_979 ();
 sg13g2_decap_8 FILLER_173_986 ();
 sg13g2_decap_8 FILLER_173_993 ();
 sg13g2_decap_4 FILLER_173_1000 ();
 sg13g2_fill_1 FILLER_173_1004 ();
 sg13g2_decap_4 FILLER_173_1009 ();
 sg13g2_fill_2 FILLER_173_1013 ();
 sg13g2_fill_1 FILLER_173_1036 ();
 sg13g2_fill_1 FILLER_173_1042 ();
 sg13g2_decap_8 FILLER_173_1069 ();
 sg13g2_decap_8 FILLER_173_1076 ();
 sg13g2_fill_2 FILLER_173_1083 ();
 sg13g2_decap_8 FILLER_173_1093 ();
 sg13g2_fill_1 FILLER_173_1105 ();
 sg13g2_decap_8 FILLER_173_1112 ();
 sg13g2_decap_8 FILLER_173_1119 ();
 sg13g2_fill_2 FILLER_173_1126 ();
 sg13g2_fill_1 FILLER_173_1128 ();
 sg13g2_fill_2 FILLER_173_1161 ();
 sg13g2_fill_1 FILLER_173_1189 ();
 sg13g2_fill_1 FILLER_173_1202 ();
 sg13g2_decap_8 FILLER_173_1209 ();
 sg13g2_decap_8 FILLER_173_1216 ();
 sg13g2_fill_2 FILLER_173_1223 ();
 sg13g2_fill_1 FILLER_173_1225 ();
 sg13g2_decap_8 FILLER_173_1230 ();
 sg13g2_decap_8 FILLER_173_1237 ();
 sg13g2_decap_4 FILLER_173_1244 ();
 sg13g2_fill_2 FILLER_173_1248 ();
 sg13g2_fill_1 FILLER_173_1264 ();
 sg13g2_decap_4 FILLER_173_1269 ();
 sg13g2_fill_2 FILLER_173_1273 ();
 sg13g2_fill_2 FILLER_173_1283 ();
 sg13g2_decap_4 FILLER_173_1293 ();
 sg13g2_fill_2 FILLER_173_1297 ();
 sg13g2_decap_8 FILLER_173_1303 ();
 sg13g2_decap_8 FILLER_173_1310 ();
 sg13g2_decap_8 FILLER_173_1317 ();
 sg13g2_decap_8 FILLER_173_1324 ();
 sg13g2_decap_8 FILLER_173_1331 ();
 sg13g2_decap_8 FILLER_173_1338 ();
 sg13g2_decap_8 FILLER_173_1345 ();
 sg13g2_decap_8 FILLER_173_1352 ();
 sg13g2_decap_8 FILLER_173_1359 ();
 sg13g2_decap_8 FILLER_173_1366 ();
 sg13g2_decap_8 FILLER_173_1373 ();
 sg13g2_decap_8 FILLER_173_1380 ();
 sg13g2_decap_8 FILLER_173_1387 ();
 sg13g2_decap_8 FILLER_173_1394 ();
 sg13g2_decap_8 FILLER_173_1401 ();
 sg13g2_decap_8 FILLER_173_1408 ();
 sg13g2_decap_8 FILLER_173_1415 ();
 sg13g2_decap_8 FILLER_173_1422 ();
 sg13g2_decap_8 FILLER_173_1429 ();
 sg13g2_decap_8 FILLER_173_1436 ();
 sg13g2_decap_8 FILLER_173_1443 ();
 sg13g2_decap_8 FILLER_173_1450 ();
 sg13g2_decap_8 FILLER_173_1457 ();
 sg13g2_decap_8 FILLER_173_1464 ();
 sg13g2_decap_8 FILLER_173_1471 ();
 sg13g2_decap_8 FILLER_173_1478 ();
 sg13g2_decap_8 FILLER_173_1485 ();
 sg13g2_decap_8 FILLER_173_1492 ();
 sg13g2_decap_8 FILLER_173_1499 ();
 sg13g2_decap_8 FILLER_173_1506 ();
 sg13g2_decap_8 FILLER_173_1513 ();
 sg13g2_decap_8 FILLER_173_1520 ();
 sg13g2_decap_8 FILLER_173_1527 ();
 sg13g2_decap_8 FILLER_173_1534 ();
 sg13g2_decap_8 FILLER_173_1541 ();
 sg13g2_decap_8 FILLER_173_1548 ();
 sg13g2_decap_8 FILLER_173_1555 ();
 sg13g2_decap_8 FILLER_173_1562 ();
 sg13g2_decap_8 FILLER_173_1569 ();
 sg13g2_decap_8 FILLER_173_1576 ();
 sg13g2_decap_8 FILLER_173_1583 ();
 sg13g2_decap_8 FILLER_173_1590 ();
 sg13g2_decap_8 FILLER_173_1597 ();
 sg13g2_decap_8 FILLER_173_1604 ();
 sg13g2_decap_8 FILLER_173_1611 ();
 sg13g2_decap_8 FILLER_173_1618 ();
 sg13g2_decap_8 FILLER_174_0 ();
 sg13g2_decap_8 FILLER_174_7 ();
 sg13g2_decap_8 FILLER_174_14 ();
 sg13g2_decap_8 FILLER_174_21 ();
 sg13g2_decap_8 FILLER_174_28 ();
 sg13g2_decap_8 FILLER_174_35 ();
 sg13g2_decap_8 FILLER_174_42 ();
 sg13g2_decap_8 FILLER_174_49 ();
 sg13g2_decap_8 FILLER_174_56 ();
 sg13g2_decap_8 FILLER_174_63 ();
 sg13g2_decap_8 FILLER_174_70 ();
 sg13g2_decap_8 FILLER_174_77 ();
 sg13g2_decap_8 FILLER_174_84 ();
 sg13g2_decap_8 FILLER_174_91 ();
 sg13g2_decap_8 FILLER_174_98 ();
 sg13g2_decap_8 FILLER_174_105 ();
 sg13g2_decap_8 FILLER_174_112 ();
 sg13g2_decap_8 FILLER_174_119 ();
 sg13g2_decap_8 FILLER_174_126 ();
 sg13g2_decap_8 FILLER_174_133 ();
 sg13g2_decap_8 FILLER_174_140 ();
 sg13g2_decap_8 FILLER_174_147 ();
 sg13g2_decap_8 FILLER_174_154 ();
 sg13g2_decap_8 FILLER_174_161 ();
 sg13g2_decap_8 FILLER_174_168 ();
 sg13g2_decap_8 FILLER_174_175 ();
 sg13g2_decap_8 FILLER_174_182 ();
 sg13g2_decap_8 FILLER_174_189 ();
 sg13g2_decap_8 FILLER_174_196 ();
 sg13g2_fill_2 FILLER_174_203 ();
 sg13g2_fill_2 FILLER_174_208 ();
 sg13g2_fill_1 FILLER_174_210 ();
 sg13g2_decap_4 FILLER_174_241 ();
 sg13g2_fill_2 FILLER_174_245 ();
 sg13g2_fill_2 FILLER_174_251 ();
 sg13g2_fill_2 FILLER_174_279 ();
 sg13g2_fill_1 FILLER_174_281 ();
 sg13g2_fill_1 FILLER_174_286 ();
 sg13g2_decap_4 FILLER_174_292 ();
 sg13g2_fill_2 FILLER_174_301 ();
 sg13g2_fill_1 FILLER_174_303 ();
 sg13g2_fill_2 FILLER_174_310 ();
 sg13g2_decap_8 FILLER_174_343 ();
 sg13g2_fill_1 FILLER_174_350 ();
 sg13g2_decap_8 FILLER_174_386 ();
 sg13g2_fill_2 FILLER_174_419 ();
 sg13g2_decap_8 FILLER_174_456 ();
 sg13g2_fill_1 FILLER_174_463 ();
 sg13g2_fill_2 FILLER_174_499 ();
 sg13g2_fill_1 FILLER_174_501 ();
 sg13g2_fill_1 FILLER_174_506 ();
 sg13g2_decap_4 FILLER_174_597 ();
 sg13g2_fill_1 FILLER_174_601 ();
 sg13g2_fill_2 FILLER_174_606 ();
 sg13g2_fill_1 FILLER_174_608 ();
 sg13g2_decap_4 FILLER_174_638 ();
 sg13g2_fill_1 FILLER_174_642 ();
 sg13g2_decap_8 FILLER_174_669 ();
 sg13g2_decap_8 FILLER_174_683 ();
 sg13g2_decap_8 FILLER_174_690 ();
 sg13g2_decap_8 FILLER_174_697 ();
 sg13g2_decap_8 FILLER_174_704 ();
 sg13g2_decap_8 FILLER_174_711 ();
 sg13g2_decap_4 FILLER_174_761 ();
 sg13g2_fill_1 FILLER_174_765 ();
 sg13g2_decap_8 FILLER_174_802 ();
 sg13g2_decap_8 FILLER_174_809 ();
 sg13g2_decap_8 FILLER_174_816 ();
 sg13g2_decap_8 FILLER_174_827 ();
 sg13g2_decap_8 FILLER_174_834 ();
 sg13g2_decap_8 FILLER_174_841 ();
 sg13g2_decap_4 FILLER_174_848 ();
 sg13g2_fill_1 FILLER_174_852 ();
 sg13g2_decap_8 FILLER_174_883 ();
 sg13g2_decap_8 FILLER_174_890 ();
 sg13g2_fill_2 FILLER_174_897 ();
 sg13g2_fill_1 FILLER_174_899 ();
 sg13g2_fill_2 FILLER_174_907 ();
 sg13g2_fill_1 FILLER_174_909 ();
 sg13g2_decap_8 FILLER_174_930 ();
 sg13g2_decap_8 FILLER_174_937 ();
 sg13g2_decap_4 FILLER_174_944 ();
 sg13g2_fill_1 FILLER_174_948 ();
 sg13g2_fill_2 FILLER_174_953 ();
 sg13g2_decap_8 FILLER_174_967 ();
 sg13g2_decap_8 FILLER_174_974 ();
 sg13g2_decap_4 FILLER_174_981 ();
 sg13g2_fill_1 FILLER_174_985 ();
 sg13g2_decap_8 FILLER_174_990 ();
 sg13g2_fill_2 FILLER_174_997 ();
 sg13g2_decap_8 FILLER_174_1025 ();
 sg13g2_fill_2 FILLER_174_1032 ();
 sg13g2_fill_1 FILLER_174_1034 ();
 sg13g2_decap_8 FILLER_174_1039 ();
 sg13g2_decap_4 FILLER_174_1046 ();
 sg13g2_fill_2 FILLER_174_1054 ();
 sg13g2_decap_8 FILLER_174_1060 ();
 sg13g2_decap_4 FILLER_174_1067 ();
 sg13g2_fill_2 FILLER_174_1103 ();
 sg13g2_decap_8 FILLER_174_1115 ();
 sg13g2_fill_1 FILLER_174_1122 ();
 sg13g2_decap_8 FILLER_174_1153 ();
 sg13g2_decap_8 FILLER_174_1160 ();
 sg13g2_decap_8 FILLER_174_1167 ();
 sg13g2_decap_8 FILLER_174_1185 ();
 sg13g2_decap_8 FILLER_174_1192 ();
 sg13g2_decap_4 FILLER_174_1199 ();
 sg13g2_fill_2 FILLER_174_1203 ();
 sg13g2_decap_4 FILLER_174_1219 ();
 sg13g2_decap_8 FILLER_174_1227 ();
 sg13g2_decap_8 FILLER_174_1234 ();
 sg13g2_fill_1 FILLER_174_1241 ();
 sg13g2_decap_8 FILLER_174_1247 ();
 sg13g2_fill_2 FILLER_174_1254 ();
 sg13g2_decap_4 FILLER_174_1266 ();
 sg13g2_decap_4 FILLER_174_1276 ();
 sg13g2_fill_2 FILLER_174_1280 ();
 sg13g2_decap_8 FILLER_174_1290 ();
 sg13g2_decap_4 FILLER_174_1297 ();
 sg13g2_fill_2 FILLER_174_1301 ();
 sg13g2_decap_8 FILLER_174_1307 ();
 sg13g2_decap_8 FILLER_174_1314 ();
 sg13g2_decap_8 FILLER_174_1321 ();
 sg13g2_decap_8 FILLER_174_1328 ();
 sg13g2_decap_8 FILLER_174_1335 ();
 sg13g2_decap_8 FILLER_174_1342 ();
 sg13g2_decap_8 FILLER_174_1349 ();
 sg13g2_decap_8 FILLER_174_1356 ();
 sg13g2_decap_8 FILLER_174_1363 ();
 sg13g2_decap_8 FILLER_174_1370 ();
 sg13g2_decap_8 FILLER_174_1377 ();
 sg13g2_decap_8 FILLER_174_1384 ();
 sg13g2_decap_8 FILLER_174_1391 ();
 sg13g2_decap_8 FILLER_174_1398 ();
 sg13g2_decap_8 FILLER_174_1405 ();
 sg13g2_decap_8 FILLER_174_1412 ();
 sg13g2_decap_8 FILLER_174_1419 ();
 sg13g2_decap_8 FILLER_174_1426 ();
 sg13g2_decap_8 FILLER_174_1433 ();
 sg13g2_decap_8 FILLER_174_1440 ();
 sg13g2_decap_8 FILLER_174_1447 ();
 sg13g2_decap_8 FILLER_174_1454 ();
 sg13g2_decap_8 FILLER_174_1461 ();
 sg13g2_decap_8 FILLER_174_1468 ();
 sg13g2_decap_8 FILLER_174_1475 ();
 sg13g2_decap_8 FILLER_174_1482 ();
 sg13g2_decap_8 FILLER_174_1489 ();
 sg13g2_decap_8 FILLER_174_1496 ();
 sg13g2_decap_8 FILLER_174_1503 ();
 sg13g2_decap_8 FILLER_174_1510 ();
 sg13g2_decap_8 FILLER_174_1517 ();
 sg13g2_decap_8 FILLER_174_1524 ();
 sg13g2_decap_8 FILLER_174_1531 ();
 sg13g2_decap_8 FILLER_174_1538 ();
 sg13g2_decap_8 FILLER_174_1545 ();
 sg13g2_decap_8 FILLER_174_1552 ();
 sg13g2_decap_8 FILLER_174_1559 ();
 sg13g2_decap_8 FILLER_174_1566 ();
 sg13g2_decap_8 FILLER_174_1573 ();
 sg13g2_decap_8 FILLER_174_1580 ();
 sg13g2_decap_8 FILLER_174_1587 ();
 sg13g2_decap_8 FILLER_174_1594 ();
 sg13g2_decap_8 FILLER_174_1601 ();
 sg13g2_decap_8 FILLER_174_1608 ();
 sg13g2_decap_8 FILLER_174_1615 ();
 sg13g2_fill_2 FILLER_174_1622 ();
 sg13g2_fill_1 FILLER_174_1624 ();
 sg13g2_decap_8 FILLER_175_0 ();
 sg13g2_decap_8 FILLER_175_7 ();
 sg13g2_decap_8 FILLER_175_14 ();
 sg13g2_decap_8 FILLER_175_21 ();
 sg13g2_decap_8 FILLER_175_28 ();
 sg13g2_decap_8 FILLER_175_35 ();
 sg13g2_decap_8 FILLER_175_42 ();
 sg13g2_decap_8 FILLER_175_49 ();
 sg13g2_decap_8 FILLER_175_56 ();
 sg13g2_decap_8 FILLER_175_63 ();
 sg13g2_decap_8 FILLER_175_70 ();
 sg13g2_decap_8 FILLER_175_77 ();
 sg13g2_decap_8 FILLER_175_84 ();
 sg13g2_decap_8 FILLER_175_91 ();
 sg13g2_decap_8 FILLER_175_98 ();
 sg13g2_decap_8 FILLER_175_105 ();
 sg13g2_decap_8 FILLER_175_112 ();
 sg13g2_decap_8 FILLER_175_119 ();
 sg13g2_decap_8 FILLER_175_126 ();
 sg13g2_decap_8 FILLER_175_133 ();
 sg13g2_decap_8 FILLER_175_140 ();
 sg13g2_decap_8 FILLER_175_147 ();
 sg13g2_decap_8 FILLER_175_154 ();
 sg13g2_decap_8 FILLER_175_161 ();
 sg13g2_decap_8 FILLER_175_168 ();
 sg13g2_decap_8 FILLER_175_175 ();
 sg13g2_decap_8 FILLER_175_182 ();
 sg13g2_decap_8 FILLER_175_189 ();
 sg13g2_decap_8 FILLER_175_196 ();
 sg13g2_fill_2 FILLER_175_203 ();
 sg13g2_decap_4 FILLER_175_230 ();
 sg13g2_fill_2 FILLER_175_234 ();
 sg13g2_decap_8 FILLER_175_241 ();
 sg13g2_decap_8 FILLER_175_248 ();
 sg13g2_fill_2 FILLER_175_286 ();
 sg13g2_fill_2 FILLER_175_293 ();
 sg13g2_decap_4 FILLER_175_320 ();
 sg13g2_decap_8 FILLER_175_329 ();
 sg13g2_fill_2 FILLER_175_348 ();
 sg13g2_fill_1 FILLER_175_350 ();
 sg13g2_fill_2 FILLER_175_356 ();
 sg13g2_fill_1 FILLER_175_358 ();
 sg13g2_decap_8 FILLER_175_369 ();
 sg13g2_decap_4 FILLER_175_376 ();
 sg13g2_fill_2 FILLER_175_380 ();
 sg13g2_fill_2 FILLER_175_391 ();
 sg13g2_fill_1 FILLER_175_406 ();
 sg13g2_decap_4 FILLER_175_425 ();
 sg13g2_fill_2 FILLER_175_429 ();
 sg13g2_decap_8 FILLER_175_460 ();
 sg13g2_decap_4 FILLER_175_467 ();
 sg13g2_fill_1 FILLER_175_471 ();
 sg13g2_decap_8 FILLER_175_477 ();
 sg13g2_decap_8 FILLER_175_484 ();
 sg13g2_decap_8 FILLER_175_491 ();
 sg13g2_fill_1 FILLER_175_498 ();
 sg13g2_fill_1 FILLER_175_507 ();
 sg13g2_fill_2 FILLER_175_639 ();
 sg13g2_fill_1 FILLER_175_641 ();
 sg13g2_decap_4 FILLER_175_667 ();
 sg13g2_fill_1 FILLER_175_697 ();
 sg13g2_fill_1 FILLER_175_742 ();
 sg13g2_fill_2 FILLER_175_779 ();
 sg13g2_fill_1 FILLER_175_781 ();
 sg13g2_fill_2 FILLER_175_811 ();
 sg13g2_fill_1 FILLER_175_813 ();
 sg13g2_decap_8 FILLER_175_848 ();
 sg13g2_decap_4 FILLER_175_855 ();
 sg13g2_fill_2 FILLER_175_863 ();
 sg13g2_fill_1 FILLER_175_894 ();
 sg13g2_fill_2 FILLER_175_903 ();
 sg13g2_fill_1 FILLER_175_905 ();
 sg13g2_fill_2 FILLER_175_1005 ();
 sg13g2_fill_1 FILLER_175_1007 ();
 sg13g2_fill_1 FILLER_175_1034 ();
 sg13g2_fill_2 FILLER_175_1074 ();
 sg13g2_fill_2 FILLER_175_1102 ();
 sg13g2_fill_1 FILLER_175_1104 ();
 sg13g2_fill_2 FILLER_175_1113 ();
 sg13g2_fill_1 FILLER_175_1115 ();
 sg13g2_decap_8 FILLER_175_1120 ();
 sg13g2_decap_8 FILLER_175_1127 ();
 sg13g2_decap_8 FILLER_175_1138 ();
 sg13g2_decap_8 FILLER_175_1145 ();
 sg13g2_decap_4 FILLER_175_1152 ();
 sg13g2_fill_2 FILLER_175_1199 ();
 sg13g2_fill_2 FILLER_175_1213 ();
 sg13g2_fill_2 FILLER_175_1241 ();
 sg13g2_fill_1 FILLER_175_1243 ();
 sg13g2_fill_1 FILLER_175_1252 ();
 sg13g2_decap_8 FILLER_175_1258 ();
 sg13g2_fill_1 FILLER_175_1265 ();
 sg13g2_fill_2 FILLER_175_1274 ();
 sg13g2_fill_1 FILLER_175_1276 ();
 sg13g2_decap_4 FILLER_175_1281 ();
 sg13g2_fill_2 FILLER_175_1285 ();
 sg13g2_decap_4 FILLER_175_1291 ();
 sg13g2_decap_8 FILLER_175_1321 ();
 sg13g2_decap_8 FILLER_175_1328 ();
 sg13g2_decap_8 FILLER_175_1335 ();
 sg13g2_decap_8 FILLER_175_1342 ();
 sg13g2_decap_8 FILLER_175_1349 ();
 sg13g2_decap_8 FILLER_175_1356 ();
 sg13g2_decap_8 FILLER_175_1363 ();
 sg13g2_decap_8 FILLER_175_1370 ();
 sg13g2_decap_8 FILLER_175_1377 ();
 sg13g2_decap_8 FILLER_175_1384 ();
 sg13g2_decap_8 FILLER_175_1391 ();
 sg13g2_decap_8 FILLER_175_1398 ();
 sg13g2_decap_8 FILLER_175_1405 ();
 sg13g2_decap_8 FILLER_175_1412 ();
 sg13g2_decap_8 FILLER_175_1419 ();
 sg13g2_decap_8 FILLER_175_1426 ();
 sg13g2_decap_8 FILLER_175_1433 ();
 sg13g2_decap_8 FILLER_175_1440 ();
 sg13g2_decap_8 FILLER_175_1447 ();
 sg13g2_decap_8 FILLER_175_1454 ();
 sg13g2_decap_8 FILLER_175_1461 ();
 sg13g2_decap_8 FILLER_175_1468 ();
 sg13g2_decap_8 FILLER_175_1475 ();
 sg13g2_decap_8 FILLER_175_1482 ();
 sg13g2_decap_8 FILLER_175_1489 ();
 sg13g2_decap_8 FILLER_175_1496 ();
 sg13g2_decap_8 FILLER_175_1503 ();
 sg13g2_decap_8 FILLER_175_1510 ();
 sg13g2_decap_8 FILLER_175_1517 ();
 sg13g2_decap_8 FILLER_175_1524 ();
 sg13g2_decap_8 FILLER_175_1531 ();
 sg13g2_decap_8 FILLER_175_1538 ();
 sg13g2_decap_8 FILLER_175_1545 ();
 sg13g2_decap_8 FILLER_175_1552 ();
 sg13g2_decap_8 FILLER_175_1559 ();
 sg13g2_decap_8 FILLER_175_1566 ();
 sg13g2_decap_8 FILLER_175_1573 ();
 sg13g2_decap_8 FILLER_175_1580 ();
 sg13g2_decap_8 FILLER_175_1587 ();
 sg13g2_decap_8 FILLER_175_1594 ();
 sg13g2_decap_8 FILLER_175_1601 ();
 sg13g2_decap_8 FILLER_175_1608 ();
 sg13g2_decap_8 FILLER_175_1615 ();
 sg13g2_fill_2 FILLER_175_1622 ();
 sg13g2_fill_1 FILLER_175_1624 ();
 sg13g2_decap_8 FILLER_176_0 ();
 sg13g2_decap_8 FILLER_176_7 ();
 sg13g2_decap_8 FILLER_176_14 ();
 sg13g2_decap_8 FILLER_176_21 ();
 sg13g2_decap_8 FILLER_176_28 ();
 sg13g2_decap_8 FILLER_176_35 ();
 sg13g2_decap_8 FILLER_176_42 ();
 sg13g2_decap_8 FILLER_176_49 ();
 sg13g2_decap_8 FILLER_176_56 ();
 sg13g2_decap_8 FILLER_176_63 ();
 sg13g2_decap_8 FILLER_176_70 ();
 sg13g2_decap_8 FILLER_176_77 ();
 sg13g2_decap_8 FILLER_176_84 ();
 sg13g2_decap_8 FILLER_176_91 ();
 sg13g2_decap_8 FILLER_176_98 ();
 sg13g2_decap_8 FILLER_176_105 ();
 sg13g2_decap_8 FILLER_176_112 ();
 sg13g2_decap_8 FILLER_176_119 ();
 sg13g2_decap_8 FILLER_176_126 ();
 sg13g2_decap_8 FILLER_176_133 ();
 sg13g2_decap_8 FILLER_176_140 ();
 sg13g2_decap_8 FILLER_176_147 ();
 sg13g2_decap_8 FILLER_176_154 ();
 sg13g2_decap_8 FILLER_176_161 ();
 sg13g2_decap_8 FILLER_176_168 ();
 sg13g2_decap_8 FILLER_176_175 ();
 sg13g2_decap_8 FILLER_176_182 ();
 sg13g2_decap_8 FILLER_176_189 ();
 sg13g2_decap_8 FILLER_176_196 ();
 sg13g2_decap_8 FILLER_176_203 ();
 sg13g2_decap_8 FILLER_176_210 ();
 sg13g2_decap_8 FILLER_176_217 ();
 sg13g2_decap_8 FILLER_176_224 ();
 sg13g2_decap_8 FILLER_176_231 ();
 sg13g2_decap_8 FILLER_176_250 ();
 sg13g2_fill_1 FILLER_176_257 ();
 sg13g2_decap_8 FILLER_176_296 ();
 sg13g2_decap_8 FILLER_176_303 ();
 sg13g2_decap_8 FILLER_176_319 ();
 sg13g2_decap_4 FILLER_176_326 ();
 sg13g2_decap_4 FILLER_176_334 ();
 sg13g2_fill_1 FILLER_176_338 ();
 sg13g2_decap_4 FILLER_176_344 ();
 sg13g2_decap_4 FILLER_176_381 ();
 sg13g2_fill_1 FILLER_176_385 ();
 sg13g2_decap_8 FILLER_176_394 ();
 sg13g2_decap_8 FILLER_176_401 ();
 sg13g2_fill_1 FILLER_176_408 ();
 sg13g2_fill_1 FILLER_176_434 ();
 sg13g2_fill_2 FILLER_176_456 ();
 sg13g2_decap_8 FILLER_176_463 ();
 sg13g2_decap_8 FILLER_176_470 ();
 sg13g2_decap_4 FILLER_176_477 ();
 sg13g2_fill_2 FILLER_176_481 ();
 sg13g2_decap_4 FILLER_176_492 ();
 sg13g2_fill_1 FILLER_176_496 ();
 sg13g2_fill_1 FILLER_176_502 ();
 sg13g2_fill_1 FILLER_176_543 ();
 sg13g2_fill_2 FILLER_176_573 ();
 sg13g2_fill_1 FILLER_176_630 ();
 sg13g2_decap_4 FILLER_176_671 ();
 sg13g2_fill_2 FILLER_176_675 ();
 sg13g2_fill_2 FILLER_176_712 ();
 sg13g2_fill_1 FILLER_176_714 ();
 sg13g2_fill_2 FILLER_176_775 ();
 sg13g2_fill_1 FILLER_176_777 ();
 sg13g2_decap_8 FILLER_176_804 ();
 sg13g2_decap_8 FILLER_176_811 ();
 sg13g2_decap_8 FILLER_176_818 ();
 sg13g2_decap_4 FILLER_176_825 ();
 sg13g2_fill_1 FILLER_176_829 ();
 sg13g2_fill_2 FILLER_176_902 ();
 sg13g2_fill_1 FILLER_176_921 ();
 sg13g2_decap_8 FILLER_176_926 ();
 sg13g2_fill_1 FILLER_176_933 ();
 sg13g2_decap_4 FILLER_176_959 ();
 sg13g2_decap_8 FILLER_176_967 ();
 sg13g2_decap_8 FILLER_176_974 ();
 sg13g2_decap_8 FILLER_176_981 ();
 sg13g2_fill_1 FILLER_176_988 ();
 sg13g2_decap_4 FILLER_176_1023 ();
 sg13g2_fill_1 FILLER_176_1027 ();
 sg13g2_fill_2 FILLER_176_1045 ();
 sg13g2_fill_1 FILLER_176_1047 ();
 sg13g2_decap_8 FILLER_176_1074 ();
 sg13g2_fill_2 FILLER_176_1081 ();
 sg13g2_decap_8 FILLER_176_1087 ();
 sg13g2_fill_2 FILLER_176_1094 ();
 sg13g2_fill_2 FILLER_176_1101 ();
 sg13g2_decap_8 FILLER_176_1133 ();
 sg13g2_decap_8 FILLER_176_1140 ();
 sg13g2_fill_2 FILLER_176_1147 ();
 sg13g2_fill_2 FILLER_176_1179 ();
 sg13g2_fill_1 FILLER_176_1189 ();
 sg13g2_decap_8 FILLER_176_1195 ();
 sg13g2_decap_8 FILLER_176_1202 ();
 sg13g2_decap_4 FILLER_176_1209 ();
 sg13g2_fill_1 FILLER_176_1213 ();
 sg13g2_decap_8 FILLER_176_1218 ();
 sg13g2_decap_8 FILLER_176_1225 ();
 sg13g2_fill_1 FILLER_176_1265 ();
 sg13g2_decap_8 FILLER_176_1299 ();
 sg13g2_decap_8 FILLER_176_1306 ();
 sg13g2_decap_8 FILLER_176_1313 ();
 sg13g2_decap_8 FILLER_176_1320 ();
 sg13g2_decap_8 FILLER_176_1327 ();
 sg13g2_decap_8 FILLER_176_1334 ();
 sg13g2_decap_8 FILLER_176_1341 ();
 sg13g2_decap_8 FILLER_176_1348 ();
 sg13g2_decap_8 FILLER_176_1355 ();
 sg13g2_decap_8 FILLER_176_1362 ();
 sg13g2_decap_8 FILLER_176_1369 ();
 sg13g2_decap_8 FILLER_176_1376 ();
 sg13g2_decap_8 FILLER_176_1383 ();
 sg13g2_decap_8 FILLER_176_1390 ();
 sg13g2_decap_8 FILLER_176_1397 ();
 sg13g2_decap_8 FILLER_176_1404 ();
 sg13g2_decap_8 FILLER_176_1411 ();
 sg13g2_decap_8 FILLER_176_1418 ();
 sg13g2_decap_8 FILLER_176_1425 ();
 sg13g2_decap_8 FILLER_176_1432 ();
 sg13g2_decap_8 FILLER_176_1439 ();
 sg13g2_decap_8 FILLER_176_1446 ();
 sg13g2_decap_8 FILLER_176_1453 ();
 sg13g2_decap_8 FILLER_176_1460 ();
 sg13g2_decap_8 FILLER_176_1467 ();
 sg13g2_decap_8 FILLER_176_1474 ();
 sg13g2_decap_8 FILLER_176_1481 ();
 sg13g2_decap_8 FILLER_176_1488 ();
 sg13g2_decap_8 FILLER_176_1495 ();
 sg13g2_decap_8 FILLER_176_1502 ();
 sg13g2_decap_8 FILLER_176_1509 ();
 sg13g2_decap_8 FILLER_176_1516 ();
 sg13g2_decap_8 FILLER_176_1523 ();
 sg13g2_decap_8 FILLER_176_1530 ();
 sg13g2_decap_8 FILLER_176_1537 ();
 sg13g2_decap_8 FILLER_176_1544 ();
 sg13g2_decap_8 FILLER_176_1551 ();
 sg13g2_decap_8 FILLER_176_1558 ();
 sg13g2_decap_8 FILLER_176_1565 ();
 sg13g2_decap_8 FILLER_176_1572 ();
 sg13g2_decap_8 FILLER_176_1579 ();
 sg13g2_decap_8 FILLER_176_1586 ();
 sg13g2_decap_8 FILLER_176_1593 ();
 sg13g2_decap_8 FILLER_176_1600 ();
 sg13g2_decap_8 FILLER_176_1607 ();
 sg13g2_decap_8 FILLER_176_1614 ();
 sg13g2_decap_4 FILLER_176_1621 ();
 sg13g2_decap_8 FILLER_177_0 ();
 sg13g2_decap_8 FILLER_177_7 ();
 sg13g2_decap_8 FILLER_177_14 ();
 sg13g2_decap_8 FILLER_177_21 ();
 sg13g2_decap_8 FILLER_177_28 ();
 sg13g2_decap_8 FILLER_177_35 ();
 sg13g2_decap_8 FILLER_177_42 ();
 sg13g2_decap_8 FILLER_177_49 ();
 sg13g2_decap_8 FILLER_177_56 ();
 sg13g2_decap_8 FILLER_177_63 ();
 sg13g2_decap_8 FILLER_177_70 ();
 sg13g2_decap_8 FILLER_177_77 ();
 sg13g2_decap_8 FILLER_177_84 ();
 sg13g2_decap_8 FILLER_177_91 ();
 sg13g2_decap_8 FILLER_177_98 ();
 sg13g2_decap_8 FILLER_177_105 ();
 sg13g2_decap_8 FILLER_177_112 ();
 sg13g2_decap_8 FILLER_177_119 ();
 sg13g2_decap_8 FILLER_177_126 ();
 sg13g2_decap_8 FILLER_177_133 ();
 sg13g2_decap_8 FILLER_177_140 ();
 sg13g2_decap_8 FILLER_177_147 ();
 sg13g2_decap_8 FILLER_177_154 ();
 sg13g2_decap_8 FILLER_177_161 ();
 sg13g2_decap_8 FILLER_177_168 ();
 sg13g2_decap_8 FILLER_177_175 ();
 sg13g2_decap_8 FILLER_177_182 ();
 sg13g2_decap_8 FILLER_177_189 ();
 sg13g2_decap_8 FILLER_177_196 ();
 sg13g2_decap_8 FILLER_177_203 ();
 sg13g2_fill_2 FILLER_177_210 ();
 sg13g2_fill_1 FILLER_177_212 ();
 sg13g2_decap_4 FILLER_177_221 ();
 sg13g2_fill_1 FILLER_177_225 ();
 sg13g2_decap_4 FILLER_177_238 ();
 sg13g2_decap_8 FILLER_177_247 ();
 sg13g2_decap_8 FILLER_177_254 ();
 sg13g2_decap_8 FILLER_177_261 ();
 sg13g2_decap_8 FILLER_177_268 ();
 sg13g2_fill_2 FILLER_177_285 ();
 sg13g2_fill_1 FILLER_177_287 ();
 sg13g2_decap_8 FILLER_177_292 ();
 sg13g2_decap_4 FILLER_177_299 ();
 sg13g2_fill_2 FILLER_177_303 ();
 sg13g2_decap_8 FILLER_177_318 ();
 sg13g2_fill_2 FILLER_177_341 ();
 sg13g2_fill_2 FILLER_177_369 ();
 sg13g2_decap_8 FILLER_177_380 ();
 sg13g2_decap_8 FILLER_177_391 ();
 sg13g2_decap_4 FILLER_177_398 ();
 sg13g2_fill_1 FILLER_177_402 ();
 sg13g2_fill_2 FILLER_177_407 ();
 sg13g2_fill_2 FILLER_177_418 ();
 sg13g2_decap_8 FILLER_177_424 ();
 sg13g2_decap_4 FILLER_177_431 ();
 sg13g2_fill_2 FILLER_177_435 ();
 sg13g2_fill_2 FILLER_177_463 ();
 sg13g2_fill_2 FILLER_177_469 ();
 sg13g2_fill_2 FILLER_177_476 ();
 sg13g2_fill_1 FILLER_177_478 ();
 sg13g2_fill_2 FILLER_177_483 ();
 sg13g2_fill_1 FILLER_177_485 ();
 sg13g2_fill_2 FILLER_177_491 ();
 sg13g2_decap_8 FILLER_177_497 ();
 sg13g2_decap_8 FILLER_177_504 ();
 sg13g2_fill_2 FILLER_177_511 ();
 sg13g2_fill_1 FILLER_177_513 ();
 sg13g2_decap_8 FILLER_177_518 ();
 sg13g2_fill_1 FILLER_177_525 ();
 sg13g2_fill_1 FILLER_177_539 ();
 sg13g2_fill_2 FILLER_177_571 ();
 sg13g2_fill_2 FILLER_177_603 ();
 sg13g2_fill_1 FILLER_177_605 ();
 sg13g2_fill_1 FILLER_177_611 ();
 sg13g2_decap_8 FILLER_177_616 ();
 sg13g2_decap_8 FILLER_177_623 ();
 sg13g2_decap_4 FILLER_177_634 ();
 sg13g2_decap_8 FILLER_177_642 ();
 sg13g2_fill_1 FILLER_177_649 ();
 sg13g2_decap_8 FILLER_177_654 ();
 sg13g2_fill_2 FILLER_177_661 ();
 sg13g2_fill_1 FILLER_177_663 ();
 sg13g2_decap_8 FILLER_177_668 ();
 sg13g2_decap_8 FILLER_177_675 ();
 sg13g2_fill_1 FILLER_177_682 ();
 sg13g2_fill_2 FILLER_177_691 ();
 sg13g2_fill_2 FILLER_177_719 ();
 sg13g2_fill_1 FILLER_177_721 ();
 sg13g2_fill_2 FILLER_177_774 ();
 sg13g2_fill_1 FILLER_177_776 ();
 sg13g2_decap_8 FILLER_177_816 ();
 sg13g2_decap_8 FILLER_177_823 ();
 sg13g2_fill_1 FILLER_177_830 ();
 sg13g2_fill_2 FILLER_177_834 ();
 sg13g2_fill_1 FILLER_177_841 ();
 sg13g2_fill_2 FILLER_177_847 ();
 sg13g2_decap_8 FILLER_177_854 ();
 sg13g2_decap_8 FILLER_177_861 ();
 sg13g2_decap_8 FILLER_177_868 ();
 sg13g2_decap_8 FILLER_177_875 ();
 sg13g2_decap_8 FILLER_177_882 ();
 sg13g2_decap_8 FILLER_177_889 ();
 sg13g2_decap_4 FILLER_177_896 ();
 sg13g2_decap_4 FILLER_177_912 ();
 sg13g2_fill_2 FILLER_177_987 ();
 sg13g2_fill_1 FILLER_177_989 ();
 sg13g2_decap_8 FILLER_177_1012 ();
 sg13g2_decap_8 FILLER_177_1025 ();
 sg13g2_decap_8 FILLER_177_1032 ();
 sg13g2_decap_8 FILLER_177_1039 ();
 sg13g2_decap_4 FILLER_177_1046 ();
 sg13g2_decap_8 FILLER_177_1054 ();
 sg13g2_fill_1 FILLER_177_1061 ();
 sg13g2_decap_4 FILLER_177_1072 ();
 sg13g2_decap_4 FILLER_177_1080 ();
 sg13g2_fill_2 FILLER_177_1109 ();
 sg13g2_decap_8 FILLER_177_1117 ();
 sg13g2_fill_2 FILLER_177_1124 ();
 sg13g2_fill_2 FILLER_177_1142 ();
 sg13g2_decap_8 FILLER_177_1153 ();
 sg13g2_decap_8 FILLER_177_1160 ();
 sg13g2_fill_2 FILLER_177_1167 ();
 sg13g2_decap_8 FILLER_177_1215 ();
 sg13g2_decap_8 FILLER_177_1222 ();
 sg13g2_fill_2 FILLER_177_1229 ();
 sg13g2_fill_1 FILLER_177_1231 ();
 sg13g2_decap_8 FILLER_177_1261 ();
 sg13g2_decap_8 FILLER_177_1268 ();
 sg13g2_decap_8 FILLER_177_1275 ();
 sg13g2_decap_4 FILLER_177_1282 ();
 sg13g2_fill_1 FILLER_177_1286 ();
 sg13g2_decap_8 FILLER_177_1312 ();
 sg13g2_decap_8 FILLER_177_1319 ();
 sg13g2_decap_8 FILLER_177_1326 ();
 sg13g2_decap_8 FILLER_177_1333 ();
 sg13g2_decap_8 FILLER_177_1340 ();
 sg13g2_decap_8 FILLER_177_1347 ();
 sg13g2_decap_8 FILLER_177_1354 ();
 sg13g2_decap_8 FILLER_177_1361 ();
 sg13g2_decap_8 FILLER_177_1368 ();
 sg13g2_decap_8 FILLER_177_1375 ();
 sg13g2_decap_8 FILLER_177_1382 ();
 sg13g2_decap_8 FILLER_177_1389 ();
 sg13g2_decap_8 FILLER_177_1396 ();
 sg13g2_decap_8 FILLER_177_1403 ();
 sg13g2_decap_8 FILLER_177_1410 ();
 sg13g2_decap_8 FILLER_177_1417 ();
 sg13g2_decap_8 FILLER_177_1424 ();
 sg13g2_decap_8 FILLER_177_1431 ();
 sg13g2_decap_8 FILLER_177_1438 ();
 sg13g2_decap_8 FILLER_177_1445 ();
 sg13g2_decap_8 FILLER_177_1452 ();
 sg13g2_decap_8 FILLER_177_1459 ();
 sg13g2_decap_8 FILLER_177_1466 ();
 sg13g2_decap_8 FILLER_177_1473 ();
 sg13g2_decap_8 FILLER_177_1480 ();
 sg13g2_decap_8 FILLER_177_1487 ();
 sg13g2_decap_8 FILLER_177_1494 ();
 sg13g2_decap_8 FILLER_177_1501 ();
 sg13g2_decap_8 FILLER_177_1508 ();
 sg13g2_decap_8 FILLER_177_1515 ();
 sg13g2_decap_8 FILLER_177_1522 ();
 sg13g2_decap_8 FILLER_177_1529 ();
 sg13g2_decap_8 FILLER_177_1536 ();
 sg13g2_decap_8 FILLER_177_1543 ();
 sg13g2_decap_8 FILLER_177_1550 ();
 sg13g2_decap_8 FILLER_177_1557 ();
 sg13g2_decap_8 FILLER_177_1564 ();
 sg13g2_decap_8 FILLER_177_1571 ();
 sg13g2_decap_8 FILLER_177_1578 ();
 sg13g2_decap_8 FILLER_177_1585 ();
 sg13g2_decap_8 FILLER_177_1592 ();
 sg13g2_decap_8 FILLER_177_1599 ();
 sg13g2_decap_8 FILLER_177_1606 ();
 sg13g2_decap_8 FILLER_177_1613 ();
 sg13g2_decap_4 FILLER_177_1620 ();
 sg13g2_fill_1 FILLER_177_1624 ();
 sg13g2_decap_8 FILLER_178_0 ();
 sg13g2_decap_8 FILLER_178_7 ();
 sg13g2_decap_8 FILLER_178_14 ();
 sg13g2_decap_8 FILLER_178_21 ();
 sg13g2_decap_8 FILLER_178_28 ();
 sg13g2_decap_8 FILLER_178_35 ();
 sg13g2_decap_8 FILLER_178_42 ();
 sg13g2_decap_8 FILLER_178_49 ();
 sg13g2_decap_8 FILLER_178_56 ();
 sg13g2_decap_8 FILLER_178_63 ();
 sg13g2_decap_8 FILLER_178_70 ();
 sg13g2_decap_8 FILLER_178_77 ();
 sg13g2_decap_8 FILLER_178_84 ();
 sg13g2_decap_8 FILLER_178_91 ();
 sg13g2_decap_8 FILLER_178_98 ();
 sg13g2_decap_8 FILLER_178_105 ();
 sg13g2_decap_8 FILLER_178_112 ();
 sg13g2_decap_8 FILLER_178_119 ();
 sg13g2_decap_8 FILLER_178_126 ();
 sg13g2_decap_8 FILLER_178_133 ();
 sg13g2_decap_8 FILLER_178_140 ();
 sg13g2_decap_8 FILLER_178_147 ();
 sg13g2_decap_8 FILLER_178_154 ();
 sg13g2_decap_8 FILLER_178_161 ();
 sg13g2_decap_8 FILLER_178_168 ();
 sg13g2_decap_8 FILLER_178_175 ();
 sg13g2_decap_8 FILLER_178_182 ();
 sg13g2_decap_8 FILLER_178_189 ();
 sg13g2_decap_8 FILLER_178_196 ();
 sg13g2_decap_8 FILLER_178_203 ();
 sg13g2_fill_1 FILLER_178_210 ();
 sg13g2_decap_4 FILLER_178_237 ();
 sg13g2_fill_2 FILLER_178_249 ();
 sg13g2_fill_1 FILLER_178_251 ();
 sg13g2_decap_8 FILLER_178_256 ();
 sg13g2_decap_8 FILLER_178_263 ();
 sg13g2_fill_2 FILLER_178_270 ();
 sg13g2_decap_4 FILLER_178_277 ();
 sg13g2_fill_2 FILLER_178_281 ();
 sg13g2_decap_8 FILLER_178_296 ();
 sg13g2_fill_2 FILLER_178_303 ();
 sg13g2_decap_8 FILLER_178_331 ();
 sg13g2_fill_1 FILLER_178_338 ();
 sg13g2_decap_8 FILLER_178_344 ();
 sg13g2_fill_2 FILLER_178_351 ();
 sg13g2_decap_8 FILLER_178_365 ();
 sg13g2_decap_8 FILLER_178_441 ();
 sg13g2_fill_1 FILLER_178_448 ();
 sg13g2_decap_4 FILLER_178_453 ();
 sg13g2_decap_4 FILLER_178_461 ();
 sg13g2_fill_1 FILLER_178_465 ();
 sg13g2_fill_1 FILLER_178_501 ();
 sg13g2_decap_4 FILLER_178_511 ();
 sg13g2_fill_1 FILLER_178_515 ();
 sg13g2_decap_8 FILLER_178_525 ();
 sg13g2_decap_8 FILLER_178_532 ();
 sg13g2_fill_2 FILLER_178_539 ();
 sg13g2_decap_8 FILLER_178_544 ();
 sg13g2_decap_8 FILLER_178_551 ();
 sg13g2_decap_4 FILLER_178_558 ();
 sg13g2_fill_2 FILLER_178_601 ();
 sg13g2_fill_2 FILLER_178_629 ();
 sg13g2_fill_1 FILLER_178_631 ();
 sg13g2_fill_2 FILLER_178_637 ();
 sg13g2_fill_1 FILLER_178_639 ();
 sg13g2_fill_2 FILLER_178_644 ();
 sg13g2_fill_1 FILLER_178_646 ();
 sg13g2_decap_8 FILLER_178_682 ();
 sg13g2_decap_4 FILLER_178_689 ();
 sg13g2_fill_2 FILLER_178_693 ();
 sg13g2_decap_4 FILLER_178_752 ();
 sg13g2_fill_1 FILLER_178_760 ();
 sg13g2_decap_8 FILLER_178_765 ();
 sg13g2_decap_8 FILLER_178_772 ();
 sg13g2_decap_4 FILLER_178_779 ();
 sg13g2_decap_8 FILLER_178_808 ();
 sg13g2_decap_8 FILLER_178_815 ();
 sg13g2_decap_8 FILLER_178_822 ();
 sg13g2_decap_8 FILLER_178_829 ();
 sg13g2_fill_2 FILLER_178_836 ();
 sg13g2_decap_8 FILLER_178_846 ();
 sg13g2_decap_4 FILLER_178_853 ();
 sg13g2_fill_2 FILLER_178_857 ();
 sg13g2_fill_2 FILLER_178_865 ();
 sg13g2_fill_1 FILLER_178_867 ();
 sg13g2_decap_4 FILLER_178_872 ();
 sg13g2_fill_1 FILLER_178_876 ();
 sg13g2_decap_8 FILLER_178_881 ();
 sg13g2_decap_8 FILLER_178_888 ();
 sg13g2_decap_8 FILLER_178_895 ();
 sg13g2_fill_2 FILLER_178_902 ();
 sg13g2_fill_2 FILLER_178_935 ();
 sg13g2_fill_2 FILLER_178_1011 ();
 sg13g2_fill_1 FILLER_178_1013 ();
 sg13g2_decap_8 FILLER_178_1018 ();
 sg13g2_decap_8 FILLER_178_1025 ();
 sg13g2_decap_4 FILLER_178_1032 ();
 sg13g2_fill_2 FILLER_178_1036 ();
 sg13g2_fill_1 FILLER_178_1075 ();
 sg13g2_decap_4 FILLER_178_1110 ();
 sg13g2_fill_2 FILLER_178_1114 ();
 sg13g2_fill_2 FILLER_178_1122 ();
 sg13g2_fill_1 FILLER_178_1124 ();
 sg13g2_fill_2 FILLER_178_1137 ();
 sg13g2_fill_1 FILLER_178_1139 ();
 sg13g2_decap_8 FILLER_178_1229 ();
 sg13g2_decap_8 FILLER_178_1236 ();
 sg13g2_fill_2 FILLER_178_1243 ();
 sg13g2_fill_2 FILLER_178_1257 ();
 sg13g2_decap_4 FILLER_178_1263 ();
 sg13g2_fill_2 FILLER_178_1267 ();
 sg13g2_decap_4 FILLER_178_1285 ();
 sg13g2_fill_2 FILLER_178_1289 ();
 sg13g2_decap_8 FILLER_178_1295 ();
 sg13g2_decap_8 FILLER_178_1302 ();
 sg13g2_decap_8 FILLER_178_1309 ();
 sg13g2_decap_8 FILLER_178_1316 ();
 sg13g2_decap_8 FILLER_178_1323 ();
 sg13g2_decap_8 FILLER_178_1330 ();
 sg13g2_decap_8 FILLER_178_1337 ();
 sg13g2_decap_8 FILLER_178_1344 ();
 sg13g2_decap_8 FILLER_178_1351 ();
 sg13g2_decap_8 FILLER_178_1358 ();
 sg13g2_decap_8 FILLER_178_1365 ();
 sg13g2_decap_8 FILLER_178_1372 ();
 sg13g2_decap_8 FILLER_178_1379 ();
 sg13g2_decap_8 FILLER_178_1386 ();
 sg13g2_decap_8 FILLER_178_1393 ();
 sg13g2_decap_8 FILLER_178_1400 ();
 sg13g2_decap_8 FILLER_178_1407 ();
 sg13g2_decap_8 FILLER_178_1414 ();
 sg13g2_decap_8 FILLER_178_1421 ();
 sg13g2_decap_8 FILLER_178_1428 ();
 sg13g2_decap_8 FILLER_178_1435 ();
 sg13g2_decap_8 FILLER_178_1442 ();
 sg13g2_decap_8 FILLER_178_1449 ();
 sg13g2_decap_8 FILLER_178_1456 ();
 sg13g2_decap_8 FILLER_178_1463 ();
 sg13g2_decap_8 FILLER_178_1470 ();
 sg13g2_decap_8 FILLER_178_1477 ();
 sg13g2_decap_8 FILLER_178_1484 ();
 sg13g2_decap_8 FILLER_178_1491 ();
 sg13g2_decap_8 FILLER_178_1498 ();
 sg13g2_decap_8 FILLER_178_1505 ();
 sg13g2_decap_8 FILLER_178_1512 ();
 sg13g2_decap_8 FILLER_178_1519 ();
 sg13g2_decap_8 FILLER_178_1526 ();
 sg13g2_decap_8 FILLER_178_1533 ();
 sg13g2_decap_8 FILLER_178_1540 ();
 sg13g2_decap_8 FILLER_178_1547 ();
 sg13g2_decap_8 FILLER_178_1554 ();
 sg13g2_decap_8 FILLER_178_1561 ();
 sg13g2_decap_8 FILLER_178_1568 ();
 sg13g2_decap_8 FILLER_178_1575 ();
 sg13g2_decap_8 FILLER_178_1582 ();
 sg13g2_decap_8 FILLER_178_1589 ();
 sg13g2_decap_8 FILLER_178_1596 ();
 sg13g2_decap_8 FILLER_178_1603 ();
 sg13g2_decap_8 FILLER_178_1610 ();
 sg13g2_decap_8 FILLER_178_1617 ();
 sg13g2_fill_1 FILLER_178_1624 ();
 sg13g2_decap_8 FILLER_179_0 ();
 sg13g2_decap_8 FILLER_179_7 ();
 sg13g2_decap_8 FILLER_179_14 ();
 sg13g2_decap_8 FILLER_179_21 ();
 sg13g2_decap_8 FILLER_179_28 ();
 sg13g2_decap_8 FILLER_179_35 ();
 sg13g2_decap_8 FILLER_179_42 ();
 sg13g2_decap_8 FILLER_179_49 ();
 sg13g2_decap_8 FILLER_179_56 ();
 sg13g2_decap_8 FILLER_179_63 ();
 sg13g2_decap_8 FILLER_179_70 ();
 sg13g2_decap_8 FILLER_179_77 ();
 sg13g2_decap_8 FILLER_179_84 ();
 sg13g2_decap_8 FILLER_179_91 ();
 sg13g2_decap_8 FILLER_179_98 ();
 sg13g2_decap_8 FILLER_179_105 ();
 sg13g2_decap_8 FILLER_179_112 ();
 sg13g2_decap_8 FILLER_179_119 ();
 sg13g2_decap_8 FILLER_179_126 ();
 sg13g2_decap_8 FILLER_179_133 ();
 sg13g2_decap_8 FILLER_179_140 ();
 sg13g2_decap_8 FILLER_179_147 ();
 sg13g2_decap_8 FILLER_179_154 ();
 sg13g2_decap_8 FILLER_179_161 ();
 sg13g2_decap_8 FILLER_179_168 ();
 sg13g2_decap_8 FILLER_179_175 ();
 sg13g2_decap_8 FILLER_179_182 ();
 sg13g2_decap_8 FILLER_179_189 ();
 sg13g2_decap_8 FILLER_179_196 ();
 sg13g2_decap_8 FILLER_179_203 ();
 sg13g2_decap_8 FILLER_179_210 ();
 sg13g2_decap_8 FILLER_179_217 ();
 sg13g2_decap_8 FILLER_179_224 ();
 sg13g2_decap_8 FILLER_179_231 ();
 sg13g2_fill_2 FILLER_179_238 ();
 sg13g2_decap_4 FILLER_179_270 ();
 sg13g2_fill_1 FILLER_179_274 ();
 sg13g2_decap_4 FILLER_179_306 ();
 sg13g2_fill_2 FILLER_179_310 ();
 sg13g2_decap_8 FILLER_179_316 ();
 sg13g2_decap_8 FILLER_179_323 ();
 sg13g2_decap_4 FILLER_179_330 ();
 sg13g2_fill_1 FILLER_179_334 ();
 sg13g2_fill_2 FILLER_179_343 ();
 sg13g2_decap_8 FILLER_179_354 ();
 sg13g2_fill_1 FILLER_179_361 ();
 sg13g2_decap_4 FILLER_179_366 ();
 sg13g2_fill_2 FILLER_179_370 ();
 sg13g2_decap_4 FILLER_179_405 ();
 sg13g2_fill_2 FILLER_179_414 ();
 sg13g2_decap_4 FILLER_179_445 ();
 sg13g2_fill_2 FILLER_179_453 ();
 sg13g2_decap_8 FILLER_179_459 ();
 sg13g2_fill_1 FILLER_179_466 ();
 sg13g2_fill_1 FILLER_179_472 ();
 sg13g2_decap_8 FILLER_179_477 ();
 sg13g2_decap_4 FILLER_179_484 ();
 sg13g2_decap_4 FILLER_179_492 ();
 sg13g2_decap_8 FILLER_179_526 ();
 sg13g2_decap_8 FILLER_179_538 ();
 sg13g2_decap_8 FILLER_179_545 ();
 sg13g2_fill_2 FILLER_179_552 ();
 sg13g2_decap_8 FILLER_179_563 ();
 sg13g2_decap_4 FILLER_179_570 ();
 sg13g2_decap_8 FILLER_179_583 ();
 sg13g2_decap_4 FILLER_179_590 ();
 sg13g2_fill_2 FILLER_179_594 ();
 sg13g2_decap_8 FILLER_179_601 ();
 sg13g2_decap_8 FILLER_179_608 ();
 sg13g2_decap_8 FILLER_179_615 ();
 sg13g2_fill_2 FILLER_179_622 ();
 sg13g2_fill_2 FILLER_179_659 ();
 sg13g2_decap_8 FILLER_179_665 ();
 sg13g2_decap_8 FILLER_179_672 ();
 sg13g2_fill_2 FILLER_179_679 ();
 sg13g2_fill_1 FILLER_179_681 ();
 sg13g2_decap_4 FILLER_179_724 ();
 sg13g2_fill_2 FILLER_179_728 ();
 sg13g2_fill_2 FILLER_179_734 ();
 sg13g2_fill_1 FILLER_179_736 ();
 sg13g2_decap_8 FILLER_179_791 ();
 sg13g2_decap_8 FILLER_179_798 ();
 sg13g2_decap_8 FILLER_179_805 ();
 sg13g2_decap_8 FILLER_179_812 ();
 sg13g2_decap_8 FILLER_179_819 ();
 sg13g2_decap_8 FILLER_179_826 ();
 sg13g2_decap_8 FILLER_179_833 ();
 sg13g2_decap_8 FILLER_179_840 ();
 sg13g2_decap_8 FILLER_179_847 ();
 sg13g2_decap_4 FILLER_179_854 ();
 sg13g2_fill_2 FILLER_179_858 ();
 sg13g2_decap_8 FILLER_179_898 ();
 sg13g2_decap_4 FILLER_179_905 ();
 sg13g2_fill_2 FILLER_179_909 ();
 sg13g2_decap_8 FILLER_179_915 ();
 sg13g2_decap_4 FILLER_179_922 ();
 sg13g2_fill_1 FILLER_179_951 ();
 sg13g2_fill_1 FILLER_179_957 ();
 sg13g2_decap_8 FILLER_179_994 ();
 sg13g2_fill_1 FILLER_179_1031 ();
 sg13g2_decap_8 FILLER_179_1046 ();
 sg13g2_decap_8 FILLER_179_1053 ();
 sg13g2_decap_8 FILLER_179_1060 ();
 sg13g2_decap_8 FILLER_179_1067 ();
 sg13g2_fill_2 FILLER_179_1074 ();
 sg13g2_fill_2 FILLER_179_1109 ();
 sg13g2_fill_1 FILLER_179_1168 ();
 sg13g2_decap_8 FILLER_179_1235 ();
 sg13g2_decap_8 FILLER_179_1242 ();
 sg13g2_fill_2 FILLER_179_1249 ();
 sg13g2_decap_4 FILLER_179_1277 ();
 sg13g2_fill_2 FILLER_179_1281 ();
 sg13g2_decap_8 FILLER_179_1309 ();
 sg13g2_decap_8 FILLER_179_1316 ();
 sg13g2_decap_8 FILLER_179_1323 ();
 sg13g2_decap_8 FILLER_179_1330 ();
 sg13g2_decap_8 FILLER_179_1337 ();
 sg13g2_decap_8 FILLER_179_1344 ();
 sg13g2_decap_8 FILLER_179_1351 ();
 sg13g2_decap_8 FILLER_179_1358 ();
 sg13g2_decap_8 FILLER_179_1365 ();
 sg13g2_decap_8 FILLER_179_1372 ();
 sg13g2_decap_8 FILLER_179_1379 ();
 sg13g2_decap_8 FILLER_179_1386 ();
 sg13g2_decap_8 FILLER_179_1393 ();
 sg13g2_decap_8 FILLER_179_1400 ();
 sg13g2_decap_8 FILLER_179_1407 ();
 sg13g2_decap_8 FILLER_179_1414 ();
 sg13g2_decap_8 FILLER_179_1421 ();
 sg13g2_decap_8 FILLER_179_1428 ();
 sg13g2_decap_8 FILLER_179_1435 ();
 sg13g2_decap_8 FILLER_179_1442 ();
 sg13g2_decap_8 FILLER_179_1449 ();
 sg13g2_decap_8 FILLER_179_1456 ();
 sg13g2_decap_8 FILLER_179_1463 ();
 sg13g2_decap_8 FILLER_179_1470 ();
 sg13g2_decap_8 FILLER_179_1477 ();
 sg13g2_decap_8 FILLER_179_1484 ();
 sg13g2_decap_8 FILLER_179_1491 ();
 sg13g2_decap_8 FILLER_179_1498 ();
 sg13g2_decap_8 FILLER_179_1505 ();
 sg13g2_decap_8 FILLER_179_1512 ();
 sg13g2_decap_8 FILLER_179_1519 ();
 sg13g2_decap_8 FILLER_179_1526 ();
 sg13g2_decap_8 FILLER_179_1533 ();
 sg13g2_decap_8 FILLER_179_1540 ();
 sg13g2_decap_8 FILLER_179_1547 ();
 sg13g2_decap_8 FILLER_179_1554 ();
 sg13g2_decap_8 FILLER_179_1561 ();
 sg13g2_decap_8 FILLER_179_1568 ();
 sg13g2_decap_8 FILLER_179_1575 ();
 sg13g2_decap_8 FILLER_179_1582 ();
 sg13g2_decap_8 FILLER_179_1589 ();
 sg13g2_decap_8 FILLER_179_1596 ();
 sg13g2_decap_8 FILLER_179_1603 ();
 sg13g2_decap_8 FILLER_179_1610 ();
 sg13g2_decap_8 FILLER_179_1617 ();
 sg13g2_fill_1 FILLER_179_1624 ();
 sg13g2_decap_8 FILLER_180_0 ();
 sg13g2_decap_8 FILLER_180_7 ();
 sg13g2_decap_8 FILLER_180_14 ();
 sg13g2_decap_8 FILLER_180_21 ();
 sg13g2_decap_8 FILLER_180_28 ();
 sg13g2_decap_8 FILLER_180_35 ();
 sg13g2_decap_8 FILLER_180_42 ();
 sg13g2_decap_8 FILLER_180_49 ();
 sg13g2_decap_8 FILLER_180_56 ();
 sg13g2_decap_8 FILLER_180_63 ();
 sg13g2_decap_8 FILLER_180_70 ();
 sg13g2_decap_8 FILLER_180_77 ();
 sg13g2_decap_8 FILLER_180_84 ();
 sg13g2_decap_8 FILLER_180_91 ();
 sg13g2_decap_8 FILLER_180_98 ();
 sg13g2_decap_8 FILLER_180_105 ();
 sg13g2_decap_8 FILLER_180_112 ();
 sg13g2_decap_8 FILLER_180_119 ();
 sg13g2_decap_8 FILLER_180_126 ();
 sg13g2_decap_8 FILLER_180_133 ();
 sg13g2_decap_8 FILLER_180_140 ();
 sg13g2_decap_8 FILLER_180_147 ();
 sg13g2_decap_8 FILLER_180_154 ();
 sg13g2_decap_8 FILLER_180_161 ();
 sg13g2_decap_8 FILLER_180_168 ();
 sg13g2_decap_8 FILLER_180_175 ();
 sg13g2_decap_8 FILLER_180_182 ();
 sg13g2_decap_8 FILLER_180_189 ();
 sg13g2_decap_8 FILLER_180_196 ();
 sg13g2_decap_8 FILLER_180_203 ();
 sg13g2_decap_8 FILLER_180_210 ();
 sg13g2_decap_8 FILLER_180_217 ();
 sg13g2_decap_8 FILLER_180_224 ();
 sg13g2_decap_8 FILLER_180_231 ();
 sg13g2_decap_8 FILLER_180_238 ();
 sg13g2_decap_8 FILLER_180_245 ();
 sg13g2_decap_8 FILLER_180_252 ();
 sg13g2_decap_4 FILLER_180_259 ();
 sg13g2_decap_8 FILLER_180_283 ();
 sg13g2_decap_8 FILLER_180_290 ();
 sg13g2_fill_2 FILLER_180_297 ();
 sg13g2_fill_2 FILLER_180_303 ();
 sg13g2_decap_8 FILLER_180_310 ();
 sg13g2_decap_4 FILLER_180_317 ();
 sg13g2_fill_2 FILLER_180_325 ();
 sg13g2_fill_1 FILLER_180_331 ();
 sg13g2_fill_2 FILLER_180_358 ();
 sg13g2_fill_1 FILLER_180_360 ();
 sg13g2_fill_2 FILLER_180_461 ();
 sg13g2_fill_1 FILLER_180_463 ();
 sg13g2_decap_8 FILLER_180_509 ();
 sg13g2_decap_8 FILLER_180_516 ();
 sg13g2_decap_8 FILLER_180_580 ();
 sg13g2_decap_4 FILLER_180_587 ();
 sg13g2_fill_1 FILLER_180_591 ();
 sg13g2_decap_8 FILLER_180_596 ();
 sg13g2_decap_8 FILLER_180_603 ();
 sg13g2_decap_8 FILLER_180_610 ();
 sg13g2_decap_8 FILLER_180_617 ();
 sg13g2_decap_4 FILLER_180_624 ();
 sg13g2_fill_1 FILLER_180_628 ();
 sg13g2_decap_8 FILLER_180_634 ();
 sg13g2_decap_8 FILLER_180_641 ();
 sg13g2_fill_2 FILLER_180_648 ();
 sg13g2_fill_1 FILLER_180_650 ();
 sg13g2_decap_8 FILLER_180_702 ();
 sg13g2_decap_8 FILLER_180_709 ();
 sg13g2_decap_4 FILLER_180_716 ();
 sg13g2_fill_2 FILLER_180_720 ();
 sg13g2_fill_2 FILLER_180_753 ();
 sg13g2_decap_8 FILLER_180_781 ();
 sg13g2_decap_8 FILLER_180_788 ();
 sg13g2_decap_8 FILLER_180_795 ();
 sg13g2_decap_8 FILLER_180_802 ();
 sg13g2_decap_4 FILLER_180_809 ();
 sg13g2_decap_8 FILLER_180_817 ();
 sg13g2_fill_1 FILLER_180_854 ();
 sg13g2_fill_1 FILLER_180_871 ();
 sg13g2_fill_1 FILLER_180_880 ();
 sg13g2_fill_1 FILLER_180_885 ();
 sg13g2_decap_8 FILLER_180_912 ();
 sg13g2_decap_8 FILLER_180_919 ();
 sg13g2_decap_8 FILLER_180_926 ();
 sg13g2_decap_4 FILLER_180_988 ();
 sg13g2_decap_8 FILLER_180_998 ();
 sg13g2_decap_8 FILLER_180_1005 ();
 sg13g2_decap_4 FILLER_180_1022 ();
 sg13g2_fill_1 FILLER_180_1026 ();
 sg13g2_decap_8 FILLER_180_1033 ();
 sg13g2_decap_4 FILLER_180_1044 ();
 sg13g2_fill_1 FILLER_180_1048 ();
 sg13g2_fill_1 FILLER_180_1055 ();
 sg13g2_fill_1 FILLER_180_1062 ();
 sg13g2_fill_1 FILLER_180_1069 ();
 sg13g2_fill_1 FILLER_180_1075 ();
 sg13g2_fill_2 FILLER_180_1082 ();
 sg13g2_fill_2 FILLER_180_1193 ();
 sg13g2_decap_8 FILLER_180_1234 ();
 sg13g2_decap_8 FILLER_180_1241 ();
 sg13g2_decap_8 FILLER_180_1248 ();
 sg13g2_decap_8 FILLER_180_1255 ();
 sg13g2_decap_8 FILLER_180_1262 ();
 sg13g2_fill_2 FILLER_180_1269 ();
 sg13g2_fill_1 FILLER_180_1271 ();
 sg13g2_decap_8 FILLER_180_1297 ();
 sg13g2_decap_8 FILLER_180_1304 ();
 sg13g2_decap_8 FILLER_180_1311 ();
 sg13g2_decap_8 FILLER_180_1318 ();
 sg13g2_decap_8 FILLER_180_1325 ();
 sg13g2_decap_8 FILLER_180_1332 ();
 sg13g2_decap_8 FILLER_180_1339 ();
 sg13g2_decap_8 FILLER_180_1346 ();
 sg13g2_decap_8 FILLER_180_1353 ();
 sg13g2_decap_8 FILLER_180_1360 ();
 sg13g2_decap_8 FILLER_180_1367 ();
 sg13g2_decap_8 FILLER_180_1374 ();
 sg13g2_decap_8 FILLER_180_1381 ();
 sg13g2_decap_8 FILLER_180_1388 ();
 sg13g2_decap_8 FILLER_180_1395 ();
 sg13g2_decap_8 FILLER_180_1402 ();
 sg13g2_decap_8 FILLER_180_1409 ();
 sg13g2_decap_8 FILLER_180_1416 ();
 sg13g2_decap_8 FILLER_180_1423 ();
 sg13g2_decap_8 FILLER_180_1430 ();
 sg13g2_decap_8 FILLER_180_1437 ();
 sg13g2_decap_8 FILLER_180_1444 ();
 sg13g2_decap_8 FILLER_180_1451 ();
 sg13g2_decap_8 FILLER_180_1458 ();
 sg13g2_decap_8 FILLER_180_1465 ();
 sg13g2_decap_8 FILLER_180_1472 ();
 sg13g2_decap_8 FILLER_180_1479 ();
 sg13g2_decap_8 FILLER_180_1486 ();
 sg13g2_decap_8 FILLER_180_1493 ();
 sg13g2_decap_8 FILLER_180_1500 ();
 sg13g2_decap_8 FILLER_180_1507 ();
 sg13g2_decap_8 FILLER_180_1514 ();
 sg13g2_decap_8 FILLER_180_1521 ();
 sg13g2_decap_8 FILLER_180_1528 ();
 sg13g2_decap_8 FILLER_180_1535 ();
 sg13g2_decap_8 FILLER_180_1542 ();
 sg13g2_decap_8 FILLER_180_1549 ();
 sg13g2_decap_8 FILLER_180_1556 ();
 sg13g2_decap_8 FILLER_180_1563 ();
 sg13g2_decap_8 FILLER_180_1570 ();
 sg13g2_decap_8 FILLER_180_1577 ();
 sg13g2_decap_8 FILLER_180_1584 ();
 sg13g2_decap_8 FILLER_180_1591 ();
 sg13g2_decap_8 FILLER_180_1598 ();
 sg13g2_decap_8 FILLER_180_1605 ();
 sg13g2_decap_8 FILLER_180_1612 ();
 sg13g2_decap_4 FILLER_180_1619 ();
 sg13g2_fill_2 FILLER_180_1623 ();
 sg13g2_decap_8 FILLER_181_0 ();
 sg13g2_decap_8 FILLER_181_7 ();
 sg13g2_decap_8 FILLER_181_14 ();
 sg13g2_decap_8 FILLER_181_21 ();
 sg13g2_decap_8 FILLER_181_28 ();
 sg13g2_decap_8 FILLER_181_35 ();
 sg13g2_decap_8 FILLER_181_42 ();
 sg13g2_decap_8 FILLER_181_49 ();
 sg13g2_decap_8 FILLER_181_56 ();
 sg13g2_decap_8 FILLER_181_63 ();
 sg13g2_decap_8 FILLER_181_70 ();
 sg13g2_decap_8 FILLER_181_77 ();
 sg13g2_decap_8 FILLER_181_84 ();
 sg13g2_decap_8 FILLER_181_91 ();
 sg13g2_decap_8 FILLER_181_98 ();
 sg13g2_decap_8 FILLER_181_105 ();
 sg13g2_decap_8 FILLER_181_112 ();
 sg13g2_decap_8 FILLER_181_119 ();
 sg13g2_decap_8 FILLER_181_126 ();
 sg13g2_decap_8 FILLER_181_133 ();
 sg13g2_decap_8 FILLER_181_140 ();
 sg13g2_decap_8 FILLER_181_147 ();
 sg13g2_decap_8 FILLER_181_154 ();
 sg13g2_decap_8 FILLER_181_161 ();
 sg13g2_decap_8 FILLER_181_168 ();
 sg13g2_decap_8 FILLER_181_175 ();
 sg13g2_decap_8 FILLER_181_182 ();
 sg13g2_decap_8 FILLER_181_189 ();
 sg13g2_decap_8 FILLER_181_196 ();
 sg13g2_decap_8 FILLER_181_203 ();
 sg13g2_decap_8 FILLER_181_210 ();
 sg13g2_decap_8 FILLER_181_217 ();
 sg13g2_decap_8 FILLER_181_224 ();
 sg13g2_decap_8 FILLER_181_231 ();
 sg13g2_decap_8 FILLER_181_238 ();
 sg13g2_fill_2 FILLER_181_274 ();
 sg13g2_fill_1 FILLER_181_276 ();
 sg13g2_fill_2 FILLER_181_287 ();
 sg13g2_fill_1 FILLER_181_289 ();
 sg13g2_fill_1 FILLER_181_299 ();
 sg13g2_fill_1 FILLER_181_315 ();
 sg13g2_fill_2 FILLER_181_330 ();
 sg13g2_fill_1 FILLER_181_332 ();
 sg13g2_fill_2 FILLER_181_343 ();
 sg13g2_decap_8 FILLER_181_376 ();
 sg13g2_fill_2 FILLER_181_383 ();
 sg13g2_fill_1 FILLER_181_385 ();
 sg13g2_decap_8 FILLER_181_392 ();
 sg13g2_fill_2 FILLER_181_399 ();
 sg13g2_decap_8 FILLER_181_431 ();
 sg13g2_decap_8 FILLER_181_438 ();
 sg13g2_fill_1 FILLER_181_445 ();
 sg13g2_fill_1 FILLER_181_451 ();
 sg13g2_fill_1 FILLER_181_491 ();
 sg13g2_decap_8 FILLER_181_504 ();
 sg13g2_decap_8 FILLER_181_511 ();
 sg13g2_fill_2 FILLER_181_518 ();
 sg13g2_fill_1 FILLER_181_520 ();
 sg13g2_fill_1 FILLER_181_552 ();
 sg13g2_decap_4 FILLER_181_557 ();
 sg13g2_fill_1 FILLER_181_561 ();
 sg13g2_decap_8 FILLER_181_566 ();
 sg13g2_fill_2 FILLER_181_573 ();
 sg13g2_decap_4 FILLER_181_580 ();
 sg13g2_fill_1 FILLER_181_584 ();
 sg13g2_decap_8 FILLER_181_624 ();
 sg13g2_decap_8 FILLER_181_631 ();
 sg13g2_decap_8 FILLER_181_638 ();
 sg13g2_decap_4 FILLER_181_645 ();
 sg13g2_fill_1 FILLER_181_649 ();
 sg13g2_fill_2 FILLER_181_685 ();
 sg13g2_fill_1 FILLER_181_687 ();
 sg13g2_decap_4 FILLER_181_717 ();
 sg13g2_decap_8 FILLER_181_730 ();
 sg13g2_fill_2 FILLER_181_737 ();
 sg13g2_fill_1 FILLER_181_739 ();
 sg13g2_fill_2 FILLER_181_749 ();
 sg13g2_decap_8 FILLER_181_777 ();
 sg13g2_decap_8 FILLER_181_784 ();
 sg13g2_decap_8 FILLER_181_791 ();
 sg13g2_decap_8 FILLER_181_798 ();
 sg13g2_fill_1 FILLER_181_805 ();
 sg13g2_fill_1 FILLER_181_841 ();
 sg13g2_decap_4 FILLER_181_846 ();
 sg13g2_fill_1 FILLER_181_850 ();
 sg13g2_decap_4 FILLER_181_877 ();
 sg13g2_decap_4 FILLER_181_884 ();
 sg13g2_fill_2 FILLER_181_888 ();
 sg13g2_decap_8 FILLER_181_897 ();
 sg13g2_fill_1 FILLER_181_904 ();
 sg13g2_decap_8 FILLER_181_930 ();
 sg13g2_fill_2 FILLER_181_937 ();
 sg13g2_decap_4 FILLER_181_943 ();
 sg13g2_fill_1 FILLER_181_947 ();
 sg13g2_fill_1 FILLER_181_952 ();
 sg13g2_decap_4 FILLER_181_1037 ();
 sg13g2_fill_1 FILLER_181_1041 ();
 sg13g2_decap_4 FILLER_181_1059 ();
 sg13g2_fill_2 FILLER_181_1063 ();
 sg13g2_decap_8 FILLER_181_1069 ();
 sg13g2_decap_4 FILLER_181_1076 ();
 sg13g2_fill_2 FILLER_181_1080 ();
 sg13g2_fill_2 FILLER_181_1094 ();
 sg13g2_fill_1 FILLER_181_1130 ();
 sg13g2_fill_2 FILLER_181_1163 ();
 sg13g2_fill_1 FILLER_181_1165 ();
 sg13g2_fill_2 FILLER_181_1214 ();
 sg13g2_fill_1 FILLER_181_1216 ();
 sg13g2_decap_8 FILLER_181_1221 ();
 sg13g2_decap_8 FILLER_181_1228 ();
 sg13g2_decap_8 FILLER_181_1235 ();
 sg13g2_decap_8 FILLER_181_1242 ();
 sg13g2_decap_8 FILLER_181_1249 ();
 sg13g2_decap_8 FILLER_181_1256 ();
 sg13g2_decap_8 FILLER_181_1263 ();
 sg13g2_decap_8 FILLER_181_1270 ();
 sg13g2_decap_8 FILLER_181_1277 ();
 sg13g2_decap_8 FILLER_181_1284 ();
 sg13g2_decap_8 FILLER_181_1291 ();
 sg13g2_decap_8 FILLER_181_1298 ();
 sg13g2_decap_8 FILLER_181_1305 ();
 sg13g2_decap_8 FILLER_181_1312 ();
 sg13g2_decap_8 FILLER_181_1319 ();
 sg13g2_decap_8 FILLER_181_1326 ();
 sg13g2_decap_8 FILLER_181_1333 ();
 sg13g2_decap_8 FILLER_181_1340 ();
 sg13g2_decap_8 FILLER_181_1347 ();
 sg13g2_decap_8 FILLER_181_1354 ();
 sg13g2_decap_8 FILLER_181_1361 ();
 sg13g2_decap_8 FILLER_181_1368 ();
 sg13g2_decap_8 FILLER_181_1375 ();
 sg13g2_decap_8 FILLER_181_1382 ();
 sg13g2_decap_8 FILLER_181_1389 ();
 sg13g2_decap_8 FILLER_181_1396 ();
 sg13g2_decap_8 FILLER_181_1403 ();
 sg13g2_decap_8 FILLER_181_1410 ();
 sg13g2_decap_8 FILLER_181_1417 ();
 sg13g2_decap_8 FILLER_181_1424 ();
 sg13g2_decap_8 FILLER_181_1431 ();
 sg13g2_decap_8 FILLER_181_1438 ();
 sg13g2_decap_8 FILLER_181_1445 ();
 sg13g2_decap_8 FILLER_181_1452 ();
 sg13g2_decap_8 FILLER_181_1459 ();
 sg13g2_decap_8 FILLER_181_1466 ();
 sg13g2_decap_8 FILLER_181_1473 ();
 sg13g2_decap_8 FILLER_181_1480 ();
 sg13g2_decap_8 FILLER_181_1487 ();
 sg13g2_decap_8 FILLER_181_1494 ();
 sg13g2_decap_8 FILLER_181_1501 ();
 sg13g2_decap_8 FILLER_181_1508 ();
 sg13g2_decap_8 FILLER_181_1515 ();
 sg13g2_decap_8 FILLER_181_1522 ();
 sg13g2_decap_8 FILLER_181_1529 ();
 sg13g2_decap_8 FILLER_181_1536 ();
 sg13g2_decap_8 FILLER_181_1543 ();
 sg13g2_decap_8 FILLER_181_1550 ();
 sg13g2_decap_8 FILLER_181_1557 ();
 sg13g2_decap_8 FILLER_181_1564 ();
 sg13g2_decap_8 FILLER_181_1571 ();
 sg13g2_decap_8 FILLER_181_1578 ();
 sg13g2_decap_8 FILLER_181_1585 ();
 sg13g2_decap_8 FILLER_181_1592 ();
 sg13g2_decap_8 FILLER_181_1599 ();
 sg13g2_decap_8 FILLER_181_1606 ();
 sg13g2_decap_8 FILLER_181_1613 ();
 sg13g2_decap_4 FILLER_181_1620 ();
 sg13g2_fill_1 FILLER_181_1624 ();
 sg13g2_decap_8 FILLER_182_0 ();
 sg13g2_decap_8 FILLER_182_7 ();
 sg13g2_decap_8 FILLER_182_14 ();
 sg13g2_decap_8 FILLER_182_21 ();
 sg13g2_decap_8 FILLER_182_28 ();
 sg13g2_decap_8 FILLER_182_35 ();
 sg13g2_decap_8 FILLER_182_42 ();
 sg13g2_decap_8 FILLER_182_49 ();
 sg13g2_decap_8 FILLER_182_56 ();
 sg13g2_decap_8 FILLER_182_63 ();
 sg13g2_decap_8 FILLER_182_70 ();
 sg13g2_decap_8 FILLER_182_77 ();
 sg13g2_decap_8 FILLER_182_84 ();
 sg13g2_decap_8 FILLER_182_91 ();
 sg13g2_decap_8 FILLER_182_98 ();
 sg13g2_decap_8 FILLER_182_105 ();
 sg13g2_decap_8 FILLER_182_112 ();
 sg13g2_decap_8 FILLER_182_119 ();
 sg13g2_decap_8 FILLER_182_126 ();
 sg13g2_decap_8 FILLER_182_133 ();
 sg13g2_decap_8 FILLER_182_140 ();
 sg13g2_decap_8 FILLER_182_147 ();
 sg13g2_decap_8 FILLER_182_154 ();
 sg13g2_decap_8 FILLER_182_161 ();
 sg13g2_decap_8 FILLER_182_168 ();
 sg13g2_decap_8 FILLER_182_175 ();
 sg13g2_decap_8 FILLER_182_182 ();
 sg13g2_decap_8 FILLER_182_189 ();
 sg13g2_decap_8 FILLER_182_196 ();
 sg13g2_decap_8 FILLER_182_203 ();
 sg13g2_decap_8 FILLER_182_210 ();
 sg13g2_decap_8 FILLER_182_217 ();
 sg13g2_decap_8 FILLER_182_224 ();
 sg13g2_decap_8 FILLER_182_231 ();
 sg13g2_decap_8 FILLER_182_238 ();
 sg13g2_fill_2 FILLER_182_277 ();
 sg13g2_fill_2 FILLER_182_318 ();
 sg13g2_fill_1 FILLER_182_351 ();
 sg13g2_decap_8 FILLER_182_386 ();
 sg13g2_fill_1 FILLER_182_393 ();
 sg13g2_fill_1 FILLER_182_412 ();
 sg13g2_decap_4 FILLER_182_438 ();
 sg13g2_decap_8 FILLER_182_446 ();
 sg13g2_decap_8 FILLER_182_453 ();
 sg13g2_decap_8 FILLER_182_460 ();
 sg13g2_decap_8 FILLER_182_467 ();
 sg13g2_decap_4 FILLER_182_474 ();
 sg13g2_fill_1 FILLER_182_483 ();
 sg13g2_decap_8 FILLER_182_494 ();
 sg13g2_decap_4 FILLER_182_501 ();
 sg13g2_fill_1 FILLER_182_505 ();
 sg13g2_fill_1 FILLER_182_534 ();
 sg13g2_decap_8 FILLER_182_539 ();
 sg13g2_fill_1 FILLER_182_546 ();
 sg13g2_fill_2 FILLER_182_572 ();
 sg13g2_fill_1 FILLER_182_595 ();
 sg13g2_fill_2 FILLER_182_601 ();
 sg13g2_fill_1 FILLER_182_612 ();
 sg13g2_fill_2 FILLER_182_644 ();
 sg13g2_fill_1 FILLER_182_650 ();
 sg13g2_decap_8 FILLER_182_656 ();
 sg13g2_decap_8 FILLER_182_663 ();
 sg13g2_decap_4 FILLER_182_670 ();
 sg13g2_fill_2 FILLER_182_674 ();
 sg13g2_decap_8 FILLER_182_680 ();
 sg13g2_decap_8 FILLER_182_687 ();
 sg13g2_fill_1 FILLER_182_694 ();
 sg13g2_decap_8 FILLER_182_705 ();
 sg13g2_fill_1 FILLER_182_712 ();
 sg13g2_decap_8 FILLER_182_745 ();
 sg13g2_fill_2 FILLER_182_752 ();
 sg13g2_decap_8 FILLER_182_783 ();
 sg13g2_decap_8 FILLER_182_790 ();
 sg13g2_decap_8 FILLER_182_797 ();
 sg13g2_decap_4 FILLER_182_804 ();
 sg13g2_fill_2 FILLER_182_808 ();
 sg13g2_decap_8 FILLER_182_847 ();
 sg13g2_fill_2 FILLER_182_854 ();
 sg13g2_fill_1 FILLER_182_856 ();
 sg13g2_fill_1 FILLER_182_889 ();
 sg13g2_fill_1 FILLER_182_915 ();
 sg13g2_fill_1 FILLER_182_941 ();
 sg13g2_fill_1 FILLER_182_993 ();
 sg13g2_decap_8 FILLER_182_1024 ();
 sg13g2_decap_8 FILLER_182_1031 ();
 sg13g2_decap_4 FILLER_182_1038 ();
 sg13g2_decap_8 FILLER_182_1048 ();
 sg13g2_fill_1 FILLER_182_1055 ();
 sg13g2_decap_8 FILLER_182_1082 ();
 sg13g2_fill_2 FILLER_182_1089 ();
 sg13g2_fill_1 FILLER_182_1091 ();
 sg13g2_fill_2 FILLER_182_1096 ();
 sg13g2_decap_8 FILLER_182_1106 ();
 sg13g2_decap_4 FILLER_182_1113 ();
 sg13g2_decap_8 FILLER_182_1121 ();
 sg13g2_decap_4 FILLER_182_1128 ();
 sg13g2_fill_1 FILLER_182_1132 ();
 sg13g2_decap_8 FILLER_182_1137 ();
 sg13g2_fill_1 FILLER_182_1144 ();
 sg13g2_decap_8 FILLER_182_1149 ();
 sg13g2_decap_4 FILLER_182_1156 ();
 sg13g2_fill_2 FILLER_182_1160 ();
 sg13g2_fill_2 FILLER_182_1188 ();
 sg13g2_decap_8 FILLER_182_1216 ();
 sg13g2_decap_8 FILLER_182_1223 ();
 sg13g2_decap_8 FILLER_182_1230 ();
 sg13g2_decap_8 FILLER_182_1237 ();
 sg13g2_decap_8 FILLER_182_1244 ();
 sg13g2_decap_8 FILLER_182_1251 ();
 sg13g2_decap_8 FILLER_182_1258 ();
 sg13g2_decap_8 FILLER_182_1265 ();
 sg13g2_decap_8 FILLER_182_1272 ();
 sg13g2_decap_8 FILLER_182_1279 ();
 sg13g2_decap_8 FILLER_182_1286 ();
 sg13g2_decap_8 FILLER_182_1293 ();
 sg13g2_decap_8 FILLER_182_1300 ();
 sg13g2_decap_8 FILLER_182_1307 ();
 sg13g2_decap_8 FILLER_182_1314 ();
 sg13g2_decap_8 FILLER_182_1321 ();
 sg13g2_decap_8 FILLER_182_1328 ();
 sg13g2_decap_8 FILLER_182_1335 ();
 sg13g2_decap_8 FILLER_182_1342 ();
 sg13g2_decap_8 FILLER_182_1349 ();
 sg13g2_decap_8 FILLER_182_1356 ();
 sg13g2_decap_8 FILLER_182_1363 ();
 sg13g2_decap_8 FILLER_182_1370 ();
 sg13g2_decap_8 FILLER_182_1377 ();
 sg13g2_decap_8 FILLER_182_1384 ();
 sg13g2_decap_8 FILLER_182_1391 ();
 sg13g2_decap_8 FILLER_182_1398 ();
 sg13g2_decap_8 FILLER_182_1405 ();
 sg13g2_decap_8 FILLER_182_1412 ();
 sg13g2_decap_8 FILLER_182_1419 ();
 sg13g2_decap_8 FILLER_182_1426 ();
 sg13g2_decap_8 FILLER_182_1433 ();
 sg13g2_decap_8 FILLER_182_1440 ();
 sg13g2_decap_8 FILLER_182_1447 ();
 sg13g2_decap_8 FILLER_182_1454 ();
 sg13g2_decap_8 FILLER_182_1461 ();
 sg13g2_decap_8 FILLER_182_1468 ();
 sg13g2_decap_8 FILLER_182_1475 ();
 sg13g2_decap_8 FILLER_182_1482 ();
 sg13g2_decap_8 FILLER_182_1489 ();
 sg13g2_decap_8 FILLER_182_1496 ();
 sg13g2_decap_8 FILLER_182_1503 ();
 sg13g2_decap_8 FILLER_182_1510 ();
 sg13g2_decap_8 FILLER_182_1517 ();
 sg13g2_decap_8 FILLER_182_1524 ();
 sg13g2_decap_8 FILLER_182_1531 ();
 sg13g2_decap_8 FILLER_182_1538 ();
 sg13g2_decap_8 FILLER_182_1545 ();
 sg13g2_decap_8 FILLER_182_1552 ();
 sg13g2_decap_8 FILLER_182_1559 ();
 sg13g2_decap_8 FILLER_182_1566 ();
 sg13g2_decap_8 FILLER_182_1573 ();
 sg13g2_decap_8 FILLER_182_1580 ();
 sg13g2_decap_8 FILLER_182_1587 ();
 sg13g2_decap_8 FILLER_182_1594 ();
 sg13g2_decap_8 FILLER_182_1601 ();
 sg13g2_decap_8 FILLER_182_1608 ();
 sg13g2_decap_8 FILLER_182_1615 ();
 sg13g2_fill_2 FILLER_182_1622 ();
 sg13g2_fill_1 FILLER_182_1624 ();
 sg13g2_decap_8 FILLER_183_0 ();
 sg13g2_decap_8 FILLER_183_7 ();
 sg13g2_decap_8 FILLER_183_14 ();
 sg13g2_decap_8 FILLER_183_21 ();
 sg13g2_decap_8 FILLER_183_28 ();
 sg13g2_decap_8 FILLER_183_35 ();
 sg13g2_decap_8 FILLER_183_42 ();
 sg13g2_decap_8 FILLER_183_49 ();
 sg13g2_decap_8 FILLER_183_56 ();
 sg13g2_decap_8 FILLER_183_63 ();
 sg13g2_decap_8 FILLER_183_70 ();
 sg13g2_decap_8 FILLER_183_77 ();
 sg13g2_decap_8 FILLER_183_84 ();
 sg13g2_decap_8 FILLER_183_91 ();
 sg13g2_decap_8 FILLER_183_98 ();
 sg13g2_decap_8 FILLER_183_105 ();
 sg13g2_decap_8 FILLER_183_112 ();
 sg13g2_decap_8 FILLER_183_119 ();
 sg13g2_decap_8 FILLER_183_126 ();
 sg13g2_decap_8 FILLER_183_133 ();
 sg13g2_decap_8 FILLER_183_140 ();
 sg13g2_decap_8 FILLER_183_147 ();
 sg13g2_decap_8 FILLER_183_154 ();
 sg13g2_decap_8 FILLER_183_161 ();
 sg13g2_decap_8 FILLER_183_168 ();
 sg13g2_decap_8 FILLER_183_175 ();
 sg13g2_decap_8 FILLER_183_182 ();
 sg13g2_decap_8 FILLER_183_189 ();
 sg13g2_decap_8 FILLER_183_196 ();
 sg13g2_decap_8 FILLER_183_203 ();
 sg13g2_decap_8 FILLER_183_210 ();
 sg13g2_decap_8 FILLER_183_217 ();
 sg13g2_decap_8 FILLER_183_224 ();
 sg13g2_decap_8 FILLER_183_231 ();
 sg13g2_decap_8 FILLER_183_238 ();
 sg13g2_fill_2 FILLER_183_245 ();
 sg13g2_fill_1 FILLER_183_247 ();
 sg13g2_decap_8 FILLER_183_252 ();
 sg13g2_decap_8 FILLER_183_259 ();
 sg13g2_decap_4 FILLER_183_266 ();
 sg13g2_fill_2 FILLER_183_270 ();
 sg13g2_decap_4 FILLER_183_278 ();
 sg13g2_fill_1 FILLER_183_282 ();
 sg13g2_fill_1 FILLER_183_287 ();
 sg13g2_fill_2 FILLER_183_292 ();
 sg13g2_decap_8 FILLER_183_372 ();
 sg13g2_decap_8 FILLER_183_379 ();
 sg13g2_decap_8 FILLER_183_386 ();
 sg13g2_fill_1 FILLER_183_393 ();
 sg13g2_fill_2 FILLER_183_399 ();
 sg13g2_fill_1 FILLER_183_401 ();
 sg13g2_fill_1 FILLER_183_447 ();
 sg13g2_fill_2 FILLER_183_453 ();
 sg13g2_decap_8 FILLER_183_496 ();
 sg13g2_fill_2 FILLER_183_503 ();
 sg13g2_fill_1 FILLER_183_535 ();
 sg13g2_fill_2 FILLER_183_571 ();
 sg13g2_fill_1 FILLER_183_573 ();
 sg13g2_fill_1 FILLER_183_638 ();
 sg13g2_fill_2 FILLER_183_643 ();
 sg13g2_fill_2 FILLER_183_654 ();
 sg13g2_fill_1 FILLER_183_656 ();
 sg13g2_fill_1 FILLER_183_662 ();
 sg13g2_decap_8 FILLER_183_668 ();
 sg13g2_fill_2 FILLER_183_675 ();
 sg13g2_fill_1 FILLER_183_677 ();
 sg13g2_decap_8 FILLER_183_682 ();
 sg13g2_fill_2 FILLER_183_689 ();
 sg13g2_fill_2 FILLER_183_700 ();
 sg13g2_fill_1 FILLER_183_702 ();
 sg13g2_decap_8 FILLER_183_734 ();
 sg13g2_decap_4 FILLER_183_741 ();
 sg13g2_fill_1 FILLER_183_745 ();
 sg13g2_decap_8 FILLER_183_751 ();
 sg13g2_fill_2 FILLER_183_758 ();
 sg13g2_fill_1 FILLER_183_760 ();
 sg13g2_decap_8 FILLER_183_765 ();
 sg13g2_decap_8 FILLER_183_772 ();
 sg13g2_decap_8 FILLER_183_779 ();
 sg13g2_decap_8 FILLER_183_786 ();
 sg13g2_decap_8 FILLER_183_793 ();
 sg13g2_decap_8 FILLER_183_800 ();
 sg13g2_fill_2 FILLER_183_807 ();
 sg13g2_fill_1 FILLER_183_809 ();
 sg13g2_decap_8 FILLER_183_843 ();
 sg13g2_decap_4 FILLER_183_850 ();
 sg13g2_fill_2 FILLER_183_854 ();
 sg13g2_decap_8 FILLER_183_860 ();
 sg13g2_decap_8 FILLER_183_867 ();
 sg13g2_fill_1 FILLER_183_874 ();
 sg13g2_decap_4 FILLER_183_911 ();
 sg13g2_fill_1 FILLER_183_915 ();
 sg13g2_decap_8 FILLER_183_926 ();
 sg13g2_decap_8 FILLER_183_933 ();
 sg13g2_decap_8 FILLER_183_940 ();
 sg13g2_fill_2 FILLER_183_947 ();
 sg13g2_decap_4 FILLER_183_953 ();
 sg13g2_decap_4 FILLER_183_1029 ();
 sg13g2_fill_1 FILLER_183_1033 ();
 sg13g2_fill_2 FILLER_183_1046 ();
 sg13g2_decap_8 FILLER_183_1051 ();
 sg13g2_decap_8 FILLER_183_1058 ();
 sg13g2_decap_8 FILLER_183_1065 ();
 sg13g2_decap_8 FILLER_183_1072 ();
 sg13g2_decap_4 FILLER_183_1079 ();
 sg13g2_decap_4 FILLER_183_1105 ();
 sg13g2_decap_8 FILLER_183_1135 ();
 sg13g2_decap_8 FILLER_183_1142 ();
 sg13g2_decap_8 FILLER_183_1149 ();
 sg13g2_decap_8 FILLER_183_1156 ();
 sg13g2_decap_4 FILLER_183_1163 ();
 sg13g2_fill_2 FILLER_183_1167 ();
 sg13g2_decap_8 FILLER_183_1173 ();
 sg13g2_decap_8 FILLER_183_1180 ();
 sg13g2_fill_2 FILLER_183_1187 ();
 sg13g2_decap_8 FILLER_183_1197 ();
 sg13g2_decap_8 FILLER_183_1204 ();
 sg13g2_decap_8 FILLER_183_1211 ();
 sg13g2_decap_8 FILLER_183_1218 ();
 sg13g2_decap_8 FILLER_183_1225 ();
 sg13g2_decap_8 FILLER_183_1232 ();
 sg13g2_decap_8 FILLER_183_1239 ();
 sg13g2_decap_8 FILLER_183_1246 ();
 sg13g2_decap_8 FILLER_183_1253 ();
 sg13g2_decap_8 FILLER_183_1260 ();
 sg13g2_decap_8 FILLER_183_1267 ();
 sg13g2_decap_8 FILLER_183_1274 ();
 sg13g2_decap_8 FILLER_183_1281 ();
 sg13g2_decap_8 FILLER_183_1288 ();
 sg13g2_decap_8 FILLER_183_1295 ();
 sg13g2_decap_8 FILLER_183_1302 ();
 sg13g2_decap_8 FILLER_183_1309 ();
 sg13g2_decap_8 FILLER_183_1316 ();
 sg13g2_decap_8 FILLER_183_1323 ();
 sg13g2_decap_8 FILLER_183_1330 ();
 sg13g2_decap_8 FILLER_183_1337 ();
 sg13g2_decap_8 FILLER_183_1344 ();
 sg13g2_decap_8 FILLER_183_1351 ();
 sg13g2_decap_8 FILLER_183_1358 ();
 sg13g2_decap_8 FILLER_183_1365 ();
 sg13g2_decap_8 FILLER_183_1372 ();
 sg13g2_decap_8 FILLER_183_1379 ();
 sg13g2_decap_8 FILLER_183_1386 ();
 sg13g2_decap_8 FILLER_183_1393 ();
 sg13g2_decap_8 FILLER_183_1400 ();
 sg13g2_decap_8 FILLER_183_1407 ();
 sg13g2_decap_8 FILLER_183_1414 ();
 sg13g2_decap_8 FILLER_183_1421 ();
 sg13g2_decap_8 FILLER_183_1428 ();
 sg13g2_decap_8 FILLER_183_1435 ();
 sg13g2_decap_8 FILLER_183_1442 ();
 sg13g2_decap_8 FILLER_183_1449 ();
 sg13g2_decap_8 FILLER_183_1456 ();
 sg13g2_decap_8 FILLER_183_1463 ();
 sg13g2_decap_8 FILLER_183_1470 ();
 sg13g2_decap_8 FILLER_183_1477 ();
 sg13g2_decap_8 FILLER_183_1484 ();
 sg13g2_decap_8 FILLER_183_1491 ();
 sg13g2_decap_8 FILLER_183_1498 ();
 sg13g2_decap_8 FILLER_183_1505 ();
 sg13g2_decap_8 FILLER_183_1512 ();
 sg13g2_decap_8 FILLER_183_1519 ();
 sg13g2_decap_8 FILLER_183_1526 ();
 sg13g2_decap_8 FILLER_183_1533 ();
 sg13g2_decap_8 FILLER_183_1540 ();
 sg13g2_decap_8 FILLER_183_1547 ();
 sg13g2_decap_8 FILLER_183_1554 ();
 sg13g2_decap_8 FILLER_183_1561 ();
 sg13g2_decap_8 FILLER_183_1568 ();
 sg13g2_decap_8 FILLER_183_1575 ();
 sg13g2_decap_8 FILLER_183_1582 ();
 sg13g2_decap_8 FILLER_183_1589 ();
 sg13g2_decap_8 FILLER_183_1596 ();
 sg13g2_decap_8 FILLER_183_1603 ();
 sg13g2_decap_8 FILLER_183_1610 ();
 sg13g2_decap_8 FILLER_183_1617 ();
 sg13g2_fill_1 FILLER_183_1624 ();
 sg13g2_decap_8 FILLER_184_0 ();
 sg13g2_decap_8 FILLER_184_7 ();
 sg13g2_decap_8 FILLER_184_14 ();
 sg13g2_decap_8 FILLER_184_21 ();
 sg13g2_decap_8 FILLER_184_28 ();
 sg13g2_decap_8 FILLER_184_35 ();
 sg13g2_decap_8 FILLER_184_42 ();
 sg13g2_decap_8 FILLER_184_49 ();
 sg13g2_decap_8 FILLER_184_56 ();
 sg13g2_decap_8 FILLER_184_63 ();
 sg13g2_decap_8 FILLER_184_70 ();
 sg13g2_decap_8 FILLER_184_77 ();
 sg13g2_decap_8 FILLER_184_84 ();
 sg13g2_decap_8 FILLER_184_91 ();
 sg13g2_decap_8 FILLER_184_98 ();
 sg13g2_decap_8 FILLER_184_105 ();
 sg13g2_decap_8 FILLER_184_112 ();
 sg13g2_decap_8 FILLER_184_119 ();
 sg13g2_decap_8 FILLER_184_126 ();
 sg13g2_decap_8 FILLER_184_133 ();
 sg13g2_decap_8 FILLER_184_140 ();
 sg13g2_decap_8 FILLER_184_147 ();
 sg13g2_decap_8 FILLER_184_154 ();
 sg13g2_decap_8 FILLER_184_161 ();
 sg13g2_decap_8 FILLER_184_168 ();
 sg13g2_decap_8 FILLER_184_175 ();
 sg13g2_decap_8 FILLER_184_182 ();
 sg13g2_decap_8 FILLER_184_189 ();
 sg13g2_decap_8 FILLER_184_196 ();
 sg13g2_decap_8 FILLER_184_203 ();
 sg13g2_decap_8 FILLER_184_210 ();
 sg13g2_decap_8 FILLER_184_217 ();
 sg13g2_decap_8 FILLER_184_224 ();
 sg13g2_decap_8 FILLER_184_231 ();
 sg13g2_decap_4 FILLER_184_238 ();
 sg13g2_decap_4 FILLER_184_301 ();
 sg13g2_fill_1 FILLER_184_309 ();
 sg13g2_fill_2 FILLER_184_320 ();
 sg13g2_fill_2 FILLER_184_365 ();
 sg13g2_decap_8 FILLER_184_376 ();
 sg13g2_fill_2 FILLER_184_383 ();
 sg13g2_fill_1 FILLER_184_385 ();
 sg13g2_fill_2 FILLER_184_392 ();
 sg13g2_fill_2 FILLER_184_442 ();
 sg13g2_decap_4 FILLER_184_449 ();
 sg13g2_fill_2 FILLER_184_505 ();
 sg13g2_fill_1 FILLER_184_516 ();
 sg13g2_fill_2 FILLER_184_521 ();
 sg13g2_fill_1 FILLER_184_523 ();
 sg13g2_fill_2 FILLER_184_529 ();
 sg13g2_fill_1 FILLER_184_531 ();
 sg13g2_fill_1 FILLER_184_540 ();
 sg13g2_decap_8 FILLER_184_545 ();
 sg13g2_fill_2 FILLER_184_552 ();
 sg13g2_decap_8 FILLER_184_558 ();
 sg13g2_decap_4 FILLER_184_565 ();
 sg13g2_fill_1 FILLER_184_603 ();
 sg13g2_decap_4 FILLER_184_607 ();
 sg13g2_fill_1 FILLER_184_611 ();
 sg13g2_fill_1 FILLER_184_616 ();
 sg13g2_fill_2 FILLER_184_622 ();
 sg13g2_fill_2 FILLER_184_663 ();
 sg13g2_fill_1 FILLER_184_665 ();
 sg13g2_fill_2 FILLER_184_709 ();
 sg13g2_fill_1 FILLER_184_711 ();
 sg13g2_fill_2 FILLER_184_746 ();
 sg13g2_decap_8 FILLER_184_778 ();
 sg13g2_decap_8 FILLER_184_785 ();
 sg13g2_fill_1 FILLER_184_792 ();
 sg13g2_decap_4 FILLER_184_797 ();
 sg13g2_fill_1 FILLER_184_801 ();
 sg13g2_decap_8 FILLER_184_806 ();
 sg13g2_decap_4 FILLER_184_813 ();
 sg13g2_fill_2 FILLER_184_817 ();
 sg13g2_decap_8 FILLER_184_823 ();
 sg13g2_decap_8 FILLER_184_830 ();
 sg13g2_fill_1 FILLER_184_837 ();
 sg13g2_decap_4 FILLER_184_844 ();
 sg13g2_fill_2 FILLER_184_848 ();
 sg13g2_fill_2 FILLER_184_880 ();
 sg13g2_decap_8 FILLER_184_894 ();
 sg13g2_decap_4 FILLER_184_901 ();
 sg13g2_decap_8 FILLER_184_909 ();
 sg13g2_decap_8 FILLER_184_916 ();
 sg13g2_decap_8 FILLER_184_923 ();
 sg13g2_decap_8 FILLER_184_930 ();
 sg13g2_decap_8 FILLER_184_937 ();
 sg13g2_decap_8 FILLER_184_944 ();
 sg13g2_decap_8 FILLER_184_951 ();
 sg13g2_decap_4 FILLER_184_958 ();
 sg13g2_fill_1 FILLER_184_962 ();
 sg13g2_decap_8 FILLER_184_975 ();
 sg13g2_fill_1 FILLER_184_982 ();
 sg13g2_decap_4 FILLER_184_1007 ();
 sg13g2_decap_8 FILLER_184_1015 ();
 sg13g2_decap_8 FILLER_184_1022 ();
 sg13g2_fill_2 FILLER_184_1029 ();
 sg13g2_decap_8 FILLER_184_1057 ();
 sg13g2_decap_4 FILLER_184_1064 ();
 sg13g2_fill_1 FILLER_184_1068 ();
 sg13g2_decap_8 FILLER_184_1081 ();
 sg13g2_fill_1 FILLER_184_1088 ();
 sg13g2_decap_4 FILLER_184_1101 ();
 sg13g2_decap_8 FILLER_184_1134 ();
 sg13g2_decap_8 FILLER_184_1141 ();
 sg13g2_decap_8 FILLER_184_1148 ();
 sg13g2_decap_8 FILLER_184_1155 ();
 sg13g2_decap_8 FILLER_184_1162 ();
 sg13g2_decap_8 FILLER_184_1169 ();
 sg13g2_decap_8 FILLER_184_1176 ();
 sg13g2_decap_8 FILLER_184_1183 ();
 sg13g2_decap_8 FILLER_184_1190 ();
 sg13g2_decap_8 FILLER_184_1197 ();
 sg13g2_decap_8 FILLER_184_1204 ();
 sg13g2_decap_8 FILLER_184_1211 ();
 sg13g2_decap_8 FILLER_184_1218 ();
 sg13g2_decap_8 FILLER_184_1225 ();
 sg13g2_decap_8 FILLER_184_1232 ();
 sg13g2_decap_8 FILLER_184_1239 ();
 sg13g2_decap_8 FILLER_184_1246 ();
 sg13g2_decap_8 FILLER_184_1253 ();
 sg13g2_decap_8 FILLER_184_1260 ();
 sg13g2_decap_8 FILLER_184_1267 ();
 sg13g2_decap_8 FILLER_184_1274 ();
 sg13g2_decap_8 FILLER_184_1281 ();
 sg13g2_decap_8 FILLER_184_1288 ();
 sg13g2_decap_8 FILLER_184_1295 ();
 sg13g2_decap_8 FILLER_184_1302 ();
 sg13g2_decap_8 FILLER_184_1309 ();
 sg13g2_decap_8 FILLER_184_1316 ();
 sg13g2_decap_8 FILLER_184_1323 ();
 sg13g2_decap_8 FILLER_184_1330 ();
 sg13g2_decap_8 FILLER_184_1337 ();
 sg13g2_decap_8 FILLER_184_1344 ();
 sg13g2_decap_8 FILLER_184_1351 ();
 sg13g2_decap_8 FILLER_184_1358 ();
 sg13g2_decap_8 FILLER_184_1365 ();
 sg13g2_decap_8 FILLER_184_1372 ();
 sg13g2_decap_8 FILLER_184_1379 ();
 sg13g2_decap_8 FILLER_184_1386 ();
 sg13g2_decap_8 FILLER_184_1393 ();
 sg13g2_decap_8 FILLER_184_1400 ();
 sg13g2_decap_8 FILLER_184_1407 ();
 sg13g2_decap_8 FILLER_184_1414 ();
 sg13g2_decap_8 FILLER_184_1421 ();
 sg13g2_decap_8 FILLER_184_1428 ();
 sg13g2_decap_8 FILLER_184_1435 ();
 sg13g2_decap_8 FILLER_184_1442 ();
 sg13g2_decap_8 FILLER_184_1449 ();
 sg13g2_decap_8 FILLER_184_1456 ();
 sg13g2_decap_8 FILLER_184_1463 ();
 sg13g2_decap_8 FILLER_184_1470 ();
 sg13g2_decap_8 FILLER_184_1477 ();
 sg13g2_decap_8 FILLER_184_1484 ();
 sg13g2_decap_8 FILLER_184_1491 ();
 sg13g2_decap_8 FILLER_184_1498 ();
 sg13g2_decap_8 FILLER_184_1505 ();
 sg13g2_decap_8 FILLER_184_1512 ();
 sg13g2_decap_8 FILLER_184_1519 ();
 sg13g2_decap_8 FILLER_184_1526 ();
 sg13g2_decap_8 FILLER_184_1533 ();
 sg13g2_decap_8 FILLER_184_1540 ();
 sg13g2_decap_8 FILLER_184_1547 ();
 sg13g2_decap_8 FILLER_184_1554 ();
 sg13g2_decap_8 FILLER_184_1561 ();
 sg13g2_decap_8 FILLER_184_1568 ();
 sg13g2_decap_8 FILLER_184_1575 ();
 sg13g2_decap_8 FILLER_184_1582 ();
 sg13g2_decap_8 FILLER_184_1589 ();
 sg13g2_decap_8 FILLER_184_1596 ();
 sg13g2_decap_8 FILLER_184_1603 ();
 sg13g2_decap_8 FILLER_184_1610 ();
 sg13g2_decap_8 FILLER_184_1617 ();
 sg13g2_fill_1 FILLER_184_1624 ();
 sg13g2_decap_8 FILLER_185_0 ();
 sg13g2_decap_8 FILLER_185_7 ();
 sg13g2_decap_8 FILLER_185_14 ();
 sg13g2_decap_8 FILLER_185_21 ();
 sg13g2_decap_8 FILLER_185_28 ();
 sg13g2_decap_8 FILLER_185_35 ();
 sg13g2_decap_8 FILLER_185_42 ();
 sg13g2_decap_8 FILLER_185_49 ();
 sg13g2_decap_8 FILLER_185_56 ();
 sg13g2_decap_8 FILLER_185_63 ();
 sg13g2_decap_8 FILLER_185_70 ();
 sg13g2_decap_8 FILLER_185_77 ();
 sg13g2_decap_8 FILLER_185_84 ();
 sg13g2_decap_8 FILLER_185_91 ();
 sg13g2_decap_8 FILLER_185_98 ();
 sg13g2_decap_8 FILLER_185_105 ();
 sg13g2_decap_8 FILLER_185_112 ();
 sg13g2_decap_8 FILLER_185_119 ();
 sg13g2_decap_8 FILLER_185_126 ();
 sg13g2_decap_8 FILLER_185_133 ();
 sg13g2_decap_8 FILLER_185_140 ();
 sg13g2_decap_8 FILLER_185_147 ();
 sg13g2_decap_8 FILLER_185_154 ();
 sg13g2_decap_8 FILLER_185_161 ();
 sg13g2_decap_8 FILLER_185_168 ();
 sg13g2_decap_8 FILLER_185_175 ();
 sg13g2_decap_8 FILLER_185_182 ();
 sg13g2_decap_8 FILLER_185_189 ();
 sg13g2_decap_8 FILLER_185_196 ();
 sg13g2_decap_8 FILLER_185_203 ();
 sg13g2_decap_8 FILLER_185_210 ();
 sg13g2_decap_8 FILLER_185_217 ();
 sg13g2_decap_8 FILLER_185_224 ();
 sg13g2_decap_8 FILLER_185_231 ();
 sg13g2_decap_8 FILLER_185_238 ();
 sg13g2_decap_8 FILLER_185_245 ();
 sg13g2_fill_1 FILLER_185_264 ();
 sg13g2_decap_8 FILLER_185_291 ();
 sg13g2_decap_4 FILLER_185_298 ();
 sg13g2_fill_1 FILLER_185_302 ();
 sg13g2_fill_2 FILLER_185_332 ();
 sg13g2_fill_1 FILLER_185_334 ();
 sg13g2_fill_2 FILLER_185_344 ();
 sg13g2_fill_1 FILLER_185_346 ();
 sg13g2_fill_2 FILLER_185_352 ();
 sg13g2_fill_1 FILLER_185_354 ();
 sg13g2_fill_2 FILLER_185_390 ();
 sg13g2_fill_2 FILLER_185_451 ();
 sg13g2_decap_8 FILLER_185_462 ();
 sg13g2_fill_2 FILLER_185_469 ();
 sg13g2_fill_2 FILLER_185_474 ();
 sg13g2_decap_8 FILLER_185_481 ();
 sg13g2_decap_8 FILLER_185_488 ();
 sg13g2_fill_2 FILLER_185_495 ();
 sg13g2_fill_2 FILLER_185_544 ();
 sg13g2_decap_8 FILLER_185_572 ();
 sg13g2_fill_2 FILLER_185_579 ();
 sg13g2_fill_1 FILLER_185_581 ();
 sg13g2_decap_4 FILLER_185_585 ();
 sg13g2_decap_8 FILLER_185_602 ();
 sg13g2_decap_8 FILLER_185_613 ();
 sg13g2_decap_4 FILLER_185_620 ();
 sg13g2_fill_2 FILLER_185_624 ();
 sg13g2_decap_8 FILLER_185_631 ();
 sg13g2_decap_8 FILLER_185_638 ();
 sg13g2_decap_4 FILLER_185_645 ();
 sg13g2_fill_1 FILLER_185_649 ();
 sg13g2_decap_8 FILLER_185_655 ();
 sg13g2_fill_1 FILLER_185_662 ();
 sg13g2_decap_8 FILLER_185_672 ();
 sg13g2_decap_8 FILLER_185_679 ();
 sg13g2_decap_4 FILLER_185_686 ();
 sg13g2_fill_2 FILLER_185_690 ();
 sg13g2_fill_2 FILLER_185_705 ();
 sg13g2_fill_1 FILLER_185_707 ();
 sg13g2_decap_8 FILLER_185_722 ();
 sg13g2_decap_8 FILLER_185_759 ();
 sg13g2_decap_8 FILLER_185_766 ();
 sg13g2_decap_8 FILLER_185_773 ();
 sg13g2_decap_8 FILLER_185_780 ();
 sg13g2_decap_8 FILLER_185_821 ();
 sg13g2_decap_8 FILLER_185_828 ();
 sg13g2_decap_8 FILLER_185_839 ();
 sg13g2_decap_8 FILLER_185_846 ();
 sg13g2_decap_8 FILLER_185_853 ();
 sg13g2_decap_8 FILLER_185_860 ();
 sg13g2_fill_2 FILLER_185_867 ();
 sg13g2_fill_1 FILLER_185_869 ();
 sg13g2_decap_4 FILLER_185_890 ();
 sg13g2_fill_2 FILLER_185_894 ();
 sg13g2_decap_8 FILLER_185_922 ();
 sg13g2_decap_8 FILLER_185_929 ();
 sg13g2_decap_8 FILLER_185_936 ();
 sg13g2_fill_2 FILLER_185_943 ();
 sg13g2_fill_1 FILLER_185_945 ();
 sg13g2_decap_8 FILLER_185_950 ();
 sg13g2_decap_4 FILLER_185_957 ();
 sg13g2_fill_1 FILLER_185_961 ();
 sg13g2_decap_4 FILLER_185_988 ();
 sg13g2_fill_2 FILLER_185_992 ();
 sg13g2_decap_8 FILLER_185_998 ();
 sg13g2_decap_8 FILLER_185_1005 ();
 sg13g2_decap_8 FILLER_185_1012 ();
 sg13g2_decap_8 FILLER_185_1019 ();
 sg13g2_decap_4 FILLER_185_1026 ();
 sg13g2_fill_2 FILLER_185_1030 ();
 sg13g2_fill_1 FILLER_185_1073 ();
 sg13g2_decap_8 FILLER_185_1078 ();
 sg13g2_decap_8 FILLER_185_1085 ();
 sg13g2_fill_2 FILLER_185_1092 ();
 sg13g2_decap_8 FILLER_185_1124 ();
 sg13g2_decap_8 FILLER_185_1131 ();
 sg13g2_decap_8 FILLER_185_1138 ();
 sg13g2_decap_8 FILLER_185_1145 ();
 sg13g2_decap_8 FILLER_185_1152 ();
 sg13g2_decap_8 FILLER_185_1159 ();
 sg13g2_decap_8 FILLER_185_1166 ();
 sg13g2_decap_8 FILLER_185_1173 ();
 sg13g2_decap_8 FILLER_185_1180 ();
 sg13g2_decap_8 FILLER_185_1187 ();
 sg13g2_decap_8 FILLER_185_1194 ();
 sg13g2_decap_8 FILLER_185_1201 ();
 sg13g2_decap_8 FILLER_185_1208 ();
 sg13g2_decap_8 FILLER_185_1215 ();
 sg13g2_decap_8 FILLER_185_1222 ();
 sg13g2_decap_8 FILLER_185_1229 ();
 sg13g2_decap_8 FILLER_185_1236 ();
 sg13g2_decap_8 FILLER_185_1243 ();
 sg13g2_decap_8 FILLER_185_1250 ();
 sg13g2_decap_8 FILLER_185_1257 ();
 sg13g2_decap_8 FILLER_185_1264 ();
 sg13g2_decap_8 FILLER_185_1271 ();
 sg13g2_decap_8 FILLER_185_1278 ();
 sg13g2_decap_8 FILLER_185_1285 ();
 sg13g2_decap_8 FILLER_185_1292 ();
 sg13g2_decap_8 FILLER_185_1299 ();
 sg13g2_decap_8 FILLER_185_1306 ();
 sg13g2_decap_8 FILLER_185_1313 ();
 sg13g2_decap_8 FILLER_185_1320 ();
 sg13g2_decap_8 FILLER_185_1327 ();
 sg13g2_decap_8 FILLER_185_1334 ();
 sg13g2_decap_8 FILLER_185_1341 ();
 sg13g2_decap_8 FILLER_185_1348 ();
 sg13g2_decap_8 FILLER_185_1355 ();
 sg13g2_decap_8 FILLER_185_1362 ();
 sg13g2_decap_8 FILLER_185_1369 ();
 sg13g2_decap_8 FILLER_185_1376 ();
 sg13g2_decap_8 FILLER_185_1383 ();
 sg13g2_decap_8 FILLER_185_1390 ();
 sg13g2_decap_8 FILLER_185_1397 ();
 sg13g2_decap_8 FILLER_185_1404 ();
 sg13g2_decap_8 FILLER_185_1411 ();
 sg13g2_decap_8 FILLER_185_1418 ();
 sg13g2_decap_8 FILLER_185_1425 ();
 sg13g2_decap_8 FILLER_185_1432 ();
 sg13g2_decap_8 FILLER_185_1439 ();
 sg13g2_decap_8 FILLER_185_1446 ();
 sg13g2_decap_8 FILLER_185_1453 ();
 sg13g2_decap_8 FILLER_185_1460 ();
 sg13g2_decap_8 FILLER_185_1467 ();
 sg13g2_decap_8 FILLER_185_1474 ();
 sg13g2_decap_8 FILLER_185_1481 ();
 sg13g2_decap_8 FILLER_185_1488 ();
 sg13g2_decap_8 FILLER_185_1495 ();
 sg13g2_decap_8 FILLER_185_1502 ();
 sg13g2_decap_8 FILLER_185_1509 ();
 sg13g2_decap_8 FILLER_185_1516 ();
 sg13g2_decap_8 FILLER_185_1523 ();
 sg13g2_decap_8 FILLER_185_1530 ();
 sg13g2_decap_8 FILLER_185_1537 ();
 sg13g2_decap_8 FILLER_185_1544 ();
 sg13g2_decap_8 FILLER_185_1551 ();
 sg13g2_decap_8 FILLER_185_1558 ();
 sg13g2_decap_8 FILLER_185_1565 ();
 sg13g2_decap_8 FILLER_185_1572 ();
 sg13g2_decap_8 FILLER_185_1579 ();
 sg13g2_decap_8 FILLER_185_1586 ();
 sg13g2_decap_8 FILLER_185_1593 ();
 sg13g2_decap_8 FILLER_185_1600 ();
 sg13g2_decap_8 FILLER_185_1607 ();
 sg13g2_decap_8 FILLER_185_1614 ();
 sg13g2_decap_4 FILLER_185_1621 ();
 sg13g2_decap_8 FILLER_186_0 ();
 sg13g2_decap_8 FILLER_186_7 ();
 sg13g2_decap_8 FILLER_186_14 ();
 sg13g2_decap_8 FILLER_186_21 ();
 sg13g2_decap_8 FILLER_186_28 ();
 sg13g2_decap_8 FILLER_186_35 ();
 sg13g2_decap_8 FILLER_186_42 ();
 sg13g2_decap_8 FILLER_186_49 ();
 sg13g2_decap_8 FILLER_186_56 ();
 sg13g2_decap_8 FILLER_186_63 ();
 sg13g2_decap_8 FILLER_186_70 ();
 sg13g2_decap_8 FILLER_186_77 ();
 sg13g2_decap_8 FILLER_186_84 ();
 sg13g2_decap_8 FILLER_186_91 ();
 sg13g2_decap_8 FILLER_186_98 ();
 sg13g2_decap_8 FILLER_186_105 ();
 sg13g2_decap_8 FILLER_186_112 ();
 sg13g2_decap_8 FILLER_186_119 ();
 sg13g2_decap_8 FILLER_186_126 ();
 sg13g2_decap_8 FILLER_186_133 ();
 sg13g2_decap_8 FILLER_186_140 ();
 sg13g2_decap_8 FILLER_186_147 ();
 sg13g2_decap_8 FILLER_186_154 ();
 sg13g2_decap_8 FILLER_186_161 ();
 sg13g2_decap_8 FILLER_186_168 ();
 sg13g2_decap_8 FILLER_186_175 ();
 sg13g2_decap_8 FILLER_186_182 ();
 sg13g2_decap_8 FILLER_186_189 ();
 sg13g2_decap_8 FILLER_186_196 ();
 sg13g2_decap_8 FILLER_186_203 ();
 sg13g2_decap_8 FILLER_186_210 ();
 sg13g2_decap_8 FILLER_186_217 ();
 sg13g2_decap_8 FILLER_186_224 ();
 sg13g2_decap_8 FILLER_186_231 ();
 sg13g2_decap_8 FILLER_186_238 ();
 sg13g2_decap_8 FILLER_186_245 ();
 sg13g2_decap_8 FILLER_186_257 ();
 sg13g2_decap_8 FILLER_186_264 ();
 sg13g2_decap_8 FILLER_186_271 ();
 sg13g2_fill_2 FILLER_186_278 ();
 sg13g2_fill_1 FILLER_186_280 ();
 sg13g2_decap_8 FILLER_186_313 ();
 sg13g2_decap_8 FILLER_186_320 ();
 sg13g2_fill_2 FILLER_186_327 ();
 sg13g2_fill_1 FILLER_186_333 ();
 sg13g2_decap_8 FILLER_186_389 ();
 sg13g2_decap_8 FILLER_186_396 ();
 sg13g2_fill_2 FILLER_186_403 ();
 sg13g2_fill_1 FILLER_186_405 ();
 sg13g2_fill_2 FILLER_186_414 ();
 sg13g2_decap_8 FILLER_186_450 ();
 sg13g2_fill_2 FILLER_186_457 ();
 sg13g2_fill_1 FILLER_186_459 ();
 sg13g2_decap_4 FILLER_186_469 ();
 sg13g2_fill_2 FILLER_186_473 ();
 sg13g2_decap_8 FILLER_186_479 ();
 sg13g2_fill_1 FILLER_186_486 ();
 sg13g2_decap_4 FILLER_186_492 ();
 sg13g2_decap_8 FILLER_186_522 ();
 sg13g2_decap_4 FILLER_186_529 ();
 sg13g2_fill_1 FILLER_186_533 ();
 sg13g2_fill_2 FILLER_186_539 ();
 sg13g2_fill_1 FILLER_186_541 ();
 sg13g2_decap_8 FILLER_186_550 ();
 sg13g2_decap_8 FILLER_186_557 ();
 sg13g2_decap_4 FILLER_186_564 ();
 sg13g2_fill_1 FILLER_186_568 ();
 sg13g2_decap_8 FILLER_186_633 ();
 sg13g2_fill_1 FILLER_186_640 ();
 sg13g2_decap_8 FILLER_186_645 ();
 sg13g2_decap_8 FILLER_186_652 ();
 sg13g2_decap_4 FILLER_186_659 ();
 sg13g2_fill_2 FILLER_186_663 ();
 sg13g2_fill_2 FILLER_186_669 ();
 sg13g2_fill_1 FILLER_186_671 ();
 sg13g2_decap_8 FILLER_186_717 ();
 sg13g2_decap_4 FILLER_186_724 ();
 sg13g2_decap_8 FILLER_186_757 ();
 sg13g2_decap_8 FILLER_186_764 ();
 sg13g2_decap_8 FILLER_186_771 ();
 sg13g2_decap_8 FILLER_186_778 ();
 sg13g2_decap_8 FILLER_186_785 ();
 sg13g2_decap_8 FILLER_186_792 ();
 sg13g2_fill_2 FILLER_186_799 ();
 sg13g2_fill_1 FILLER_186_801 ();
 sg13g2_fill_2 FILLER_186_810 ();
 sg13g2_fill_1 FILLER_186_812 ();
 sg13g2_decap_4 FILLER_186_818 ();
 sg13g2_fill_1 FILLER_186_822 ();
 sg13g2_decap_8 FILLER_186_853 ();
 sg13g2_decap_8 FILLER_186_860 ();
 sg13g2_decap_8 FILLER_186_867 ();
 sg13g2_decap_4 FILLER_186_874 ();
 sg13g2_decap_4 FILLER_186_887 ();
 sg13g2_fill_2 FILLER_186_891 ();
 sg13g2_fill_1 FILLER_186_897 ();
 sg13g2_decap_8 FILLER_186_931 ();
 sg13g2_fill_1 FILLER_186_938 ();
 sg13g2_fill_2 FILLER_186_965 ();
 sg13g2_fill_1 FILLER_186_967 ();
 sg13g2_fill_1 FILLER_186_972 ();
 sg13g2_fill_2 FILLER_186_977 ();
 sg13g2_decap_8 FILLER_186_1005 ();
 sg13g2_decap_8 FILLER_186_1012 ();
 sg13g2_decap_8 FILLER_186_1019 ();
 sg13g2_decap_8 FILLER_186_1026 ();
 sg13g2_decap_8 FILLER_186_1033 ();
 sg13g2_fill_1 FILLER_186_1066 ();
 sg13g2_decap_8 FILLER_186_1093 ();
 sg13g2_decap_8 FILLER_186_1100 ();
 sg13g2_decap_8 FILLER_186_1107 ();
 sg13g2_decap_8 FILLER_186_1114 ();
 sg13g2_decap_8 FILLER_186_1121 ();
 sg13g2_decap_8 FILLER_186_1128 ();
 sg13g2_decap_8 FILLER_186_1135 ();
 sg13g2_decap_8 FILLER_186_1142 ();
 sg13g2_decap_8 FILLER_186_1149 ();
 sg13g2_decap_8 FILLER_186_1156 ();
 sg13g2_decap_8 FILLER_186_1163 ();
 sg13g2_decap_8 FILLER_186_1170 ();
 sg13g2_decap_8 FILLER_186_1177 ();
 sg13g2_decap_8 FILLER_186_1184 ();
 sg13g2_decap_8 FILLER_186_1191 ();
 sg13g2_decap_8 FILLER_186_1198 ();
 sg13g2_decap_8 FILLER_186_1205 ();
 sg13g2_decap_8 FILLER_186_1212 ();
 sg13g2_decap_8 FILLER_186_1219 ();
 sg13g2_decap_8 FILLER_186_1226 ();
 sg13g2_decap_8 FILLER_186_1233 ();
 sg13g2_decap_8 FILLER_186_1240 ();
 sg13g2_decap_8 FILLER_186_1247 ();
 sg13g2_decap_8 FILLER_186_1254 ();
 sg13g2_decap_8 FILLER_186_1261 ();
 sg13g2_decap_8 FILLER_186_1268 ();
 sg13g2_decap_8 FILLER_186_1275 ();
 sg13g2_decap_8 FILLER_186_1282 ();
 sg13g2_decap_8 FILLER_186_1289 ();
 sg13g2_decap_8 FILLER_186_1296 ();
 sg13g2_decap_8 FILLER_186_1303 ();
 sg13g2_decap_8 FILLER_186_1310 ();
 sg13g2_decap_8 FILLER_186_1317 ();
 sg13g2_decap_8 FILLER_186_1324 ();
 sg13g2_decap_8 FILLER_186_1331 ();
 sg13g2_decap_8 FILLER_186_1338 ();
 sg13g2_decap_8 FILLER_186_1345 ();
 sg13g2_decap_8 FILLER_186_1352 ();
 sg13g2_decap_8 FILLER_186_1359 ();
 sg13g2_decap_8 FILLER_186_1366 ();
 sg13g2_decap_8 FILLER_186_1373 ();
 sg13g2_decap_8 FILLER_186_1380 ();
 sg13g2_decap_8 FILLER_186_1387 ();
 sg13g2_decap_8 FILLER_186_1394 ();
 sg13g2_decap_8 FILLER_186_1401 ();
 sg13g2_decap_8 FILLER_186_1408 ();
 sg13g2_decap_8 FILLER_186_1415 ();
 sg13g2_decap_8 FILLER_186_1422 ();
 sg13g2_decap_8 FILLER_186_1429 ();
 sg13g2_decap_8 FILLER_186_1436 ();
 sg13g2_decap_8 FILLER_186_1443 ();
 sg13g2_decap_8 FILLER_186_1450 ();
 sg13g2_decap_8 FILLER_186_1457 ();
 sg13g2_decap_8 FILLER_186_1464 ();
 sg13g2_decap_8 FILLER_186_1471 ();
 sg13g2_decap_8 FILLER_186_1478 ();
 sg13g2_decap_8 FILLER_186_1485 ();
 sg13g2_decap_8 FILLER_186_1492 ();
 sg13g2_decap_8 FILLER_186_1499 ();
 sg13g2_decap_8 FILLER_186_1506 ();
 sg13g2_decap_8 FILLER_186_1513 ();
 sg13g2_decap_8 FILLER_186_1520 ();
 sg13g2_decap_8 FILLER_186_1527 ();
 sg13g2_decap_8 FILLER_186_1534 ();
 sg13g2_decap_8 FILLER_186_1541 ();
 sg13g2_decap_8 FILLER_186_1548 ();
 sg13g2_decap_8 FILLER_186_1555 ();
 sg13g2_decap_8 FILLER_186_1562 ();
 sg13g2_decap_8 FILLER_186_1569 ();
 sg13g2_decap_8 FILLER_186_1576 ();
 sg13g2_decap_8 FILLER_186_1583 ();
 sg13g2_decap_8 FILLER_186_1590 ();
 sg13g2_decap_8 FILLER_186_1597 ();
 sg13g2_decap_8 FILLER_186_1604 ();
 sg13g2_decap_8 FILLER_186_1611 ();
 sg13g2_decap_8 FILLER_186_1618 ();
 sg13g2_decap_8 FILLER_187_0 ();
 sg13g2_decap_8 FILLER_187_7 ();
 sg13g2_decap_8 FILLER_187_14 ();
 sg13g2_decap_8 FILLER_187_21 ();
 sg13g2_decap_8 FILLER_187_28 ();
 sg13g2_decap_8 FILLER_187_35 ();
 sg13g2_decap_8 FILLER_187_42 ();
 sg13g2_decap_8 FILLER_187_49 ();
 sg13g2_decap_8 FILLER_187_56 ();
 sg13g2_decap_8 FILLER_187_63 ();
 sg13g2_decap_8 FILLER_187_70 ();
 sg13g2_decap_8 FILLER_187_77 ();
 sg13g2_decap_8 FILLER_187_84 ();
 sg13g2_decap_8 FILLER_187_91 ();
 sg13g2_decap_8 FILLER_187_98 ();
 sg13g2_decap_8 FILLER_187_105 ();
 sg13g2_decap_8 FILLER_187_112 ();
 sg13g2_decap_8 FILLER_187_119 ();
 sg13g2_decap_8 FILLER_187_126 ();
 sg13g2_decap_8 FILLER_187_133 ();
 sg13g2_decap_8 FILLER_187_140 ();
 sg13g2_decap_8 FILLER_187_147 ();
 sg13g2_decap_8 FILLER_187_154 ();
 sg13g2_decap_8 FILLER_187_161 ();
 sg13g2_decap_8 FILLER_187_168 ();
 sg13g2_decap_8 FILLER_187_175 ();
 sg13g2_decap_8 FILLER_187_182 ();
 sg13g2_decap_8 FILLER_187_189 ();
 sg13g2_decap_8 FILLER_187_196 ();
 sg13g2_decap_8 FILLER_187_203 ();
 sg13g2_decap_8 FILLER_187_210 ();
 sg13g2_decap_8 FILLER_187_217 ();
 sg13g2_decap_8 FILLER_187_224 ();
 sg13g2_decap_8 FILLER_187_231 ();
 sg13g2_decap_8 FILLER_187_238 ();
 sg13g2_decap_8 FILLER_187_245 ();
 sg13g2_decap_8 FILLER_187_252 ();
 sg13g2_decap_4 FILLER_187_259 ();
 sg13g2_fill_2 FILLER_187_263 ();
 sg13g2_decap_8 FILLER_187_269 ();
 sg13g2_fill_2 FILLER_187_276 ();
 sg13g2_fill_1 FILLER_187_278 ();
 sg13g2_decap_4 FILLER_187_328 ();
 sg13g2_decap_4 FILLER_187_336 ();
 sg13g2_fill_1 FILLER_187_340 ();
 sg13g2_decap_8 FILLER_187_345 ();
 sg13g2_decap_4 FILLER_187_352 ();
 sg13g2_decap_4 FILLER_187_386 ();
 sg13g2_fill_2 FILLER_187_390 ();
 sg13g2_fill_2 FILLER_187_396 ();
 sg13g2_fill_1 FILLER_187_424 ();
 sg13g2_decap_4 FILLER_187_451 ();
 sg13g2_decap_4 FILLER_187_494 ();
 sg13g2_fill_1 FILLER_187_498 ();
 sg13g2_fill_2 FILLER_187_516 ();
 sg13g2_fill_1 FILLER_187_518 ();
 sg13g2_fill_1 FILLER_187_529 ();
 sg13g2_fill_1 FILLER_187_534 ();
 sg13g2_fill_1 FILLER_187_541 ();
 sg13g2_fill_2 FILLER_187_552 ();
 sg13g2_fill_1 FILLER_187_558 ();
 sg13g2_fill_1 FILLER_187_576 ();
 sg13g2_fill_2 FILLER_187_582 ();
 sg13g2_fill_1 FILLER_187_584 ();
 sg13g2_decap_8 FILLER_187_594 ();
 sg13g2_decap_8 FILLER_187_601 ();
 sg13g2_decap_8 FILLER_187_608 ();
 sg13g2_decap_8 FILLER_187_615 ();
 sg13g2_decap_4 FILLER_187_622 ();
 sg13g2_fill_1 FILLER_187_660 ();
 sg13g2_decap_4 FILLER_187_713 ();
 sg13g2_decap_8 FILLER_187_747 ();
 sg13g2_decap_8 FILLER_187_754 ();
 sg13g2_decap_8 FILLER_187_761 ();
 sg13g2_decap_8 FILLER_187_768 ();
 sg13g2_decap_4 FILLER_187_775 ();
 sg13g2_decap_8 FILLER_187_819 ();
 sg13g2_decap_8 FILLER_187_826 ();
 sg13g2_fill_1 FILLER_187_841 ();
 sg13g2_decap_8 FILLER_187_856 ();
 sg13g2_fill_2 FILLER_187_863 ();
 sg13g2_fill_2 FILLER_187_874 ();
 sg13g2_fill_1 FILLER_187_910 ();
 sg13g2_decap_8 FILLER_187_937 ();
 sg13g2_fill_2 FILLER_187_948 ();
 sg13g2_decap_4 FILLER_187_958 ();
 sg13g2_decap_8 FILLER_187_995 ();
 sg13g2_decap_8 FILLER_187_1002 ();
 sg13g2_decap_8 FILLER_187_1009 ();
 sg13g2_decap_8 FILLER_187_1016 ();
 sg13g2_decap_8 FILLER_187_1023 ();
 sg13g2_decap_8 FILLER_187_1030 ();
 sg13g2_decap_8 FILLER_187_1037 ();
 sg13g2_fill_2 FILLER_187_1044 ();
 sg13g2_decap_8 FILLER_187_1050 ();
 sg13g2_decap_8 FILLER_187_1057 ();
 sg13g2_decap_8 FILLER_187_1064 ();
 sg13g2_decap_8 FILLER_187_1071 ();
 sg13g2_decap_8 FILLER_187_1078 ();
 sg13g2_decap_8 FILLER_187_1085 ();
 sg13g2_decap_8 FILLER_187_1092 ();
 sg13g2_decap_8 FILLER_187_1099 ();
 sg13g2_decap_8 FILLER_187_1106 ();
 sg13g2_decap_8 FILLER_187_1113 ();
 sg13g2_decap_8 FILLER_187_1120 ();
 sg13g2_decap_8 FILLER_187_1127 ();
 sg13g2_decap_8 FILLER_187_1134 ();
 sg13g2_decap_8 FILLER_187_1141 ();
 sg13g2_decap_8 FILLER_187_1148 ();
 sg13g2_decap_8 FILLER_187_1155 ();
 sg13g2_decap_8 FILLER_187_1162 ();
 sg13g2_decap_8 FILLER_187_1169 ();
 sg13g2_decap_8 FILLER_187_1176 ();
 sg13g2_decap_8 FILLER_187_1183 ();
 sg13g2_decap_8 FILLER_187_1190 ();
 sg13g2_decap_8 FILLER_187_1197 ();
 sg13g2_decap_8 FILLER_187_1204 ();
 sg13g2_decap_8 FILLER_187_1211 ();
 sg13g2_decap_8 FILLER_187_1218 ();
 sg13g2_decap_8 FILLER_187_1225 ();
 sg13g2_decap_8 FILLER_187_1232 ();
 sg13g2_decap_8 FILLER_187_1239 ();
 sg13g2_decap_8 FILLER_187_1246 ();
 sg13g2_decap_8 FILLER_187_1253 ();
 sg13g2_decap_8 FILLER_187_1260 ();
 sg13g2_decap_8 FILLER_187_1267 ();
 sg13g2_decap_8 FILLER_187_1274 ();
 sg13g2_decap_8 FILLER_187_1281 ();
 sg13g2_decap_8 FILLER_187_1288 ();
 sg13g2_decap_8 FILLER_187_1295 ();
 sg13g2_decap_8 FILLER_187_1302 ();
 sg13g2_decap_8 FILLER_187_1309 ();
 sg13g2_decap_8 FILLER_187_1316 ();
 sg13g2_decap_8 FILLER_187_1323 ();
 sg13g2_decap_8 FILLER_187_1330 ();
 sg13g2_decap_8 FILLER_187_1337 ();
 sg13g2_decap_8 FILLER_187_1344 ();
 sg13g2_decap_8 FILLER_187_1351 ();
 sg13g2_decap_8 FILLER_187_1358 ();
 sg13g2_decap_8 FILLER_187_1365 ();
 sg13g2_decap_8 FILLER_187_1372 ();
 sg13g2_decap_8 FILLER_187_1379 ();
 sg13g2_decap_8 FILLER_187_1386 ();
 sg13g2_decap_8 FILLER_187_1393 ();
 sg13g2_decap_8 FILLER_187_1400 ();
 sg13g2_decap_8 FILLER_187_1407 ();
 sg13g2_decap_8 FILLER_187_1414 ();
 sg13g2_decap_8 FILLER_187_1421 ();
 sg13g2_decap_8 FILLER_187_1428 ();
 sg13g2_decap_8 FILLER_187_1435 ();
 sg13g2_decap_8 FILLER_187_1442 ();
 sg13g2_decap_8 FILLER_187_1449 ();
 sg13g2_decap_8 FILLER_187_1456 ();
 sg13g2_decap_8 FILLER_187_1463 ();
 sg13g2_decap_8 FILLER_187_1470 ();
 sg13g2_decap_8 FILLER_187_1477 ();
 sg13g2_decap_8 FILLER_187_1484 ();
 sg13g2_decap_8 FILLER_187_1491 ();
 sg13g2_decap_8 FILLER_187_1498 ();
 sg13g2_decap_8 FILLER_187_1505 ();
 sg13g2_decap_8 FILLER_187_1512 ();
 sg13g2_decap_8 FILLER_187_1519 ();
 sg13g2_decap_8 FILLER_187_1526 ();
 sg13g2_decap_8 FILLER_187_1533 ();
 sg13g2_decap_8 FILLER_187_1540 ();
 sg13g2_decap_8 FILLER_187_1547 ();
 sg13g2_decap_8 FILLER_187_1554 ();
 sg13g2_decap_8 FILLER_187_1561 ();
 sg13g2_decap_8 FILLER_187_1568 ();
 sg13g2_decap_8 FILLER_187_1575 ();
 sg13g2_decap_8 FILLER_187_1582 ();
 sg13g2_decap_8 FILLER_187_1589 ();
 sg13g2_decap_8 FILLER_187_1596 ();
 sg13g2_decap_8 FILLER_187_1603 ();
 sg13g2_decap_8 FILLER_187_1610 ();
 sg13g2_decap_8 FILLER_187_1617 ();
 sg13g2_fill_1 FILLER_187_1624 ();
 sg13g2_decap_8 FILLER_188_0 ();
 sg13g2_decap_8 FILLER_188_7 ();
 sg13g2_decap_8 FILLER_188_14 ();
 sg13g2_decap_8 FILLER_188_21 ();
 sg13g2_decap_8 FILLER_188_28 ();
 sg13g2_decap_8 FILLER_188_35 ();
 sg13g2_decap_8 FILLER_188_42 ();
 sg13g2_decap_8 FILLER_188_49 ();
 sg13g2_decap_8 FILLER_188_56 ();
 sg13g2_decap_8 FILLER_188_63 ();
 sg13g2_decap_8 FILLER_188_70 ();
 sg13g2_decap_8 FILLER_188_77 ();
 sg13g2_decap_8 FILLER_188_84 ();
 sg13g2_decap_8 FILLER_188_91 ();
 sg13g2_decap_8 FILLER_188_98 ();
 sg13g2_decap_8 FILLER_188_105 ();
 sg13g2_decap_8 FILLER_188_112 ();
 sg13g2_decap_8 FILLER_188_119 ();
 sg13g2_decap_8 FILLER_188_126 ();
 sg13g2_decap_8 FILLER_188_133 ();
 sg13g2_decap_8 FILLER_188_140 ();
 sg13g2_decap_8 FILLER_188_147 ();
 sg13g2_decap_8 FILLER_188_154 ();
 sg13g2_decap_8 FILLER_188_161 ();
 sg13g2_decap_8 FILLER_188_168 ();
 sg13g2_decap_8 FILLER_188_175 ();
 sg13g2_decap_8 FILLER_188_182 ();
 sg13g2_decap_8 FILLER_188_189 ();
 sg13g2_decap_8 FILLER_188_196 ();
 sg13g2_decap_8 FILLER_188_203 ();
 sg13g2_decap_8 FILLER_188_210 ();
 sg13g2_decap_8 FILLER_188_217 ();
 sg13g2_decap_8 FILLER_188_224 ();
 sg13g2_decap_8 FILLER_188_231 ();
 sg13g2_decap_8 FILLER_188_238 ();
 sg13g2_decap_8 FILLER_188_245 ();
 sg13g2_decap_8 FILLER_188_252 ();
 sg13g2_fill_2 FILLER_188_259 ();
 sg13g2_decap_8 FILLER_188_277 ();
 sg13g2_fill_2 FILLER_188_284 ();
 sg13g2_fill_2 FILLER_188_319 ();
 sg13g2_fill_1 FILLER_188_321 ();
 sg13g2_decap_8 FILLER_188_377 ();
 sg13g2_fill_1 FILLER_188_384 ();
 sg13g2_decap_8 FILLER_188_440 ();
 sg13g2_decap_4 FILLER_188_447 ();
 sg13g2_fill_2 FILLER_188_451 ();
 sg13g2_decap_8 FILLER_188_458 ();
 sg13g2_decap_8 FILLER_188_465 ();
 sg13g2_decap_4 FILLER_188_472 ();
 sg13g2_fill_1 FILLER_188_483 ();
 sg13g2_fill_1 FILLER_188_612 ();
 sg13g2_decap_4 FILLER_188_652 ();
 sg13g2_fill_2 FILLER_188_656 ();
 sg13g2_decap_4 FILLER_188_671 ();
 sg13g2_fill_2 FILLER_188_675 ();
 sg13g2_decap_8 FILLER_188_683 ();
 sg13g2_decap_8 FILLER_188_690 ();
 sg13g2_decap_8 FILLER_188_697 ();
 sg13g2_decap_8 FILLER_188_704 ();
 sg13g2_decap_8 FILLER_188_711 ();
 sg13g2_decap_8 FILLER_188_718 ();
 sg13g2_decap_4 FILLER_188_725 ();
 sg13g2_fill_1 FILLER_188_729 ();
 sg13g2_decap_8 FILLER_188_737 ();
 sg13g2_decap_8 FILLER_188_744 ();
 sg13g2_decap_8 FILLER_188_751 ();
 sg13g2_decap_8 FILLER_188_758 ();
 sg13g2_decap_8 FILLER_188_765 ();
 sg13g2_decap_4 FILLER_188_772 ();
 sg13g2_fill_1 FILLER_188_806 ();
 sg13g2_decap_8 FILLER_188_826 ();
 sg13g2_decap_8 FILLER_188_833 ();
 sg13g2_decap_4 FILLER_188_840 ();
 sg13g2_decap_4 FILLER_188_869 ();
 sg13g2_fill_1 FILLER_188_873 ();
 sg13g2_fill_2 FILLER_188_880 ();
 sg13g2_fill_1 FILLER_188_882 ();
 sg13g2_decap_8 FILLER_188_887 ();
 sg13g2_decap_8 FILLER_188_894 ();
 sg13g2_decap_8 FILLER_188_901 ();
 sg13g2_decap_4 FILLER_188_908 ();
 sg13g2_decap_4 FILLER_188_931 ();
 sg13g2_fill_1 FILLER_188_935 ();
 sg13g2_fill_2 FILLER_188_939 ();
 sg13g2_fill_1 FILLER_188_941 ();
 sg13g2_fill_2 FILLER_188_954 ();
 sg13g2_decap_8 FILLER_188_990 ();
 sg13g2_decap_8 FILLER_188_997 ();
 sg13g2_decap_8 FILLER_188_1004 ();
 sg13g2_decap_8 FILLER_188_1011 ();
 sg13g2_decap_8 FILLER_188_1018 ();
 sg13g2_decap_8 FILLER_188_1025 ();
 sg13g2_decap_8 FILLER_188_1032 ();
 sg13g2_decap_8 FILLER_188_1039 ();
 sg13g2_decap_8 FILLER_188_1046 ();
 sg13g2_decap_8 FILLER_188_1053 ();
 sg13g2_decap_8 FILLER_188_1060 ();
 sg13g2_decap_8 FILLER_188_1067 ();
 sg13g2_decap_8 FILLER_188_1074 ();
 sg13g2_decap_8 FILLER_188_1081 ();
 sg13g2_decap_8 FILLER_188_1088 ();
 sg13g2_decap_8 FILLER_188_1095 ();
 sg13g2_decap_8 FILLER_188_1102 ();
 sg13g2_decap_8 FILLER_188_1109 ();
 sg13g2_decap_8 FILLER_188_1116 ();
 sg13g2_decap_8 FILLER_188_1123 ();
 sg13g2_decap_8 FILLER_188_1130 ();
 sg13g2_decap_8 FILLER_188_1137 ();
 sg13g2_decap_8 FILLER_188_1144 ();
 sg13g2_decap_8 FILLER_188_1151 ();
 sg13g2_decap_8 FILLER_188_1158 ();
 sg13g2_decap_8 FILLER_188_1165 ();
 sg13g2_decap_8 FILLER_188_1172 ();
 sg13g2_decap_8 FILLER_188_1179 ();
 sg13g2_decap_8 FILLER_188_1186 ();
 sg13g2_decap_8 FILLER_188_1193 ();
 sg13g2_decap_8 FILLER_188_1200 ();
 sg13g2_decap_8 FILLER_188_1207 ();
 sg13g2_decap_8 FILLER_188_1214 ();
 sg13g2_decap_8 FILLER_188_1221 ();
 sg13g2_decap_8 FILLER_188_1228 ();
 sg13g2_decap_8 FILLER_188_1235 ();
 sg13g2_decap_8 FILLER_188_1242 ();
 sg13g2_decap_8 FILLER_188_1249 ();
 sg13g2_decap_8 FILLER_188_1256 ();
 sg13g2_decap_8 FILLER_188_1263 ();
 sg13g2_decap_8 FILLER_188_1270 ();
 sg13g2_decap_8 FILLER_188_1277 ();
 sg13g2_decap_8 FILLER_188_1284 ();
 sg13g2_decap_8 FILLER_188_1291 ();
 sg13g2_decap_8 FILLER_188_1298 ();
 sg13g2_decap_8 FILLER_188_1305 ();
 sg13g2_decap_8 FILLER_188_1312 ();
 sg13g2_decap_8 FILLER_188_1319 ();
 sg13g2_decap_8 FILLER_188_1326 ();
 sg13g2_decap_8 FILLER_188_1333 ();
 sg13g2_decap_8 FILLER_188_1340 ();
 sg13g2_decap_8 FILLER_188_1347 ();
 sg13g2_decap_8 FILLER_188_1354 ();
 sg13g2_decap_8 FILLER_188_1361 ();
 sg13g2_decap_8 FILLER_188_1368 ();
 sg13g2_decap_8 FILLER_188_1375 ();
 sg13g2_decap_8 FILLER_188_1382 ();
 sg13g2_decap_8 FILLER_188_1389 ();
 sg13g2_decap_8 FILLER_188_1396 ();
 sg13g2_decap_8 FILLER_188_1403 ();
 sg13g2_decap_8 FILLER_188_1410 ();
 sg13g2_decap_8 FILLER_188_1417 ();
 sg13g2_decap_8 FILLER_188_1424 ();
 sg13g2_decap_8 FILLER_188_1431 ();
 sg13g2_decap_8 FILLER_188_1438 ();
 sg13g2_decap_8 FILLER_188_1445 ();
 sg13g2_decap_8 FILLER_188_1452 ();
 sg13g2_decap_8 FILLER_188_1459 ();
 sg13g2_decap_8 FILLER_188_1466 ();
 sg13g2_decap_8 FILLER_188_1473 ();
 sg13g2_decap_8 FILLER_188_1480 ();
 sg13g2_decap_8 FILLER_188_1487 ();
 sg13g2_decap_8 FILLER_188_1494 ();
 sg13g2_decap_8 FILLER_188_1501 ();
 sg13g2_decap_8 FILLER_188_1508 ();
 sg13g2_decap_8 FILLER_188_1515 ();
 sg13g2_decap_8 FILLER_188_1522 ();
 sg13g2_decap_8 FILLER_188_1529 ();
 sg13g2_decap_8 FILLER_188_1536 ();
 sg13g2_decap_8 FILLER_188_1543 ();
 sg13g2_decap_8 FILLER_188_1550 ();
 sg13g2_decap_8 FILLER_188_1557 ();
 sg13g2_decap_8 FILLER_188_1564 ();
 sg13g2_decap_8 FILLER_188_1571 ();
 sg13g2_decap_8 FILLER_188_1578 ();
 sg13g2_decap_8 FILLER_188_1585 ();
 sg13g2_decap_8 FILLER_188_1592 ();
 sg13g2_decap_8 FILLER_188_1599 ();
 sg13g2_decap_8 FILLER_188_1606 ();
 sg13g2_decap_8 FILLER_188_1613 ();
 sg13g2_decap_4 FILLER_188_1620 ();
 sg13g2_fill_1 FILLER_188_1624 ();
 sg13g2_decap_8 FILLER_189_0 ();
 sg13g2_decap_8 FILLER_189_7 ();
 sg13g2_decap_8 FILLER_189_14 ();
 sg13g2_decap_8 FILLER_189_21 ();
 sg13g2_decap_8 FILLER_189_28 ();
 sg13g2_decap_8 FILLER_189_35 ();
 sg13g2_decap_8 FILLER_189_42 ();
 sg13g2_decap_8 FILLER_189_49 ();
 sg13g2_decap_8 FILLER_189_56 ();
 sg13g2_decap_8 FILLER_189_63 ();
 sg13g2_decap_8 FILLER_189_70 ();
 sg13g2_decap_8 FILLER_189_77 ();
 sg13g2_decap_8 FILLER_189_84 ();
 sg13g2_decap_8 FILLER_189_91 ();
 sg13g2_decap_8 FILLER_189_98 ();
 sg13g2_decap_8 FILLER_189_105 ();
 sg13g2_decap_8 FILLER_189_112 ();
 sg13g2_decap_8 FILLER_189_119 ();
 sg13g2_decap_8 FILLER_189_126 ();
 sg13g2_decap_8 FILLER_189_133 ();
 sg13g2_decap_8 FILLER_189_140 ();
 sg13g2_decap_8 FILLER_189_147 ();
 sg13g2_decap_8 FILLER_189_154 ();
 sg13g2_decap_8 FILLER_189_161 ();
 sg13g2_decap_8 FILLER_189_168 ();
 sg13g2_decap_8 FILLER_189_175 ();
 sg13g2_decap_8 FILLER_189_182 ();
 sg13g2_decap_8 FILLER_189_189 ();
 sg13g2_decap_8 FILLER_189_196 ();
 sg13g2_decap_8 FILLER_189_203 ();
 sg13g2_decap_8 FILLER_189_210 ();
 sg13g2_decap_8 FILLER_189_217 ();
 sg13g2_decap_8 FILLER_189_224 ();
 sg13g2_decap_8 FILLER_189_231 ();
 sg13g2_decap_8 FILLER_189_238 ();
 sg13g2_decap_8 FILLER_189_245 ();
 sg13g2_decap_8 FILLER_189_252 ();
 sg13g2_decap_4 FILLER_189_259 ();
 sg13g2_fill_1 FILLER_189_263 ();
 sg13g2_decap_4 FILLER_189_316 ();
 sg13g2_fill_2 FILLER_189_320 ();
 sg13g2_decap_8 FILLER_189_325 ();
 sg13g2_decap_8 FILLER_189_332 ();
 sg13g2_decap_4 FILLER_189_339 ();
 sg13g2_fill_2 FILLER_189_343 ();
 sg13g2_decap_4 FILLER_189_355 ();
 sg13g2_decap_4 FILLER_189_363 ();
 sg13g2_decap_8 FILLER_189_371 ();
 sg13g2_decap_8 FILLER_189_378 ();
 sg13g2_decap_8 FILLER_189_385 ();
 sg13g2_decap_4 FILLER_189_392 ();
 sg13g2_decap_8 FILLER_189_399 ();
 sg13g2_fill_2 FILLER_189_406 ();
 sg13g2_decap_8 FILLER_189_434 ();
 sg13g2_fill_2 FILLER_189_441 ();
 sg13g2_fill_1 FILLER_189_443 ();
 sg13g2_fill_1 FILLER_189_462 ();
 sg13g2_fill_1 FILLER_189_543 ();
 sg13g2_fill_1 FILLER_189_570 ();
 sg13g2_decap_4 FILLER_189_607 ();
 sg13g2_fill_1 FILLER_189_615 ();
 sg13g2_decap_8 FILLER_189_642 ();
 sg13g2_fill_2 FILLER_189_649 ();
 sg13g2_fill_1 FILLER_189_651 ();
 sg13g2_fill_1 FILLER_189_690 ();
 sg13g2_fill_2 FILLER_189_695 ();
 sg13g2_fill_1 FILLER_189_697 ();
 sg13g2_fill_1 FILLER_189_717 ();
 sg13g2_fill_2 FILLER_189_722 ();
 sg13g2_decap_8 FILLER_189_750 ();
 sg13g2_decap_8 FILLER_189_757 ();
 sg13g2_decap_8 FILLER_189_764 ();
 sg13g2_decap_4 FILLER_189_771 ();
 sg13g2_fill_1 FILLER_189_775 ();
 sg13g2_fill_1 FILLER_189_805 ();
 sg13g2_fill_1 FILLER_189_814 ();
 sg13g2_fill_1 FILLER_189_823 ();
 sg13g2_fill_1 FILLER_189_828 ();
 sg13g2_decap_4 FILLER_189_833 ();
 sg13g2_fill_2 FILLER_189_837 ();
 sg13g2_decap_8 FILLER_189_844 ();
 sg13g2_decap_8 FILLER_189_851 ();
 sg13g2_fill_2 FILLER_189_858 ();
 sg13g2_decap_8 FILLER_189_866 ();
 sg13g2_decap_8 FILLER_189_873 ();
 sg13g2_decap_8 FILLER_189_880 ();
 sg13g2_fill_2 FILLER_189_887 ();
 sg13g2_fill_1 FILLER_189_889 ();
 sg13g2_fill_2 FILLER_189_895 ();
 sg13g2_fill_1 FILLER_189_897 ();
 sg13g2_decap_8 FILLER_189_902 ();
 sg13g2_decap_8 FILLER_189_909 ();
 sg13g2_fill_2 FILLER_189_916 ();
 sg13g2_decap_8 FILLER_189_925 ();
 sg13g2_decap_8 FILLER_189_932 ();
 sg13g2_decap_8 FILLER_189_939 ();
 sg13g2_decap_8 FILLER_189_946 ();
 sg13g2_decap_4 FILLER_189_953 ();
 sg13g2_decap_8 FILLER_189_962 ();
 sg13g2_decap_8 FILLER_189_969 ();
 sg13g2_decap_8 FILLER_189_976 ();
 sg13g2_decap_8 FILLER_189_983 ();
 sg13g2_decap_8 FILLER_189_990 ();
 sg13g2_decap_8 FILLER_189_997 ();
 sg13g2_decap_8 FILLER_189_1004 ();
 sg13g2_decap_8 FILLER_189_1011 ();
 sg13g2_decap_8 FILLER_189_1018 ();
 sg13g2_decap_8 FILLER_189_1025 ();
 sg13g2_decap_8 FILLER_189_1032 ();
 sg13g2_decap_8 FILLER_189_1039 ();
 sg13g2_decap_8 FILLER_189_1046 ();
 sg13g2_decap_8 FILLER_189_1053 ();
 sg13g2_decap_8 FILLER_189_1060 ();
 sg13g2_decap_8 FILLER_189_1067 ();
 sg13g2_decap_8 FILLER_189_1074 ();
 sg13g2_decap_8 FILLER_189_1081 ();
 sg13g2_decap_8 FILLER_189_1088 ();
 sg13g2_decap_8 FILLER_189_1095 ();
 sg13g2_decap_8 FILLER_189_1102 ();
 sg13g2_decap_8 FILLER_189_1109 ();
 sg13g2_decap_8 FILLER_189_1116 ();
 sg13g2_decap_8 FILLER_189_1123 ();
 sg13g2_decap_8 FILLER_189_1130 ();
 sg13g2_decap_8 FILLER_189_1137 ();
 sg13g2_decap_8 FILLER_189_1144 ();
 sg13g2_decap_8 FILLER_189_1151 ();
 sg13g2_decap_8 FILLER_189_1158 ();
 sg13g2_decap_8 FILLER_189_1165 ();
 sg13g2_decap_8 FILLER_189_1172 ();
 sg13g2_decap_8 FILLER_189_1179 ();
 sg13g2_decap_8 FILLER_189_1186 ();
 sg13g2_decap_8 FILLER_189_1193 ();
 sg13g2_decap_8 FILLER_189_1200 ();
 sg13g2_decap_8 FILLER_189_1207 ();
 sg13g2_decap_8 FILLER_189_1214 ();
 sg13g2_decap_8 FILLER_189_1221 ();
 sg13g2_decap_8 FILLER_189_1228 ();
 sg13g2_decap_8 FILLER_189_1235 ();
 sg13g2_decap_8 FILLER_189_1242 ();
 sg13g2_decap_8 FILLER_189_1249 ();
 sg13g2_decap_8 FILLER_189_1256 ();
 sg13g2_decap_8 FILLER_189_1263 ();
 sg13g2_decap_8 FILLER_189_1270 ();
 sg13g2_decap_8 FILLER_189_1277 ();
 sg13g2_decap_8 FILLER_189_1284 ();
 sg13g2_decap_8 FILLER_189_1291 ();
 sg13g2_decap_8 FILLER_189_1298 ();
 sg13g2_decap_8 FILLER_189_1305 ();
 sg13g2_decap_8 FILLER_189_1312 ();
 sg13g2_decap_8 FILLER_189_1319 ();
 sg13g2_decap_8 FILLER_189_1326 ();
 sg13g2_decap_8 FILLER_189_1333 ();
 sg13g2_decap_8 FILLER_189_1340 ();
 sg13g2_decap_8 FILLER_189_1347 ();
 sg13g2_decap_8 FILLER_189_1354 ();
 sg13g2_decap_8 FILLER_189_1361 ();
 sg13g2_decap_8 FILLER_189_1368 ();
 sg13g2_decap_8 FILLER_189_1375 ();
 sg13g2_decap_8 FILLER_189_1382 ();
 sg13g2_decap_8 FILLER_189_1389 ();
 sg13g2_decap_8 FILLER_189_1396 ();
 sg13g2_decap_8 FILLER_189_1403 ();
 sg13g2_decap_8 FILLER_189_1410 ();
 sg13g2_decap_8 FILLER_189_1417 ();
 sg13g2_decap_8 FILLER_189_1424 ();
 sg13g2_decap_8 FILLER_189_1431 ();
 sg13g2_decap_8 FILLER_189_1438 ();
 sg13g2_decap_8 FILLER_189_1445 ();
 sg13g2_decap_8 FILLER_189_1452 ();
 sg13g2_decap_8 FILLER_189_1459 ();
 sg13g2_decap_8 FILLER_189_1466 ();
 sg13g2_decap_8 FILLER_189_1473 ();
 sg13g2_decap_8 FILLER_189_1480 ();
 sg13g2_decap_8 FILLER_189_1487 ();
 sg13g2_decap_8 FILLER_189_1494 ();
 sg13g2_decap_8 FILLER_189_1501 ();
 sg13g2_decap_8 FILLER_189_1508 ();
 sg13g2_decap_8 FILLER_189_1515 ();
 sg13g2_decap_8 FILLER_189_1522 ();
 sg13g2_decap_8 FILLER_189_1529 ();
 sg13g2_decap_8 FILLER_189_1536 ();
 sg13g2_decap_8 FILLER_189_1543 ();
 sg13g2_decap_8 FILLER_189_1550 ();
 sg13g2_decap_8 FILLER_189_1557 ();
 sg13g2_decap_8 FILLER_189_1564 ();
 sg13g2_decap_8 FILLER_189_1571 ();
 sg13g2_decap_8 FILLER_189_1578 ();
 sg13g2_decap_8 FILLER_189_1585 ();
 sg13g2_decap_8 FILLER_189_1592 ();
 sg13g2_decap_8 FILLER_189_1599 ();
 sg13g2_decap_8 FILLER_189_1606 ();
 sg13g2_decap_8 FILLER_189_1613 ();
 sg13g2_decap_4 FILLER_189_1620 ();
 sg13g2_fill_1 FILLER_189_1624 ();
 sg13g2_decap_8 FILLER_190_0 ();
 sg13g2_decap_8 FILLER_190_7 ();
 sg13g2_decap_8 FILLER_190_14 ();
 sg13g2_decap_8 FILLER_190_21 ();
 sg13g2_decap_8 FILLER_190_28 ();
 sg13g2_decap_8 FILLER_190_35 ();
 sg13g2_decap_8 FILLER_190_42 ();
 sg13g2_decap_8 FILLER_190_49 ();
 sg13g2_decap_8 FILLER_190_56 ();
 sg13g2_decap_8 FILLER_190_63 ();
 sg13g2_decap_8 FILLER_190_70 ();
 sg13g2_decap_8 FILLER_190_77 ();
 sg13g2_decap_8 FILLER_190_84 ();
 sg13g2_decap_8 FILLER_190_91 ();
 sg13g2_decap_8 FILLER_190_98 ();
 sg13g2_decap_8 FILLER_190_105 ();
 sg13g2_decap_8 FILLER_190_112 ();
 sg13g2_decap_8 FILLER_190_119 ();
 sg13g2_decap_8 FILLER_190_126 ();
 sg13g2_decap_8 FILLER_190_133 ();
 sg13g2_decap_8 FILLER_190_140 ();
 sg13g2_decap_8 FILLER_190_147 ();
 sg13g2_decap_8 FILLER_190_154 ();
 sg13g2_decap_8 FILLER_190_161 ();
 sg13g2_decap_8 FILLER_190_168 ();
 sg13g2_decap_8 FILLER_190_175 ();
 sg13g2_decap_8 FILLER_190_182 ();
 sg13g2_decap_8 FILLER_190_189 ();
 sg13g2_decap_8 FILLER_190_196 ();
 sg13g2_decap_8 FILLER_190_203 ();
 sg13g2_decap_8 FILLER_190_210 ();
 sg13g2_decap_8 FILLER_190_217 ();
 sg13g2_decap_8 FILLER_190_224 ();
 sg13g2_decap_8 FILLER_190_231 ();
 sg13g2_decap_8 FILLER_190_238 ();
 sg13g2_decap_8 FILLER_190_245 ();
 sg13g2_decap_8 FILLER_190_252 ();
 sg13g2_decap_8 FILLER_190_259 ();
 sg13g2_decap_8 FILLER_190_266 ();
 sg13g2_decap_8 FILLER_190_273 ();
 sg13g2_decap_8 FILLER_190_280 ();
 sg13g2_decap_8 FILLER_190_287 ();
 sg13g2_decap_8 FILLER_190_294 ();
 sg13g2_decap_8 FILLER_190_301 ();
 sg13g2_decap_8 FILLER_190_308 ();
 sg13g2_decap_4 FILLER_190_315 ();
 sg13g2_fill_2 FILLER_190_319 ();
 sg13g2_fill_2 FILLER_190_330 ();
 sg13g2_fill_1 FILLER_190_332 ();
 sg13g2_decap_8 FILLER_190_336 ();
 sg13g2_fill_2 FILLER_190_343 ();
 sg13g2_fill_1 FILLER_190_350 ();
 sg13g2_fill_1 FILLER_190_356 ();
 sg13g2_fill_1 FILLER_190_362 ();
 sg13g2_fill_1 FILLER_190_367 ();
 sg13g2_fill_2 FILLER_190_392 ();
 sg13g2_decap_4 FILLER_190_399 ();
 sg13g2_decap_8 FILLER_190_408 ();
 sg13g2_decap_8 FILLER_190_419 ();
 sg13g2_decap_4 FILLER_190_426 ();
 sg13g2_fill_1 FILLER_190_430 ();
 sg13g2_fill_2 FILLER_190_435 ();
 sg13g2_decap_8 FILLER_190_445 ();
 sg13g2_fill_1 FILLER_190_452 ();
 sg13g2_decap_4 FILLER_190_457 ();
 sg13g2_fill_2 FILLER_190_500 ();
 sg13g2_decap_8 FILLER_190_532 ();
 sg13g2_fill_1 FILLER_190_539 ();
 sg13g2_decap_8 FILLER_190_609 ();
 sg13g2_decap_8 FILLER_190_616 ();
 sg13g2_decap_8 FILLER_190_629 ();
 sg13g2_decap_8 FILLER_190_636 ();
 sg13g2_fill_2 FILLER_190_643 ();
 sg13g2_fill_1 FILLER_190_659 ();
 sg13g2_fill_2 FILLER_190_692 ();
 sg13g2_decap_4 FILLER_190_703 ();
 sg13g2_decap_8 FILLER_190_751 ();
 sg13g2_decap_8 FILLER_190_758 ();
 sg13g2_decap_8 FILLER_190_765 ();
 sg13g2_decap_8 FILLER_190_772 ();
 sg13g2_decap_4 FILLER_190_779 ();
 sg13g2_fill_2 FILLER_190_783 ();
 sg13g2_decap_8 FILLER_190_814 ();
 sg13g2_decap_8 FILLER_190_847 ();
 sg13g2_decap_4 FILLER_190_866 ();
 sg13g2_fill_1 FILLER_190_870 ();
 sg13g2_decap_8 FILLER_190_875 ();
 sg13g2_decap_8 FILLER_190_882 ();
 sg13g2_fill_2 FILLER_190_889 ();
 sg13g2_decap_8 FILLER_190_925 ();
 sg13g2_fill_1 FILLER_190_932 ();
 sg13g2_fill_2 FILLER_190_941 ();
 sg13g2_fill_1 FILLER_190_943 ();
 sg13g2_decap_4 FILLER_190_952 ();
 sg13g2_decap_8 FILLER_190_968 ();
 sg13g2_decap_8 FILLER_190_975 ();
 sg13g2_decap_8 FILLER_190_982 ();
 sg13g2_decap_8 FILLER_190_989 ();
 sg13g2_decap_8 FILLER_190_996 ();
 sg13g2_decap_8 FILLER_190_1003 ();
 sg13g2_decap_8 FILLER_190_1010 ();
 sg13g2_decap_8 FILLER_190_1017 ();
 sg13g2_decap_8 FILLER_190_1024 ();
 sg13g2_decap_8 FILLER_190_1031 ();
 sg13g2_decap_8 FILLER_190_1038 ();
 sg13g2_decap_8 FILLER_190_1045 ();
 sg13g2_decap_8 FILLER_190_1052 ();
 sg13g2_decap_8 FILLER_190_1059 ();
 sg13g2_decap_8 FILLER_190_1066 ();
 sg13g2_decap_8 FILLER_190_1073 ();
 sg13g2_decap_8 FILLER_190_1080 ();
 sg13g2_decap_8 FILLER_190_1087 ();
 sg13g2_decap_8 FILLER_190_1094 ();
 sg13g2_decap_8 FILLER_190_1101 ();
 sg13g2_decap_8 FILLER_190_1108 ();
 sg13g2_decap_8 FILLER_190_1115 ();
 sg13g2_decap_8 FILLER_190_1122 ();
 sg13g2_decap_8 FILLER_190_1129 ();
 sg13g2_decap_8 FILLER_190_1136 ();
 sg13g2_decap_8 FILLER_190_1143 ();
 sg13g2_decap_8 FILLER_190_1150 ();
 sg13g2_decap_8 FILLER_190_1157 ();
 sg13g2_decap_8 FILLER_190_1164 ();
 sg13g2_decap_8 FILLER_190_1171 ();
 sg13g2_decap_8 FILLER_190_1178 ();
 sg13g2_decap_8 FILLER_190_1185 ();
 sg13g2_decap_8 FILLER_190_1192 ();
 sg13g2_decap_8 FILLER_190_1199 ();
 sg13g2_decap_8 FILLER_190_1206 ();
 sg13g2_decap_8 FILLER_190_1213 ();
 sg13g2_decap_8 FILLER_190_1220 ();
 sg13g2_decap_8 FILLER_190_1227 ();
 sg13g2_decap_8 FILLER_190_1234 ();
 sg13g2_decap_8 FILLER_190_1241 ();
 sg13g2_decap_8 FILLER_190_1248 ();
 sg13g2_decap_8 FILLER_190_1255 ();
 sg13g2_decap_8 FILLER_190_1262 ();
 sg13g2_decap_8 FILLER_190_1269 ();
 sg13g2_decap_8 FILLER_190_1276 ();
 sg13g2_decap_8 FILLER_190_1283 ();
 sg13g2_decap_8 FILLER_190_1290 ();
 sg13g2_decap_8 FILLER_190_1297 ();
 sg13g2_decap_8 FILLER_190_1304 ();
 sg13g2_decap_8 FILLER_190_1311 ();
 sg13g2_decap_8 FILLER_190_1318 ();
 sg13g2_decap_8 FILLER_190_1325 ();
 sg13g2_decap_8 FILLER_190_1332 ();
 sg13g2_decap_8 FILLER_190_1339 ();
 sg13g2_decap_8 FILLER_190_1346 ();
 sg13g2_decap_8 FILLER_190_1353 ();
 sg13g2_decap_8 FILLER_190_1360 ();
 sg13g2_decap_8 FILLER_190_1367 ();
 sg13g2_decap_8 FILLER_190_1374 ();
 sg13g2_decap_8 FILLER_190_1381 ();
 sg13g2_decap_8 FILLER_190_1388 ();
 sg13g2_decap_8 FILLER_190_1395 ();
 sg13g2_decap_8 FILLER_190_1402 ();
 sg13g2_decap_8 FILLER_190_1409 ();
 sg13g2_decap_8 FILLER_190_1416 ();
 sg13g2_decap_8 FILLER_190_1423 ();
 sg13g2_decap_8 FILLER_190_1430 ();
 sg13g2_decap_8 FILLER_190_1437 ();
 sg13g2_decap_8 FILLER_190_1444 ();
 sg13g2_decap_8 FILLER_190_1451 ();
 sg13g2_decap_8 FILLER_190_1458 ();
 sg13g2_decap_8 FILLER_190_1465 ();
 sg13g2_decap_8 FILLER_190_1472 ();
 sg13g2_decap_8 FILLER_190_1479 ();
 sg13g2_decap_8 FILLER_190_1486 ();
 sg13g2_decap_8 FILLER_190_1493 ();
 sg13g2_decap_8 FILLER_190_1500 ();
 sg13g2_decap_8 FILLER_190_1507 ();
 sg13g2_decap_8 FILLER_190_1514 ();
 sg13g2_decap_8 FILLER_190_1521 ();
 sg13g2_decap_8 FILLER_190_1528 ();
 sg13g2_decap_8 FILLER_190_1535 ();
 sg13g2_decap_8 FILLER_190_1542 ();
 sg13g2_decap_8 FILLER_190_1549 ();
 sg13g2_decap_8 FILLER_190_1556 ();
 sg13g2_decap_8 FILLER_190_1563 ();
 sg13g2_decap_8 FILLER_190_1570 ();
 sg13g2_decap_8 FILLER_190_1577 ();
 sg13g2_decap_8 FILLER_190_1584 ();
 sg13g2_decap_8 FILLER_190_1591 ();
 sg13g2_decap_8 FILLER_190_1598 ();
 sg13g2_decap_8 FILLER_190_1605 ();
 sg13g2_decap_8 FILLER_190_1612 ();
 sg13g2_decap_4 FILLER_190_1619 ();
 sg13g2_fill_2 FILLER_190_1623 ();
 sg13g2_decap_8 FILLER_191_0 ();
 sg13g2_decap_8 FILLER_191_7 ();
 sg13g2_decap_8 FILLER_191_14 ();
 sg13g2_decap_8 FILLER_191_21 ();
 sg13g2_decap_8 FILLER_191_28 ();
 sg13g2_decap_8 FILLER_191_35 ();
 sg13g2_decap_8 FILLER_191_42 ();
 sg13g2_decap_8 FILLER_191_49 ();
 sg13g2_decap_8 FILLER_191_56 ();
 sg13g2_decap_8 FILLER_191_63 ();
 sg13g2_decap_8 FILLER_191_70 ();
 sg13g2_decap_8 FILLER_191_77 ();
 sg13g2_decap_8 FILLER_191_84 ();
 sg13g2_decap_8 FILLER_191_91 ();
 sg13g2_decap_8 FILLER_191_98 ();
 sg13g2_decap_8 FILLER_191_105 ();
 sg13g2_decap_8 FILLER_191_112 ();
 sg13g2_decap_8 FILLER_191_119 ();
 sg13g2_decap_8 FILLER_191_126 ();
 sg13g2_decap_8 FILLER_191_133 ();
 sg13g2_decap_8 FILLER_191_140 ();
 sg13g2_decap_8 FILLER_191_147 ();
 sg13g2_decap_8 FILLER_191_154 ();
 sg13g2_decap_8 FILLER_191_161 ();
 sg13g2_decap_8 FILLER_191_168 ();
 sg13g2_decap_8 FILLER_191_175 ();
 sg13g2_decap_8 FILLER_191_182 ();
 sg13g2_decap_8 FILLER_191_189 ();
 sg13g2_decap_8 FILLER_191_196 ();
 sg13g2_decap_8 FILLER_191_203 ();
 sg13g2_decap_8 FILLER_191_210 ();
 sg13g2_decap_8 FILLER_191_217 ();
 sg13g2_decap_8 FILLER_191_224 ();
 sg13g2_decap_8 FILLER_191_231 ();
 sg13g2_decap_8 FILLER_191_238 ();
 sg13g2_decap_8 FILLER_191_245 ();
 sg13g2_decap_8 FILLER_191_252 ();
 sg13g2_decap_8 FILLER_191_259 ();
 sg13g2_decap_8 FILLER_191_266 ();
 sg13g2_decap_8 FILLER_191_273 ();
 sg13g2_decap_8 FILLER_191_280 ();
 sg13g2_decap_8 FILLER_191_287 ();
 sg13g2_decap_8 FILLER_191_294 ();
 sg13g2_fill_1 FILLER_191_301 ();
 sg13g2_decap_8 FILLER_191_306 ();
 sg13g2_decap_4 FILLER_191_313 ();
 sg13g2_fill_1 FILLER_191_317 ();
 sg13g2_decap_4 FILLER_191_326 ();
 sg13g2_fill_2 FILLER_191_330 ();
 sg13g2_decap_8 FILLER_191_336 ();
 sg13g2_fill_2 FILLER_191_343 ();
 sg13g2_fill_2 FILLER_191_356 ();
 sg13g2_fill_2 FILLER_191_368 ();
 sg13g2_decap_8 FILLER_191_384 ();
 sg13g2_fill_2 FILLER_191_391 ();
 sg13g2_decap_8 FILLER_191_415 ();
 sg13g2_decap_8 FILLER_191_422 ();
 sg13g2_fill_2 FILLER_191_481 ();
 sg13g2_decap_8 FILLER_191_487 ();
 sg13g2_decap_8 FILLER_191_494 ();
 sg13g2_decap_4 FILLER_191_515 ();
 sg13g2_fill_2 FILLER_191_519 ();
 sg13g2_fill_2 FILLER_191_572 ();
 sg13g2_fill_1 FILLER_191_574 ();
 sg13g2_fill_2 FILLER_191_609 ();
 sg13g2_fill_1 FILLER_191_611 ();
 sg13g2_fill_2 FILLER_191_616 ();
 sg13g2_decap_8 FILLER_191_623 ();
 sg13g2_decap_8 FILLER_191_630 ();
 sg13g2_decap_4 FILLER_191_637 ();
 sg13g2_fill_2 FILLER_191_641 ();
 sg13g2_decap_4 FILLER_191_652 ();
 sg13g2_fill_1 FILLER_191_656 ();
 sg13g2_decap_4 FILLER_191_661 ();
 sg13g2_fill_1 FILLER_191_665 ();
 sg13g2_decap_8 FILLER_191_671 ();
 sg13g2_fill_1 FILLER_191_678 ();
 sg13g2_fill_2 FILLER_191_708 ();
 sg13g2_decap_8 FILLER_191_749 ();
 sg13g2_decap_8 FILLER_191_756 ();
 sg13g2_decap_8 FILLER_191_763 ();
 sg13g2_decap_8 FILLER_191_770 ();
 sg13g2_decap_8 FILLER_191_777 ();
 sg13g2_fill_2 FILLER_191_784 ();
 sg13g2_fill_1 FILLER_191_786 ();
 sg13g2_decap_8 FILLER_191_813 ();
 sg13g2_fill_2 FILLER_191_820 ();
 sg13g2_fill_1 FILLER_191_822 ();
 sg13g2_decap_8 FILLER_191_827 ();
 sg13g2_decap_4 FILLER_191_834 ();
 sg13g2_fill_2 FILLER_191_838 ();
 sg13g2_fill_2 FILLER_191_848 ();
 sg13g2_fill_2 FILLER_191_860 ();
 sg13g2_fill_1 FILLER_191_862 ();
 sg13g2_fill_2 FILLER_191_914 ();
 sg13g2_fill_1 FILLER_191_916 ();
 sg13g2_decap_4 FILLER_191_925 ();
 sg13g2_fill_2 FILLER_191_929 ();
 sg13g2_fill_2 FILLER_191_957 ();
 sg13g2_decap_4 FILLER_191_963 ();
 sg13g2_fill_1 FILLER_191_967 ();
 sg13g2_decap_8 FILLER_191_972 ();
 sg13g2_decap_8 FILLER_191_979 ();
 sg13g2_decap_8 FILLER_191_986 ();
 sg13g2_decap_8 FILLER_191_993 ();
 sg13g2_decap_8 FILLER_191_1000 ();
 sg13g2_decap_8 FILLER_191_1007 ();
 sg13g2_decap_8 FILLER_191_1014 ();
 sg13g2_decap_8 FILLER_191_1021 ();
 sg13g2_decap_8 FILLER_191_1028 ();
 sg13g2_decap_8 FILLER_191_1035 ();
 sg13g2_decap_8 FILLER_191_1042 ();
 sg13g2_decap_8 FILLER_191_1049 ();
 sg13g2_decap_8 FILLER_191_1056 ();
 sg13g2_decap_8 FILLER_191_1063 ();
 sg13g2_decap_8 FILLER_191_1070 ();
 sg13g2_decap_8 FILLER_191_1077 ();
 sg13g2_decap_8 FILLER_191_1084 ();
 sg13g2_decap_8 FILLER_191_1091 ();
 sg13g2_decap_8 FILLER_191_1098 ();
 sg13g2_decap_8 FILLER_191_1105 ();
 sg13g2_decap_8 FILLER_191_1112 ();
 sg13g2_decap_8 FILLER_191_1119 ();
 sg13g2_decap_8 FILLER_191_1126 ();
 sg13g2_decap_8 FILLER_191_1133 ();
 sg13g2_decap_8 FILLER_191_1140 ();
 sg13g2_decap_8 FILLER_191_1147 ();
 sg13g2_decap_8 FILLER_191_1154 ();
 sg13g2_decap_8 FILLER_191_1161 ();
 sg13g2_decap_8 FILLER_191_1168 ();
 sg13g2_decap_8 FILLER_191_1175 ();
 sg13g2_decap_8 FILLER_191_1182 ();
 sg13g2_decap_8 FILLER_191_1189 ();
 sg13g2_decap_8 FILLER_191_1196 ();
 sg13g2_decap_8 FILLER_191_1203 ();
 sg13g2_decap_8 FILLER_191_1210 ();
 sg13g2_decap_8 FILLER_191_1217 ();
 sg13g2_decap_8 FILLER_191_1224 ();
 sg13g2_decap_8 FILLER_191_1231 ();
 sg13g2_decap_8 FILLER_191_1238 ();
 sg13g2_decap_8 FILLER_191_1245 ();
 sg13g2_decap_8 FILLER_191_1252 ();
 sg13g2_decap_8 FILLER_191_1259 ();
 sg13g2_decap_8 FILLER_191_1266 ();
 sg13g2_decap_8 FILLER_191_1273 ();
 sg13g2_decap_8 FILLER_191_1280 ();
 sg13g2_decap_8 FILLER_191_1287 ();
 sg13g2_decap_8 FILLER_191_1294 ();
 sg13g2_decap_8 FILLER_191_1301 ();
 sg13g2_decap_8 FILLER_191_1308 ();
 sg13g2_decap_8 FILLER_191_1315 ();
 sg13g2_decap_8 FILLER_191_1322 ();
 sg13g2_decap_8 FILLER_191_1329 ();
 sg13g2_decap_8 FILLER_191_1336 ();
 sg13g2_decap_8 FILLER_191_1343 ();
 sg13g2_decap_8 FILLER_191_1350 ();
 sg13g2_decap_8 FILLER_191_1357 ();
 sg13g2_decap_8 FILLER_191_1364 ();
 sg13g2_decap_8 FILLER_191_1371 ();
 sg13g2_decap_8 FILLER_191_1378 ();
 sg13g2_decap_8 FILLER_191_1385 ();
 sg13g2_decap_8 FILLER_191_1392 ();
 sg13g2_decap_8 FILLER_191_1399 ();
 sg13g2_decap_8 FILLER_191_1406 ();
 sg13g2_decap_8 FILLER_191_1413 ();
 sg13g2_decap_8 FILLER_191_1420 ();
 sg13g2_decap_8 FILLER_191_1427 ();
 sg13g2_decap_8 FILLER_191_1434 ();
 sg13g2_decap_8 FILLER_191_1441 ();
 sg13g2_decap_8 FILLER_191_1448 ();
 sg13g2_decap_8 FILLER_191_1455 ();
 sg13g2_decap_8 FILLER_191_1462 ();
 sg13g2_decap_8 FILLER_191_1469 ();
 sg13g2_decap_8 FILLER_191_1476 ();
 sg13g2_decap_8 FILLER_191_1483 ();
 sg13g2_decap_8 FILLER_191_1490 ();
 sg13g2_decap_8 FILLER_191_1497 ();
 sg13g2_decap_8 FILLER_191_1504 ();
 sg13g2_decap_8 FILLER_191_1511 ();
 sg13g2_decap_8 FILLER_191_1518 ();
 sg13g2_decap_8 FILLER_191_1525 ();
 sg13g2_decap_8 FILLER_191_1532 ();
 sg13g2_decap_8 FILLER_191_1539 ();
 sg13g2_decap_8 FILLER_191_1546 ();
 sg13g2_decap_8 FILLER_191_1553 ();
 sg13g2_decap_8 FILLER_191_1560 ();
 sg13g2_decap_8 FILLER_191_1567 ();
 sg13g2_decap_8 FILLER_191_1574 ();
 sg13g2_decap_8 FILLER_191_1581 ();
 sg13g2_decap_8 FILLER_191_1588 ();
 sg13g2_decap_8 FILLER_191_1595 ();
 sg13g2_decap_8 FILLER_191_1602 ();
 sg13g2_decap_8 FILLER_191_1609 ();
 sg13g2_decap_8 FILLER_191_1616 ();
 sg13g2_fill_2 FILLER_191_1623 ();
 sg13g2_decap_8 FILLER_192_0 ();
 sg13g2_decap_8 FILLER_192_7 ();
 sg13g2_decap_8 FILLER_192_14 ();
 sg13g2_decap_8 FILLER_192_21 ();
 sg13g2_decap_8 FILLER_192_28 ();
 sg13g2_decap_8 FILLER_192_35 ();
 sg13g2_decap_8 FILLER_192_42 ();
 sg13g2_decap_8 FILLER_192_49 ();
 sg13g2_decap_8 FILLER_192_56 ();
 sg13g2_decap_8 FILLER_192_63 ();
 sg13g2_decap_8 FILLER_192_70 ();
 sg13g2_decap_8 FILLER_192_77 ();
 sg13g2_decap_8 FILLER_192_84 ();
 sg13g2_decap_8 FILLER_192_91 ();
 sg13g2_decap_8 FILLER_192_98 ();
 sg13g2_decap_8 FILLER_192_105 ();
 sg13g2_decap_8 FILLER_192_112 ();
 sg13g2_decap_8 FILLER_192_119 ();
 sg13g2_decap_8 FILLER_192_126 ();
 sg13g2_decap_8 FILLER_192_133 ();
 sg13g2_decap_8 FILLER_192_140 ();
 sg13g2_decap_8 FILLER_192_147 ();
 sg13g2_decap_8 FILLER_192_154 ();
 sg13g2_decap_8 FILLER_192_161 ();
 sg13g2_decap_8 FILLER_192_168 ();
 sg13g2_decap_8 FILLER_192_175 ();
 sg13g2_decap_8 FILLER_192_182 ();
 sg13g2_decap_8 FILLER_192_189 ();
 sg13g2_decap_8 FILLER_192_196 ();
 sg13g2_decap_8 FILLER_192_203 ();
 sg13g2_decap_8 FILLER_192_210 ();
 sg13g2_decap_8 FILLER_192_217 ();
 sg13g2_decap_8 FILLER_192_224 ();
 sg13g2_decap_8 FILLER_192_231 ();
 sg13g2_decap_8 FILLER_192_238 ();
 sg13g2_decap_8 FILLER_192_245 ();
 sg13g2_decap_8 FILLER_192_252 ();
 sg13g2_decap_8 FILLER_192_259 ();
 sg13g2_decap_8 FILLER_192_266 ();
 sg13g2_decap_8 FILLER_192_273 ();
 sg13g2_decap_8 FILLER_192_280 ();
 sg13g2_decap_8 FILLER_192_287 ();
 sg13g2_decap_8 FILLER_192_294 ();
 sg13g2_fill_2 FILLER_192_301 ();
 sg13g2_fill_1 FILLER_192_329 ();
 sg13g2_fill_2 FILLER_192_339 ();
 sg13g2_fill_1 FILLER_192_350 ();
 sg13g2_decap_8 FILLER_192_359 ();
 sg13g2_decap_4 FILLER_192_377 ();
 sg13g2_decap_8 FILLER_192_385 ();
 sg13g2_decap_8 FILLER_192_392 ();
 sg13g2_decap_8 FILLER_192_399 ();
 sg13g2_fill_1 FILLER_192_406 ();
 sg13g2_decap_8 FILLER_192_422 ();
 sg13g2_fill_2 FILLER_192_434 ();
 sg13g2_fill_1 FILLER_192_469 ();
 sg13g2_fill_2 FILLER_192_473 ();
 sg13g2_decap_8 FILLER_192_501 ();
 sg13g2_decap_8 FILLER_192_508 ();
 sg13g2_decap_8 FILLER_192_515 ();
 sg13g2_decap_8 FILLER_192_522 ();
 sg13g2_decap_8 FILLER_192_529 ();
 sg13g2_fill_2 FILLER_192_536 ();
 sg13g2_fill_1 FILLER_192_538 ();
 sg13g2_decap_8 FILLER_192_551 ();
 sg13g2_decap_4 FILLER_192_558 ();
 sg13g2_fill_2 FILLER_192_597 ();
 sg13g2_decap_8 FILLER_192_603 ();
 sg13g2_fill_2 FILLER_192_640 ();
 sg13g2_fill_1 FILLER_192_642 ();
 sg13g2_fill_1 FILLER_192_647 ();
 sg13g2_decap_8 FILLER_192_652 ();
 sg13g2_decap_4 FILLER_192_659 ();
 sg13g2_fill_2 FILLER_192_663 ();
 sg13g2_decap_4 FILLER_192_669 ();
 sg13g2_decap_8 FILLER_192_677 ();
 sg13g2_decap_4 FILLER_192_684 ();
 sg13g2_fill_1 FILLER_192_688 ();
 sg13g2_fill_1 FILLER_192_715 ();
 sg13g2_decap_8 FILLER_192_742 ();
 sg13g2_decap_4 FILLER_192_749 ();
 sg13g2_decap_8 FILLER_192_778 ();
 sg13g2_decap_4 FILLER_192_785 ();
 sg13g2_decap_8 FILLER_192_799 ();
 sg13g2_decap_8 FILLER_192_806 ();
 sg13g2_fill_2 FILLER_192_813 ();
 sg13g2_fill_1 FILLER_192_815 ();
 sg13g2_decap_4 FILLER_192_846 ();
 sg13g2_fill_1 FILLER_192_850 ();
 sg13g2_decap_8 FILLER_192_855 ();
 sg13g2_decap_4 FILLER_192_862 ();
 sg13g2_decap_8 FILLER_192_878 ();
 sg13g2_decap_4 FILLER_192_885 ();
 sg13g2_decap_4 FILLER_192_902 ();
 sg13g2_fill_1 FILLER_192_906 ();
 sg13g2_fill_1 FILLER_192_915 ();
 sg13g2_decap_8 FILLER_192_928 ();
 sg13g2_fill_1 FILLER_192_935 ();
 sg13g2_decap_4 FILLER_192_940 ();
 sg13g2_fill_1 FILLER_192_944 ();
 sg13g2_decap_8 FILLER_192_948 ();
 sg13g2_decap_4 FILLER_192_955 ();
 sg13g2_fill_1 FILLER_192_959 ();
 sg13g2_decap_8 FILLER_192_986 ();
 sg13g2_decap_8 FILLER_192_993 ();
 sg13g2_decap_8 FILLER_192_1000 ();
 sg13g2_decap_8 FILLER_192_1007 ();
 sg13g2_decap_8 FILLER_192_1014 ();
 sg13g2_decap_8 FILLER_192_1021 ();
 sg13g2_decap_8 FILLER_192_1028 ();
 sg13g2_decap_8 FILLER_192_1035 ();
 sg13g2_decap_8 FILLER_192_1042 ();
 sg13g2_decap_8 FILLER_192_1049 ();
 sg13g2_decap_8 FILLER_192_1056 ();
 sg13g2_decap_8 FILLER_192_1063 ();
 sg13g2_decap_8 FILLER_192_1070 ();
 sg13g2_decap_8 FILLER_192_1077 ();
 sg13g2_decap_8 FILLER_192_1084 ();
 sg13g2_decap_8 FILLER_192_1091 ();
 sg13g2_decap_8 FILLER_192_1098 ();
 sg13g2_decap_8 FILLER_192_1105 ();
 sg13g2_decap_8 FILLER_192_1112 ();
 sg13g2_decap_8 FILLER_192_1119 ();
 sg13g2_decap_8 FILLER_192_1126 ();
 sg13g2_decap_8 FILLER_192_1133 ();
 sg13g2_decap_8 FILLER_192_1140 ();
 sg13g2_decap_8 FILLER_192_1147 ();
 sg13g2_decap_8 FILLER_192_1154 ();
 sg13g2_decap_8 FILLER_192_1161 ();
 sg13g2_decap_8 FILLER_192_1168 ();
 sg13g2_decap_8 FILLER_192_1175 ();
 sg13g2_decap_8 FILLER_192_1182 ();
 sg13g2_decap_8 FILLER_192_1189 ();
 sg13g2_decap_8 FILLER_192_1196 ();
 sg13g2_decap_8 FILLER_192_1203 ();
 sg13g2_decap_8 FILLER_192_1210 ();
 sg13g2_decap_8 FILLER_192_1217 ();
 sg13g2_decap_8 FILLER_192_1224 ();
 sg13g2_decap_8 FILLER_192_1231 ();
 sg13g2_decap_8 FILLER_192_1238 ();
 sg13g2_decap_8 FILLER_192_1245 ();
 sg13g2_decap_8 FILLER_192_1252 ();
 sg13g2_decap_8 FILLER_192_1259 ();
 sg13g2_decap_8 FILLER_192_1266 ();
 sg13g2_decap_8 FILLER_192_1273 ();
 sg13g2_decap_8 FILLER_192_1280 ();
 sg13g2_decap_8 FILLER_192_1287 ();
 sg13g2_decap_8 FILLER_192_1294 ();
 sg13g2_decap_8 FILLER_192_1301 ();
 sg13g2_decap_8 FILLER_192_1308 ();
 sg13g2_decap_8 FILLER_192_1315 ();
 sg13g2_decap_8 FILLER_192_1322 ();
 sg13g2_decap_8 FILLER_192_1329 ();
 sg13g2_decap_8 FILLER_192_1336 ();
 sg13g2_decap_8 FILLER_192_1343 ();
 sg13g2_decap_8 FILLER_192_1350 ();
 sg13g2_decap_8 FILLER_192_1357 ();
 sg13g2_decap_8 FILLER_192_1364 ();
 sg13g2_decap_8 FILLER_192_1371 ();
 sg13g2_decap_8 FILLER_192_1378 ();
 sg13g2_decap_8 FILLER_192_1385 ();
 sg13g2_decap_8 FILLER_192_1392 ();
 sg13g2_decap_8 FILLER_192_1399 ();
 sg13g2_decap_8 FILLER_192_1406 ();
 sg13g2_decap_8 FILLER_192_1413 ();
 sg13g2_decap_8 FILLER_192_1420 ();
 sg13g2_decap_8 FILLER_192_1427 ();
 sg13g2_decap_8 FILLER_192_1434 ();
 sg13g2_decap_8 FILLER_192_1441 ();
 sg13g2_decap_8 FILLER_192_1448 ();
 sg13g2_decap_8 FILLER_192_1455 ();
 sg13g2_decap_8 FILLER_192_1462 ();
 sg13g2_decap_8 FILLER_192_1469 ();
 sg13g2_decap_8 FILLER_192_1476 ();
 sg13g2_decap_8 FILLER_192_1483 ();
 sg13g2_decap_8 FILLER_192_1490 ();
 sg13g2_decap_8 FILLER_192_1497 ();
 sg13g2_decap_8 FILLER_192_1504 ();
 sg13g2_decap_8 FILLER_192_1511 ();
 sg13g2_decap_8 FILLER_192_1518 ();
 sg13g2_decap_8 FILLER_192_1525 ();
 sg13g2_decap_8 FILLER_192_1532 ();
 sg13g2_decap_8 FILLER_192_1539 ();
 sg13g2_decap_8 FILLER_192_1546 ();
 sg13g2_decap_8 FILLER_192_1553 ();
 sg13g2_decap_8 FILLER_192_1560 ();
 sg13g2_decap_8 FILLER_192_1567 ();
 sg13g2_decap_8 FILLER_192_1574 ();
 sg13g2_decap_8 FILLER_192_1581 ();
 sg13g2_decap_8 FILLER_192_1588 ();
 sg13g2_decap_8 FILLER_192_1595 ();
 sg13g2_decap_8 FILLER_192_1602 ();
 sg13g2_decap_8 FILLER_192_1609 ();
 sg13g2_decap_8 FILLER_192_1616 ();
 sg13g2_fill_2 FILLER_192_1623 ();
 sg13g2_decap_8 FILLER_193_0 ();
 sg13g2_decap_8 FILLER_193_7 ();
 sg13g2_decap_8 FILLER_193_14 ();
 sg13g2_decap_8 FILLER_193_21 ();
 sg13g2_decap_8 FILLER_193_28 ();
 sg13g2_decap_8 FILLER_193_35 ();
 sg13g2_decap_8 FILLER_193_42 ();
 sg13g2_decap_8 FILLER_193_49 ();
 sg13g2_decap_8 FILLER_193_56 ();
 sg13g2_decap_8 FILLER_193_63 ();
 sg13g2_decap_8 FILLER_193_70 ();
 sg13g2_decap_8 FILLER_193_77 ();
 sg13g2_decap_8 FILLER_193_84 ();
 sg13g2_decap_8 FILLER_193_91 ();
 sg13g2_decap_8 FILLER_193_98 ();
 sg13g2_decap_8 FILLER_193_105 ();
 sg13g2_decap_8 FILLER_193_112 ();
 sg13g2_decap_8 FILLER_193_119 ();
 sg13g2_decap_8 FILLER_193_126 ();
 sg13g2_decap_8 FILLER_193_133 ();
 sg13g2_decap_8 FILLER_193_140 ();
 sg13g2_decap_8 FILLER_193_147 ();
 sg13g2_decap_8 FILLER_193_154 ();
 sg13g2_decap_8 FILLER_193_161 ();
 sg13g2_decap_8 FILLER_193_168 ();
 sg13g2_decap_8 FILLER_193_175 ();
 sg13g2_decap_8 FILLER_193_182 ();
 sg13g2_decap_8 FILLER_193_189 ();
 sg13g2_decap_8 FILLER_193_196 ();
 sg13g2_decap_8 FILLER_193_203 ();
 sg13g2_decap_8 FILLER_193_210 ();
 sg13g2_decap_8 FILLER_193_217 ();
 sg13g2_decap_8 FILLER_193_224 ();
 sg13g2_decap_8 FILLER_193_231 ();
 sg13g2_decap_8 FILLER_193_238 ();
 sg13g2_decap_8 FILLER_193_245 ();
 sg13g2_decap_8 FILLER_193_252 ();
 sg13g2_decap_8 FILLER_193_259 ();
 sg13g2_decap_8 FILLER_193_266 ();
 sg13g2_decap_8 FILLER_193_273 ();
 sg13g2_decap_8 FILLER_193_280 ();
 sg13g2_decap_8 FILLER_193_287 ();
 sg13g2_decap_8 FILLER_193_294 ();
 sg13g2_decap_8 FILLER_193_301 ();
 sg13g2_decap_4 FILLER_193_308 ();
 sg13g2_decap_8 FILLER_193_316 ();
 sg13g2_decap_8 FILLER_193_323 ();
 sg13g2_decap_8 FILLER_193_330 ();
 sg13g2_fill_1 FILLER_193_337 ();
 sg13g2_fill_1 FILLER_193_343 ();
 sg13g2_fill_2 FILLER_193_360 ();
 sg13g2_fill_1 FILLER_193_362 ();
 sg13g2_fill_1 FILLER_193_369 ();
 sg13g2_decap_4 FILLER_193_379 ();
 sg13g2_fill_2 FILLER_193_383 ();
 sg13g2_decap_4 FILLER_193_390 ();
 sg13g2_fill_2 FILLER_193_394 ();
 sg13g2_fill_2 FILLER_193_467 ();
 sg13g2_fill_1 FILLER_193_469 ();
 sg13g2_decap_8 FILLER_193_495 ();
 sg13g2_decap_8 FILLER_193_502 ();
 sg13g2_fill_1 FILLER_193_514 ();
 sg13g2_fill_2 FILLER_193_520 ();
 sg13g2_fill_1 FILLER_193_522 ();
 sg13g2_decap_4 FILLER_193_528 ();
 sg13g2_fill_2 FILLER_193_548 ();
 sg13g2_fill_1 FILLER_193_550 ();
 sg13g2_decap_4 FILLER_193_560 ();
 sg13g2_fill_2 FILLER_193_564 ();
 sg13g2_fill_2 FILLER_193_604 ();
 sg13g2_fill_1 FILLER_193_606 ();
 sg13g2_fill_1 FILLER_193_611 ();
 sg13g2_fill_2 FILLER_193_637 ();
 sg13g2_decap_4 FILLER_193_694 ();
 sg13g2_decap_4 FILLER_193_703 ();
 sg13g2_fill_1 FILLER_193_707 ();
 sg13g2_decap_8 FILLER_193_758 ();
 sg13g2_decap_8 FILLER_193_765 ();
 sg13g2_decap_8 FILLER_193_772 ();
 sg13g2_decap_8 FILLER_193_779 ();
 sg13g2_decap_8 FILLER_193_786 ();
 sg13g2_decap_8 FILLER_193_793 ();
 sg13g2_decap_8 FILLER_193_800 ();
 sg13g2_decap_8 FILLER_193_807 ();
 sg13g2_decap_8 FILLER_193_814 ();
 sg13g2_decap_8 FILLER_193_821 ();
 sg13g2_decap_8 FILLER_193_828 ();
 sg13g2_decap_8 FILLER_193_835 ();
 sg13g2_fill_2 FILLER_193_842 ();
 sg13g2_fill_1 FILLER_193_844 ();
 sg13g2_fill_1 FILLER_193_857 ();
 sg13g2_fill_1 FILLER_193_916 ();
 sg13g2_fill_2 FILLER_193_926 ();
 sg13g2_decap_8 FILLER_193_954 ();
 sg13g2_decap_8 FILLER_193_961 ();
 sg13g2_decap_8 FILLER_193_968 ();
 sg13g2_decap_8 FILLER_193_975 ();
 sg13g2_decap_8 FILLER_193_982 ();
 sg13g2_decap_8 FILLER_193_989 ();
 sg13g2_decap_8 FILLER_193_996 ();
 sg13g2_decap_8 FILLER_193_1003 ();
 sg13g2_decap_8 FILLER_193_1010 ();
 sg13g2_decap_8 FILLER_193_1017 ();
 sg13g2_decap_8 FILLER_193_1024 ();
 sg13g2_decap_8 FILLER_193_1031 ();
 sg13g2_decap_8 FILLER_193_1038 ();
 sg13g2_decap_8 FILLER_193_1045 ();
 sg13g2_decap_8 FILLER_193_1052 ();
 sg13g2_decap_8 FILLER_193_1059 ();
 sg13g2_decap_8 FILLER_193_1066 ();
 sg13g2_decap_8 FILLER_193_1073 ();
 sg13g2_decap_8 FILLER_193_1080 ();
 sg13g2_decap_8 FILLER_193_1087 ();
 sg13g2_decap_8 FILLER_193_1094 ();
 sg13g2_decap_8 FILLER_193_1101 ();
 sg13g2_decap_8 FILLER_193_1108 ();
 sg13g2_decap_8 FILLER_193_1115 ();
 sg13g2_decap_8 FILLER_193_1122 ();
 sg13g2_decap_8 FILLER_193_1129 ();
 sg13g2_decap_8 FILLER_193_1136 ();
 sg13g2_decap_8 FILLER_193_1143 ();
 sg13g2_decap_8 FILLER_193_1150 ();
 sg13g2_decap_8 FILLER_193_1157 ();
 sg13g2_decap_8 FILLER_193_1164 ();
 sg13g2_decap_8 FILLER_193_1171 ();
 sg13g2_decap_8 FILLER_193_1178 ();
 sg13g2_decap_8 FILLER_193_1185 ();
 sg13g2_decap_8 FILLER_193_1192 ();
 sg13g2_decap_8 FILLER_193_1199 ();
 sg13g2_decap_8 FILLER_193_1206 ();
 sg13g2_decap_8 FILLER_193_1213 ();
 sg13g2_decap_8 FILLER_193_1220 ();
 sg13g2_decap_8 FILLER_193_1227 ();
 sg13g2_decap_8 FILLER_193_1234 ();
 sg13g2_decap_8 FILLER_193_1241 ();
 sg13g2_decap_8 FILLER_193_1248 ();
 sg13g2_decap_8 FILLER_193_1255 ();
 sg13g2_decap_8 FILLER_193_1262 ();
 sg13g2_decap_8 FILLER_193_1269 ();
 sg13g2_decap_8 FILLER_193_1276 ();
 sg13g2_decap_8 FILLER_193_1283 ();
 sg13g2_decap_8 FILLER_193_1290 ();
 sg13g2_decap_8 FILLER_193_1297 ();
 sg13g2_decap_8 FILLER_193_1304 ();
 sg13g2_decap_8 FILLER_193_1311 ();
 sg13g2_decap_8 FILLER_193_1318 ();
 sg13g2_decap_8 FILLER_193_1325 ();
 sg13g2_decap_8 FILLER_193_1332 ();
 sg13g2_decap_8 FILLER_193_1339 ();
 sg13g2_decap_8 FILLER_193_1346 ();
 sg13g2_decap_8 FILLER_193_1353 ();
 sg13g2_decap_8 FILLER_193_1360 ();
 sg13g2_decap_8 FILLER_193_1367 ();
 sg13g2_decap_8 FILLER_193_1374 ();
 sg13g2_decap_8 FILLER_193_1381 ();
 sg13g2_decap_8 FILLER_193_1388 ();
 sg13g2_decap_8 FILLER_193_1395 ();
 sg13g2_decap_8 FILLER_193_1402 ();
 sg13g2_decap_8 FILLER_193_1409 ();
 sg13g2_decap_8 FILLER_193_1416 ();
 sg13g2_decap_8 FILLER_193_1423 ();
 sg13g2_decap_8 FILLER_193_1430 ();
 sg13g2_decap_8 FILLER_193_1437 ();
 sg13g2_decap_8 FILLER_193_1444 ();
 sg13g2_decap_8 FILLER_193_1451 ();
 sg13g2_decap_8 FILLER_193_1458 ();
 sg13g2_decap_8 FILLER_193_1465 ();
 sg13g2_decap_8 FILLER_193_1472 ();
 sg13g2_decap_8 FILLER_193_1479 ();
 sg13g2_decap_8 FILLER_193_1486 ();
 sg13g2_decap_8 FILLER_193_1493 ();
 sg13g2_decap_8 FILLER_193_1500 ();
 sg13g2_decap_8 FILLER_193_1507 ();
 sg13g2_decap_8 FILLER_193_1514 ();
 sg13g2_decap_8 FILLER_193_1521 ();
 sg13g2_decap_8 FILLER_193_1528 ();
 sg13g2_decap_8 FILLER_193_1535 ();
 sg13g2_decap_8 FILLER_193_1542 ();
 sg13g2_decap_8 FILLER_193_1549 ();
 sg13g2_decap_8 FILLER_193_1556 ();
 sg13g2_decap_8 FILLER_193_1563 ();
 sg13g2_decap_8 FILLER_193_1570 ();
 sg13g2_decap_8 FILLER_193_1577 ();
 sg13g2_decap_8 FILLER_193_1584 ();
 sg13g2_decap_8 FILLER_193_1591 ();
 sg13g2_decap_8 FILLER_193_1598 ();
 sg13g2_decap_8 FILLER_193_1605 ();
 sg13g2_decap_8 FILLER_193_1612 ();
 sg13g2_decap_4 FILLER_193_1619 ();
 sg13g2_fill_2 FILLER_193_1623 ();
 sg13g2_decap_8 FILLER_194_0 ();
 sg13g2_decap_8 FILLER_194_7 ();
 sg13g2_decap_8 FILLER_194_14 ();
 sg13g2_decap_8 FILLER_194_21 ();
 sg13g2_decap_8 FILLER_194_28 ();
 sg13g2_decap_8 FILLER_194_35 ();
 sg13g2_decap_8 FILLER_194_42 ();
 sg13g2_decap_8 FILLER_194_49 ();
 sg13g2_decap_8 FILLER_194_56 ();
 sg13g2_decap_8 FILLER_194_63 ();
 sg13g2_decap_8 FILLER_194_70 ();
 sg13g2_decap_8 FILLER_194_77 ();
 sg13g2_decap_8 FILLER_194_84 ();
 sg13g2_decap_8 FILLER_194_91 ();
 sg13g2_decap_8 FILLER_194_98 ();
 sg13g2_decap_8 FILLER_194_105 ();
 sg13g2_decap_8 FILLER_194_112 ();
 sg13g2_decap_8 FILLER_194_119 ();
 sg13g2_decap_8 FILLER_194_126 ();
 sg13g2_decap_8 FILLER_194_133 ();
 sg13g2_decap_8 FILLER_194_140 ();
 sg13g2_decap_8 FILLER_194_147 ();
 sg13g2_decap_8 FILLER_194_154 ();
 sg13g2_decap_8 FILLER_194_161 ();
 sg13g2_decap_8 FILLER_194_168 ();
 sg13g2_decap_8 FILLER_194_175 ();
 sg13g2_decap_8 FILLER_194_182 ();
 sg13g2_decap_8 FILLER_194_189 ();
 sg13g2_decap_8 FILLER_194_196 ();
 sg13g2_decap_8 FILLER_194_203 ();
 sg13g2_decap_8 FILLER_194_210 ();
 sg13g2_decap_8 FILLER_194_217 ();
 sg13g2_decap_8 FILLER_194_224 ();
 sg13g2_decap_8 FILLER_194_231 ();
 sg13g2_decap_8 FILLER_194_238 ();
 sg13g2_decap_8 FILLER_194_245 ();
 sg13g2_decap_8 FILLER_194_252 ();
 sg13g2_decap_8 FILLER_194_259 ();
 sg13g2_decap_8 FILLER_194_266 ();
 sg13g2_decap_8 FILLER_194_273 ();
 sg13g2_decap_8 FILLER_194_280 ();
 sg13g2_decap_8 FILLER_194_287 ();
 sg13g2_decap_8 FILLER_194_294 ();
 sg13g2_decap_4 FILLER_194_301 ();
 sg13g2_decap_4 FILLER_194_342 ();
 sg13g2_fill_2 FILLER_194_346 ();
 sg13g2_decap_8 FILLER_194_353 ();
 sg13g2_decap_8 FILLER_194_360 ();
 sg13g2_decap_8 FILLER_194_367 ();
 sg13g2_decap_4 FILLER_194_374 ();
 sg13g2_fill_2 FILLER_194_378 ();
 sg13g2_decap_8 FILLER_194_410 ();
 sg13g2_fill_2 FILLER_194_417 ();
 sg13g2_fill_1 FILLER_194_424 ();
 sg13g2_fill_2 FILLER_194_430 ();
 sg13g2_decap_8 FILLER_194_437 ();
 sg13g2_decap_8 FILLER_194_444 ();
 sg13g2_decap_8 FILLER_194_451 ();
 sg13g2_decap_8 FILLER_194_458 ();
 sg13g2_decap_4 FILLER_194_465 ();
 sg13g2_fill_1 FILLER_194_469 ();
 sg13g2_decap_8 FILLER_194_479 ();
 sg13g2_decap_8 FILLER_194_486 ();
 sg13g2_fill_1 FILLER_194_493 ();
 sg13g2_fill_2 FILLER_194_500 ();
 sg13g2_fill_1 FILLER_194_502 ();
 sg13g2_fill_2 FILLER_194_527 ();
 sg13g2_fill_2 FILLER_194_533 ();
 sg13g2_fill_1 FILLER_194_535 ();
 sg13g2_fill_2 FILLER_194_541 ();
 sg13g2_fill_1 FILLER_194_543 ();
 sg13g2_decap_8 FILLER_194_549 ();
 sg13g2_decap_8 FILLER_194_556 ();
 sg13g2_decap_8 FILLER_194_563 ();
 sg13g2_fill_1 FILLER_194_570 ();
 sg13g2_decap_8 FILLER_194_633 ();
 sg13g2_decap_8 FILLER_194_640 ();
 sg13g2_decap_8 FILLER_194_647 ();
 sg13g2_fill_2 FILLER_194_654 ();
 sg13g2_fill_1 FILLER_194_656 ();
 sg13g2_fill_2 FILLER_194_682 ();
 sg13g2_fill_1 FILLER_194_709 ();
 sg13g2_decap_8 FILLER_194_722 ();
 sg13g2_decap_8 FILLER_194_729 ();
 sg13g2_decap_8 FILLER_194_736 ();
 sg13g2_decap_8 FILLER_194_743 ();
 sg13g2_decap_8 FILLER_194_750 ();
 sg13g2_decap_8 FILLER_194_757 ();
 sg13g2_decap_8 FILLER_194_764 ();
 sg13g2_decap_8 FILLER_194_771 ();
 sg13g2_decap_8 FILLER_194_778 ();
 sg13g2_decap_8 FILLER_194_785 ();
 sg13g2_decap_8 FILLER_194_792 ();
 sg13g2_decap_8 FILLER_194_799 ();
 sg13g2_decap_8 FILLER_194_806 ();
 sg13g2_decap_8 FILLER_194_813 ();
 sg13g2_decap_8 FILLER_194_820 ();
 sg13g2_decap_8 FILLER_194_827 ();
 sg13g2_decap_4 FILLER_194_864 ();
 sg13g2_decap_8 FILLER_194_894 ();
 sg13g2_decap_8 FILLER_194_901 ();
 sg13g2_decap_8 FILLER_194_908 ();
 sg13g2_fill_1 FILLER_194_915 ();
 sg13g2_decap_8 FILLER_194_920 ();
 sg13g2_decap_4 FILLER_194_927 ();
 sg13g2_decap_8 FILLER_194_935 ();
 sg13g2_fill_2 FILLER_194_942 ();
 sg13g2_fill_1 FILLER_194_944 ();
 sg13g2_decap_8 FILLER_194_970 ();
 sg13g2_decap_8 FILLER_194_977 ();
 sg13g2_decap_8 FILLER_194_984 ();
 sg13g2_decap_8 FILLER_194_991 ();
 sg13g2_decap_8 FILLER_194_998 ();
 sg13g2_decap_8 FILLER_194_1005 ();
 sg13g2_decap_8 FILLER_194_1012 ();
 sg13g2_decap_8 FILLER_194_1019 ();
 sg13g2_decap_8 FILLER_194_1026 ();
 sg13g2_decap_8 FILLER_194_1033 ();
 sg13g2_decap_8 FILLER_194_1040 ();
 sg13g2_decap_8 FILLER_194_1047 ();
 sg13g2_decap_8 FILLER_194_1054 ();
 sg13g2_decap_8 FILLER_194_1061 ();
 sg13g2_decap_8 FILLER_194_1068 ();
 sg13g2_decap_8 FILLER_194_1075 ();
 sg13g2_decap_8 FILLER_194_1082 ();
 sg13g2_decap_8 FILLER_194_1089 ();
 sg13g2_decap_8 FILLER_194_1096 ();
 sg13g2_decap_8 FILLER_194_1103 ();
 sg13g2_decap_8 FILLER_194_1110 ();
 sg13g2_decap_8 FILLER_194_1117 ();
 sg13g2_decap_8 FILLER_194_1124 ();
 sg13g2_decap_8 FILLER_194_1131 ();
 sg13g2_decap_8 FILLER_194_1138 ();
 sg13g2_decap_8 FILLER_194_1145 ();
 sg13g2_decap_8 FILLER_194_1152 ();
 sg13g2_decap_8 FILLER_194_1159 ();
 sg13g2_decap_8 FILLER_194_1166 ();
 sg13g2_decap_8 FILLER_194_1173 ();
 sg13g2_decap_8 FILLER_194_1180 ();
 sg13g2_decap_8 FILLER_194_1187 ();
 sg13g2_decap_8 FILLER_194_1194 ();
 sg13g2_decap_8 FILLER_194_1201 ();
 sg13g2_decap_8 FILLER_194_1208 ();
 sg13g2_decap_8 FILLER_194_1215 ();
 sg13g2_decap_8 FILLER_194_1222 ();
 sg13g2_decap_8 FILLER_194_1229 ();
 sg13g2_decap_8 FILLER_194_1236 ();
 sg13g2_decap_8 FILLER_194_1243 ();
 sg13g2_decap_8 FILLER_194_1250 ();
 sg13g2_decap_8 FILLER_194_1257 ();
 sg13g2_decap_8 FILLER_194_1264 ();
 sg13g2_decap_8 FILLER_194_1271 ();
 sg13g2_decap_8 FILLER_194_1278 ();
 sg13g2_decap_8 FILLER_194_1285 ();
 sg13g2_decap_8 FILLER_194_1292 ();
 sg13g2_decap_8 FILLER_194_1299 ();
 sg13g2_decap_8 FILLER_194_1306 ();
 sg13g2_decap_8 FILLER_194_1313 ();
 sg13g2_decap_8 FILLER_194_1320 ();
 sg13g2_decap_8 FILLER_194_1327 ();
 sg13g2_decap_8 FILLER_194_1334 ();
 sg13g2_decap_8 FILLER_194_1341 ();
 sg13g2_decap_8 FILLER_194_1348 ();
 sg13g2_decap_8 FILLER_194_1355 ();
 sg13g2_decap_8 FILLER_194_1362 ();
 sg13g2_decap_8 FILLER_194_1369 ();
 sg13g2_decap_8 FILLER_194_1376 ();
 sg13g2_decap_8 FILLER_194_1383 ();
 sg13g2_decap_8 FILLER_194_1390 ();
 sg13g2_decap_8 FILLER_194_1397 ();
 sg13g2_decap_8 FILLER_194_1404 ();
 sg13g2_decap_8 FILLER_194_1411 ();
 sg13g2_decap_8 FILLER_194_1418 ();
 sg13g2_decap_8 FILLER_194_1425 ();
 sg13g2_decap_8 FILLER_194_1432 ();
 sg13g2_decap_8 FILLER_194_1439 ();
 sg13g2_decap_8 FILLER_194_1446 ();
 sg13g2_decap_8 FILLER_194_1453 ();
 sg13g2_decap_8 FILLER_194_1460 ();
 sg13g2_decap_8 FILLER_194_1467 ();
 sg13g2_decap_8 FILLER_194_1474 ();
 sg13g2_decap_8 FILLER_194_1481 ();
 sg13g2_decap_8 FILLER_194_1488 ();
 sg13g2_decap_8 FILLER_194_1495 ();
 sg13g2_decap_8 FILLER_194_1502 ();
 sg13g2_decap_8 FILLER_194_1509 ();
 sg13g2_decap_8 FILLER_194_1516 ();
 sg13g2_decap_8 FILLER_194_1523 ();
 sg13g2_decap_8 FILLER_194_1530 ();
 sg13g2_decap_8 FILLER_194_1537 ();
 sg13g2_decap_8 FILLER_194_1544 ();
 sg13g2_decap_8 FILLER_194_1551 ();
 sg13g2_decap_8 FILLER_194_1558 ();
 sg13g2_decap_8 FILLER_194_1565 ();
 sg13g2_decap_8 FILLER_194_1572 ();
 sg13g2_decap_8 FILLER_194_1579 ();
 sg13g2_decap_8 FILLER_194_1586 ();
 sg13g2_decap_8 FILLER_194_1593 ();
 sg13g2_decap_8 FILLER_194_1600 ();
 sg13g2_decap_8 FILLER_194_1607 ();
 sg13g2_decap_8 FILLER_194_1614 ();
 sg13g2_decap_4 FILLER_194_1621 ();
 sg13g2_decap_8 FILLER_195_0 ();
 sg13g2_decap_8 FILLER_195_7 ();
 sg13g2_decap_8 FILLER_195_14 ();
 sg13g2_decap_8 FILLER_195_21 ();
 sg13g2_decap_8 FILLER_195_28 ();
 sg13g2_decap_8 FILLER_195_35 ();
 sg13g2_decap_8 FILLER_195_42 ();
 sg13g2_decap_8 FILLER_195_49 ();
 sg13g2_decap_8 FILLER_195_56 ();
 sg13g2_decap_8 FILLER_195_63 ();
 sg13g2_decap_8 FILLER_195_70 ();
 sg13g2_decap_8 FILLER_195_77 ();
 sg13g2_decap_8 FILLER_195_84 ();
 sg13g2_decap_8 FILLER_195_91 ();
 sg13g2_decap_8 FILLER_195_98 ();
 sg13g2_decap_8 FILLER_195_105 ();
 sg13g2_decap_8 FILLER_195_112 ();
 sg13g2_decap_8 FILLER_195_119 ();
 sg13g2_decap_8 FILLER_195_126 ();
 sg13g2_decap_8 FILLER_195_133 ();
 sg13g2_decap_8 FILLER_195_140 ();
 sg13g2_decap_8 FILLER_195_147 ();
 sg13g2_decap_8 FILLER_195_154 ();
 sg13g2_decap_8 FILLER_195_161 ();
 sg13g2_decap_8 FILLER_195_168 ();
 sg13g2_decap_8 FILLER_195_175 ();
 sg13g2_decap_8 FILLER_195_182 ();
 sg13g2_decap_8 FILLER_195_189 ();
 sg13g2_decap_8 FILLER_195_196 ();
 sg13g2_decap_8 FILLER_195_203 ();
 sg13g2_decap_8 FILLER_195_210 ();
 sg13g2_decap_8 FILLER_195_217 ();
 sg13g2_decap_8 FILLER_195_224 ();
 sg13g2_decap_8 FILLER_195_231 ();
 sg13g2_decap_8 FILLER_195_238 ();
 sg13g2_decap_8 FILLER_195_245 ();
 sg13g2_decap_8 FILLER_195_252 ();
 sg13g2_decap_8 FILLER_195_259 ();
 sg13g2_decap_8 FILLER_195_266 ();
 sg13g2_decap_8 FILLER_195_273 ();
 sg13g2_decap_8 FILLER_195_280 ();
 sg13g2_decap_8 FILLER_195_287 ();
 sg13g2_decap_8 FILLER_195_294 ();
 sg13g2_decap_4 FILLER_195_349 ();
 sg13g2_fill_2 FILLER_195_353 ();
 sg13g2_decap_8 FILLER_195_359 ();
 sg13g2_decap_4 FILLER_195_366 ();
 sg13g2_decap_8 FILLER_195_382 ();
 sg13g2_decap_8 FILLER_195_393 ();
 sg13g2_decap_8 FILLER_195_400 ();
 sg13g2_decap_8 FILLER_195_419 ();
 sg13g2_decap_4 FILLER_195_426 ();
 sg13g2_decap_8 FILLER_195_434 ();
 sg13g2_decap_8 FILLER_195_441 ();
 sg13g2_decap_8 FILLER_195_448 ();
 sg13g2_decap_8 FILLER_195_455 ();
 sg13g2_fill_2 FILLER_195_462 ();
 sg13g2_fill_1 FILLER_195_480 ();
 sg13g2_fill_1 FILLER_195_486 ();
 sg13g2_fill_2 FILLER_195_492 ();
 sg13g2_fill_2 FILLER_195_499 ();
 sg13g2_fill_2 FILLER_195_506 ();
 sg13g2_decap_8 FILLER_195_516 ();
 sg13g2_fill_1 FILLER_195_523 ();
 sg13g2_fill_2 FILLER_195_532 ();
 sg13g2_fill_1 FILLER_195_534 ();
 sg13g2_fill_2 FILLER_195_553 ();
 sg13g2_fill_1 FILLER_195_555 ();
 sg13g2_decap_8 FILLER_195_563 ();
 sg13g2_decap_8 FILLER_195_570 ();
 sg13g2_fill_1 FILLER_195_577 ();
 sg13g2_fill_2 FILLER_195_603 ();
 sg13g2_decap_8 FILLER_195_613 ();
 sg13g2_fill_1 FILLER_195_623 ();
 sg13g2_fill_2 FILLER_195_631 ();
 sg13g2_fill_1 FILLER_195_638 ();
 sg13g2_decap_4 FILLER_195_655 ();
 sg13g2_decap_4 FILLER_195_672 ();
 sg13g2_fill_2 FILLER_195_682 ();
 sg13g2_fill_1 FILLER_195_684 ();
 sg13g2_fill_2 FILLER_195_698 ();
 sg13g2_decap_8 FILLER_195_722 ();
 sg13g2_decap_8 FILLER_195_729 ();
 sg13g2_decap_8 FILLER_195_736 ();
 sg13g2_decap_8 FILLER_195_743 ();
 sg13g2_decap_8 FILLER_195_750 ();
 sg13g2_decap_8 FILLER_195_757 ();
 sg13g2_decap_8 FILLER_195_764 ();
 sg13g2_decap_8 FILLER_195_771 ();
 sg13g2_decap_8 FILLER_195_778 ();
 sg13g2_decap_8 FILLER_195_785 ();
 sg13g2_decap_8 FILLER_195_792 ();
 sg13g2_decap_8 FILLER_195_799 ();
 sg13g2_decap_8 FILLER_195_806 ();
 sg13g2_decap_8 FILLER_195_813 ();
 sg13g2_decap_8 FILLER_195_820 ();
 sg13g2_decap_8 FILLER_195_827 ();
 sg13g2_decap_8 FILLER_195_834 ();
 sg13g2_decap_8 FILLER_195_841 ();
 sg13g2_decap_8 FILLER_195_848 ();
 sg13g2_decap_8 FILLER_195_855 ();
 sg13g2_decap_8 FILLER_195_862 ();
 sg13g2_decap_4 FILLER_195_869 ();
 sg13g2_fill_2 FILLER_195_873 ();
 sg13g2_decap_8 FILLER_195_879 ();
 sg13g2_decap_8 FILLER_195_886 ();
 sg13g2_decap_4 FILLER_195_893 ();
 sg13g2_fill_1 FILLER_195_897 ();
 sg13g2_fill_1 FILLER_195_902 ();
 sg13g2_fill_1 FILLER_195_907 ();
 sg13g2_fill_1 FILLER_195_912 ();
 sg13g2_fill_1 FILLER_195_921 ();
 sg13g2_decap_8 FILLER_195_948 ();
 sg13g2_decap_8 FILLER_195_955 ();
 sg13g2_decap_8 FILLER_195_962 ();
 sg13g2_decap_8 FILLER_195_969 ();
 sg13g2_decap_8 FILLER_195_976 ();
 sg13g2_decap_8 FILLER_195_983 ();
 sg13g2_decap_8 FILLER_195_990 ();
 sg13g2_decap_8 FILLER_195_997 ();
 sg13g2_decap_8 FILLER_195_1004 ();
 sg13g2_decap_8 FILLER_195_1011 ();
 sg13g2_decap_8 FILLER_195_1018 ();
 sg13g2_decap_8 FILLER_195_1025 ();
 sg13g2_decap_8 FILLER_195_1032 ();
 sg13g2_decap_8 FILLER_195_1039 ();
 sg13g2_decap_8 FILLER_195_1046 ();
 sg13g2_decap_8 FILLER_195_1053 ();
 sg13g2_decap_8 FILLER_195_1060 ();
 sg13g2_decap_8 FILLER_195_1067 ();
 sg13g2_decap_8 FILLER_195_1074 ();
 sg13g2_decap_8 FILLER_195_1081 ();
 sg13g2_decap_8 FILLER_195_1088 ();
 sg13g2_decap_8 FILLER_195_1095 ();
 sg13g2_decap_8 FILLER_195_1102 ();
 sg13g2_decap_8 FILLER_195_1109 ();
 sg13g2_decap_8 FILLER_195_1116 ();
 sg13g2_decap_8 FILLER_195_1123 ();
 sg13g2_decap_8 FILLER_195_1130 ();
 sg13g2_decap_8 FILLER_195_1137 ();
 sg13g2_decap_8 FILLER_195_1144 ();
 sg13g2_decap_8 FILLER_195_1151 ();
 sg13g2_decap_8 FILLER_195_1158 ();
 sg13g2_decap_8 FILLER_195_1165 ();
 sg13g2_decap_8 FILLER_195_1172 ();
 sg13g2_decap_8 FILLER_195_1179 ();
 sg13g2_decap_8 FILLER_195_1186 ();
 sg13g2_decap_8 FILLER_195_1193 ();
 sg13g2_decap_8 FILLER_195_1200 ();
 sg13g2_decap_8 FILLER_195_1207 ();
 sg13g2_decap_8 FILLER_195_1214 ();
 sg13g2_decap_8 FILLER_195_1221 ();
 sg13g2_decap_8 FILLER_195_1228 ();
 sg13g2_decap_8 FILLER_195_1235 ();
 sg13g2_decap_8 FILLER_195_1242 ();
 sg13g2_decap_8 FILLER_195_1249 ();
 sg13g2_decap_8 FILLER_195_1256 ();
 sg13g2_decap_8 FILLER_195_1263 ();
 sg13g2_decap_8 FILLER_195_1270 ();
 sg13g2_decap_8 FILLER_195_1277 ();
 sg13g2_decap_8 FILLER_195_1284 ();
 sg13g2_decap_8 FILLER_195_1291 ();
 sg13g2_decap_8 FILLER_195_1298 ();
 sg13g2_decap_8 FILLER_195_1305 ();
 sg13g2_decap_8 FILLER_195_1312 ();
 sg13g2_decap_8 FILLER_195_1319 ();
 sg13g2_decap_8 FILLER_195_1326 ();
 sg13g2_decap_8 FILLER_195_1333 ();
 sg13g2_decap_8 FILLER_195_1340 ();
 sg13g2_decap_8 FILLER_195_1347 ();
 sg13g2_decap_8 FILLER_195_1354 ();
 sg13g2_decap_8 FILLER_195_1361 ();
 sg13g2_decap_8 FILLER_195_1368 ();
 sg13g2_decap_8 FILLER_195_1375 ();
 sg13g2_decap_8 FILLER_195_1382 ();
 sg13g2_decap_8 FILLER_195_1389 ();
 sg13g2_decap_8 FILLER_195_1396 ();
 sg13g2_decap_8 FILLER_195_1403 ();
 sg13g2_decap_8 FILLER_195_1410 ();
 sg13g2_decap_8 FILLER_195_1417 ();
 sg13g2_decap_8 FILLER_195_1424 ();
 sg13g2_decap_8 FILLER_195_1431 ();
 sg13g2_decap_8 FILLER_195_1438 ();
 sg13g2_decap_8 FILLER_195_1445 ();
 sg13g2_decap_8 FILLER_195_1452 ();
 sg13g2_decap_8 FILLER_195_1459 ();
 sg13g2_decap_8 FILLER_195_1466 ();
 sg13g2_decap_8 FILLER_195_1473 ();
 sg13g2_decap_8 FILLER_195_1480 ();
 sg13g2_decap_8 FILLER_195_1487 ();
 sg13g2_decap_8 FILLER_195_1494 ();
 sg13g2_decap_8 FILLER_195_1501 ();
 sg13g2_decap_8 FILLER_195_1508 ();
 sg13g2_decap_8 FILLER_195_1515 ();
 sg13g2_decap_8 FILLER_195_1522 ();
 sg13g2_decap_8 FILLER_195_1529 ();
 sg13g2_decap_8 FILLER_195_1536 ();
 sg13g2_decap_8 FILLER_195_1543 ();
 sg13g2_decap_8 FILLER_195_1550 ();
 sg13g2_decap_8 FILLER_195_1557 ();
 sg13g2_decap_8 FILLER_195_1564 ();
 sg13g2_decap_8 FILLER_195_1571 ();
 sg13g2_decap_8 FILLER_195_1578 ();
 sg13g2_decap_8 FILLER_195_1585 ();
 sg13g2_decap_8 FILLER_195_1592 ();
 sg13g2_decap_8 FILLER_195_1599 ();
 sg13g2_decap_8 FILLER_195_1606 ();
 sg13g2_decap_8 FILLER_195_1613 ();
 sg13g2_decap_4 FILLER_195_1620 ();
 sg13g2_fill_1 FILLER_195_1624 ();
 sg13g2_decap_8 FILLER_196_0 ();
 sg13g2_decap_8 FILLER_196_7 ();
 sg13g2_decap_8 FILLER_196_14 ();
 sg13g2_decap_8 FILLER_196_21 ();
 sg13g2_decap_8 FILLER_196_28 ();
 sg13g2_decap_8 FILLER_196_35 ();
 sg13g2_decap_8 FILLER_196_42 ();
 sg13g2_decap_8 FILLER_196_49 ();
 sg13g2_decap_8 FILLER_196_56 ();
 sg13g2_decap_8 FILLER_196_63 ();
 sg13g2_decap_8 FILLER_196_70 ();
 sg13g2_decap_8 FILLER_196_77 ();
 sg13g2_decap_8 FILLER_196_84 ();
 sg13g2_decap_8 FILLER_196_91 ();
 sg13g2_decap_8 FILLER_196_98 ();
 sg13g2_decap_8 FILLER_196_105 ();
 sg13g2_decap_8 FILLER_196_112 ();
 sg13g2_decap_8 FILLER_196_119 ();
 sg13g2_decap_8 FILLER_196_126 ();
 sg13g2_decap_8 FILLER_196_133 ();
 sg13g2_decap_8 FILLER_196_140 ();
 sg13g2_decap_8 FILLER_196_147 ();
 sg13g2_decap_8 FILLER_196_154 ();
 sg13g2_decap_8 FILLER_196_161 ();
 sg13g2_decap_8 FILLER_196_168 ();
 sg13g2_decap_8 FILLER_196_175 ();
 sg13g2_decap_8 FILLER_196_182 ();
 sg13g2_decap_8 FILLER_196_189 ();
 sg13g2_decap_8 FILLER_196_196 ();
 sg13g2_decap_8 FILLER_196_203 ();
 sg13g2_decap_8 FILLER_196_210 ();
 sg13g2_decap_8 FILLER_196_217 ();
 sg13g2_decap_8 FILLER_196_224 ();
 sg13g2_decap_8 FILLER_196_231 ();
 sg13g2_decap_8 FILLER_196_238 ();
 sg13g2_decap_8 FILLER_196_245 ();
 sg13g2_decap_8 FILLER_196_252 ();
 sg13g2_decap_8 FILLER_196_259 ();
 sg13g2_decap_8 FILLER_196_266 ();
 sg13g2_decap_8 FILLER_196_273 ();
 sg13g2_decap_8 FILLER_196_280 ();
 sg13g2_decap_8 FILLER_196_287 ();
 sg13g2_decap_8 FILLER_196_294 ();
 sg13g2_decap_8 FILLER_196_301 ();
 sg13g2_decap_8 FILLER_196_308 ();
 sg13g2_decap_8 FILLER_196_315 ();
 sg13g2_decap_8 FILLER_196_322 ();
 sg13g2_decap_4 FILLER_196_329 ();
 sg13g2_fill_2 FILLER_196_333 ();
 sg13g2_decap_8 FILLER_196_343 ();
 sg13g2_decap_8 FILLER_196_350 ();
 sg13g2_decap_8 FILLER_196_365 ();
 sg13g2_fill_2 FILLER_196_372 ();
 sg13g2_decap_8 FILLER_196_381 ();
 sg13g2_decap_8 FILLER_196_388 ();
 sg13g2_decap_8 FILLER_196_395 ();
 sg13g2_decap_8 FILLER_196_402 ();
 sg13g2_decap_8 FILLER_196_409 ();
 sg13g2_decap_8 FILLER_196_416 ();
 sg13g2_decap_8 FILLER_196_423 ();
 sg13g2_decap_8 FILLER_196_435 ();
 sg13g2_decap_8 FILLER_196_450 ();
 sg13g2_decap_8 FILLER_196_457 ();
 sg13g2_fill_2 FILLER_196_464 ();
 sg13g2_fill_1 FILLER_196_466 ();
 sg13g2_decap_8 FILLER_196_475 ();
 sg13g2_decap_8 FILLER_196_482 ();
 sg13g2_fill_1 FILLER_196_489 ();
 sg13g2_decap_4 FILLER_196_500 ();
 sg13g2_fill_2 FILLER_196_504 ();
 sg13g2_decap_4 FILLER_196_521 ();
 sg13g2_decap_4 FILLER_196_532 ();
 sg13g2_fill_1 FILLER_196_536 ();
 sg13g2_fill_1 FILLER_196_542 ();
 sg13g2_fill_2 FILLER_196_551 ();
 sg13g2_fill_2 FILLER_196_558 ();
 sg13g2_fill_1 FILLER_196_560 ();
 sg13g2_decap_8 FILLER_196_574 ();
 sg13g2_fill_2 FILLER_196_586 ();
 sg13g2_fill_1 FILLER_196_588 ();
 sg13g2_fill_2 FILLER_196_594 ();
 sg13g2_fill_1 FILLER_196_619 ();
 sg13g2_fill_2 FILLER_196_678 ();
 sg13g2_fill_2 FILLER_196_690 ();
 sg13g2_decap_4 FILLER_196_700 ();
 sg13g2_fill_2 FILLER_196_704 ();
 sg13g2_decap_8 FILLER_196_720 ();
 sg13g2_decap_8 FILLER_196_727 ();
 sg13g2_decap_8 FILLER_196_734 ();
 sg13g2_decap_8 FILLER_196_741 ();
 sg13g2_decap_8 FILLER_196_748 ();
 sg13g2_decap_8 FILLER_196_755 ();
 sg13g2_decap_8 FILLER_196_762 ();
 sg13g2_decap_8 FILLER_196_769 ();
 sg13g2_decap_8 FILLER_196_776 ();
 sg13g2_decap_8 FILLER_196_783 ();
 sg13g2_decap_8 FILLER_196_790 ();
 sg13g2_decap_8 FILLER_196_797 ();
 sg13g2_decap_8 FILLER_196_804 ();
 sg13g2_decap_8 FILLER_196_811 ();
 sg13g2_decap_8 FILLER_196_818 ();
 sg13g2_decap_8 FILLER_196_825 ();
 sg13g2_decap_8 FILLER_196_832 ();
 sg13g2_decap_8 FILLER_196_839 ();
 sg13g2_decap_4 FILLER_196_846 ();
 sg13g2_fill_1 FILLER_196_850 ();
 sg13g2_decap_8 FILLER_196_855 ();
 sg13g2_decap_8 FILLER_196_862 ();
 sg13g2_decap_4 FILLER_196_869 ();
 sg13g2_decap_4 FILLER_196_882 ();
 sg13g2_decap_8 FILLER_196_898 ();
 sg13g2_fill_2 FILLER_196_905 ();
 sg13g2_decap_8 FILLER_196_919 ();
 sg13g2_decap_8 FILLER_196_926 ();
 sg13g2_decap_8 FILLER_196_933 ();
 sg13g2_decap_8 FILLER_196_940 ();
 sg13g2_decap_8 FILLER_196_947 ();
 sg13g2_decap_8 FILLER_196_954 ();
 sg13g2_decap_8 FILLER_196_961 ();
 sg13g2_decap_8 FILLER_196_968 ();
 sg13g2_decap_8 FILLER_196_975 ();
 sg13g2_decap_8 FILLER_196_982 ();
 sg13g2_decap_8 FILLER_196_989 ();
 sg13g2_decap_8 FILLER_196_996 ();
 sg13g2_decap_8 FILLER_196_1003 ();
 sg13g2_decap_8 FILLER_196_1010 ();
 sg13g2_decap_8 FILLER_196_1017 ();
 sg13g2_decap_8 FILLER_196_1024 ();
 sg13g2_decap_8 FILLER_196_1031 ();
 sg13g2_decap_8 FILLER_196_1038 ();
 sg13g2_decap_8 FILLER_196_1045 ();
 sg13g2_decap_8 FILLER_196_1052 ();
 sg13g2_decap_8 FILLER_196_1059 ();
 sg13g2_decap_8 FILLER_196_1066 ();
 sg13g2_decap_8 FILLER_196_1073 ();
 sg13g2_decap_8 FILLER_196_1080 ();
 sg13g2_decap_8 FILLER_196_1087 ();
 sg13g2_decap_8 FILLER_196_1094 ();
 sg13g2_decap_8 FILLER_196_1101 ();
 sg13g2_decap_8 FILLER_196_1108 ();
 sg13g2_decap_8 FILLER_196_1115 ();
 sg13g2_decap_8 FILLER_196_1122 ();
 sg13g2_decap_8 FILLER_196_1129 ();
 sg13g2_decap_8 FILLER_196_1136 ();
 sg13g2_decap_8 FILLER_196_1143 ();
 sg13g2_decap_8 FILLER_196_1150 ();
 sg13g2_decap_8 FILLER_196_1157 ();
 sg13g2_decap_8 FILLER_196_1164 ();
 sg13g2_decap_8 FILLER_196_1171 ();
 sg13g2_decap_8 FILLER_196_1178 ();
 sg13g2_decap_8 FILLER_196_1185 ();
 sg13g2_decap_8 FILLER_196_1192 ();
 sg13g2_decap_8 FILLER_196_1199 ();
 sg13g2_decap_8 FILLER_196_1206 ();
 sg13g2_decap_8 FILLER_196_1213 ();
 sg13g2_decap_8 FILLER_196_1220 ();
 sg13g2_decap_8 FILLER_196_1227 ();
 sg13g2_decap_8 FILLER_196_1234 ();
 sg13g2_decap_8 FILLER_196_1241 ();
 sg13g2_decap_8 FILLER_196_1248 ();
 sg13g2_decap_8 FILLER_196_1255 ();
 sg13g2_decap_8 FILLER_196_1262 ();
 sg13g2_decap_8 FILLER_196_1269 ();
 sg13g2_decap_8 FILLER_196_1276 ();
 sg13g2_decap_8 FILLER_196_1283 ();
 sg13g2_decap_8 FILLER_196_1290 ();
 sg13g2_decap_8 FILLER_196_1297 ();
 sg13g2_decap_8 FILLER_196_1304 ();
 sg13g2_decap_8 FILLER_196_1311 ();
 sg13g2_decap_8 FILLER_196_1318 ();
 sg13g2_decap_8 FILLER_196_1325 ();
 sg13g2_decap_8 FILLER_196_1332 ();
 sg13g2_decap_8 FILLER_196_1339 ();
 sg13g2_decap_8 FILLER_196_1346 ();
 sg13g2_decap_8 FILLER_196_1353 ();
 sg13g2_decap_8 FILLER_196_1360 ();
 sg13g2_decap_8 FILLER_196_1367 ();
 sg13g2_decap_8 FILLER_196_1374 ();
 sg13g2_decap_8 FILLER_196_1381 ();
 sg13g2_decap_8 FILLER_196_1388 ();
 sg13g2_decap_8 FILLER_196_1395 ();
 sg13g2_decap_8 FILLER_196_1402 ();
 sg13g2_decap_8 FILLER_196_1409 ();
 sg13g2_decap_8 FILLER_196_1416 ();
 sg13g2_decap_8 FILLER_196_1423 ();
 sg13g2_decap_8 FILLER_196_1430 ();
 sg13g2_decap_8 FILLER_196_1437 ();
 sg13g2_decap_8 FILLER_196_1444 ();
 sg13g2_decap_8 FILLER_196_1451 ();
 sg13g2_decap_8 FILLER_196_1458 ();
 sg13g2_decap_8 FILLER_196_1465 ();
 sg13g2_decap_8 FILLER_196_1472 ();
 sg13g2_decap_8 FILLER_196_1479 ();
 sg13g2_decap_8 FILLER_196_1486 ();
 sg13g2_decap_8 FILLER_196_1493 ();
 sg13g2_decap_8 FILLER_196_1500 ();
 sg13g2_decap_8 FILLER_196_1507 ();
 sg13g2_decap_8 FILLER_196_1514 ();
 sg13g2_decap_8 FILLER_196_1521 ();
 sg13g2_decap_8 FILLER_196_1528 ();
 sg13g2_decap_8 FILLER_196_1535 ();
 sg13g2_decap_8 FILLER_196_1542 ();
 sg13g2_decap_8 FILLER_196_1549 ();
 sg13g2_decap_8 FILLER_196_1556 ();
 sg13g2_decap_8 FILLER_196_1563 ();
 sg13g2_decap_8 FILLER_196_1570 ();
 sg13g2_decap_8 FILLER_196_1577 ();
 sg13g2_decap_8 FILLER_196_1584 ();
 sg13g2_decap_8 FILLER_196_1591 ();
 sg13g2_decap_8 FILLER_196_1598 ();
 sg13g2_decap_8 FILLER_196_1605 ();
 sg13g2_decap_8 FILLER_196_1612 ();
 sg13g2_decap_4 FILLER_196_1619 ();
 sg13g2_fill_2 FILLER_196_1623 ();
 sg13g2_decap_8 FILLER_197_0 ();
 sg13g2_decap_8 FILLER_197_7 ();
 sg13g2_decap_8 FILLER_197_14 ();
 sg13g2_decap_8 FILLER_197_21 ();
 sg13g2_decap_8 FILLER_197_28 ();
 sg13g2_decap_8 FILLER_197_35 ();
 sg13g2_decap_8 FILLER_197_42 ();
 sg13g2_decap_8 FILLER_197_49 ();
 sg13g2_decap_8 FILLER_197_56 ();
 sg13g2_decap_8 FILLER_197_63 ();
 sg13g2_decap_8 FILLER_197_70 ();
 sg13g2_decap_8 FILLER_197_77 ();
 sg13g2_decap_8 FILLER_197_84 ();
 sg13g2_decap_8 FILLER_197_91 ();
 sg13g2_decap_8 FILLER_197_98 ();
 sg13g2_decap_8 FILLER_197_105 ();
 sg13g2_decap_8 FILLER_197_112 ();
 sg13g2_decap_8 FILLER_197_119 ();
 sg13g2_decap_8 FILLER_197_126 ();
 sg13g2_decap_8 FILLER_197_133 ();
 sg13g2_decap_8 FILLER_197_140 ();
 sg13g2_decap_8 FILLER_197_147 ();
 sg13g2_decap_8 FILLER_197_154 ();
 sg13g2_decap_8 FILLER_197_161 ();
 sg13g2_decap_8 FILLER_197_168 ();
 sg13g2_decap_8 FILLER_197_175 ();
 sg13g2_decap_8 FILLER_197_182 ();
 sg13g2_decap_8 FILLER_197_189 ();
 sg13g2_decap_8 FILLER_197_196 ();
 sg13g2_decap_8 FILLER_197_203 ();
 sg13g2_decap_8 FILLER_197_210 ();
 sg13g2_decap_8 FILLER_197_217 ();
 sg13g2_decap_8 FILLER_197_224 ();
 sg13g2_decap_8 FILLER_197_231 ();
 sg13g2_decap_8 FILLER_197_238 ();
 sg13g2_decap_8 FILLER_197_245 ();
 sg13g2_decap_8 FILLER_197_252 ();
 sg13g2_decap_8 FILLER_197_259 ();
 sg13g2_decap_8 FILLER_197_266 ();
 sg13g2_decap_8 FILLER_197_273 ();
 sg13g2_decap_8 FILLER_197_280 ();
 sg13g2_decap_8 FILLER_197_287 ();
 sg13g2_decap_8 FILLER_197_294 ();
 sg13g2_decap_8 FILLER_197_301 ();
 sg13g2_decap_8 FILLER_197_308 ();
 sg13g2_decap_8 FILLER_197_315 ();
 sg13g2_decap_8 FILLER_197_322 ();
 sg13g2_decap_4 FILLER_197_329 ();
 sg13g2_decap_4 FILLER_197_341 ();
 sg13g2_fill_1 FILLER_197_345 ();
 sg13g2_decap_8 FILLER_197_376 ();
 sg13g2_decap_8 FILLER_197_383 ();
 sg13g2_decap_8 FILLER_197_390 ();
 sg13g2_decap_4 FILLER_197_397 ();
 sg13g2_fill_2 FILLER_197_413 ();
 sg13g2_fill_1 FILLER_197_415 ();
 sg13g2_decap_4 FILLER_197_420 ();
 sg13g2_fill_2 FILLER_197_424 ();
 sg13g2_fill_2 FILLER_197_464 ();
 sg13g2_fill_1 FILLER_197_466 ();
 sg13g2_fill_2 FILLER_197_502 ();
 sg13g2_decap_8 FILLER_197_523 ();
 sg13g2_decap_8 FILLER_197_530 ();
 sg13g2_fill_1 FILLER_197_537 ();
 sg13g2_decap_4 FILLER_197_550 ();
 sg13g2_decap_8 FILLER_197_559 ();
 sg13g2_decap_8 FILLER_197_566 ();
 sg13g2_fill_2 FILLER_197_573 ();
 sg13g2_fill_1 FILLER_197_575 ();
 sg13g2_decap_4 FILLER_197_580 ();
 sg13g2_fill_1 FILLER_197_584 ();
 sg13g2_decap_8 FILLER_197_590 ();
 sg13g2_fill_2 FILLER_197_597 ();
 sg13g2_fill_2 FILLER_197_604 ();
 sg13g2_decap_4 FILLER_197_622 ();
 sg13g2_fill_2 FILLER_197_648 ();
 sg13g2_fill_1 FILLER_197_650 ();
 sg13g2_decap_8 FILLER_197_659 ();
 sg13g2_decap_8 FILLER_197_666 ();
 sg13g2_decap_8 FILLER_197_673 ();
 sg13g2_decap_8 FILLER_197_680 ();
 sg13g2_decap_8 FILLER_197_687 ();
 sg13g2_decap_8 FILLER_197_694 ();
 sg13g2_fill_1 FILLER_197_701 ();
 sg13g2_decap_8 FILLER_197_706 ();
 sg13g2_decap_8 FILLER_197_713 ();
 sg13g2_decap_8 FILLER_197_720 ();
 sg13g2_decap_8 FILLER_197_727 ();
 sg13g2_decap_8 FILLER_197_734 ();
 sg13g2_decap_8 FILLER_197_741 ();
 sg13g2_decap_8 FILLER_197_748 ();
 sg13g2_decap_8 FILLER_197_755 ();
 sg13g2_decap_8 FILLER_197_762 ();
 sg13g2_decap_8 FILLER_197_769 ();
 sg13g2_decap_8 FILLER_197_776 ();
 sg13g2_decap_8 FILLER_197_783 ();
 sg13g2_decap_8 FILLER_197_790 ();
 sg13g2_decap_8 FILLER_197_797 ();
 sg13g2_decap_8 FILLER_197_804 ();
 sg13g2_decap_8 FILLER_197_811 ();
 sg13g2_decap_8 FILLER_197_818 ();
 sg13g2_decap_8 FILLER_197_825 ();
 sg13g2_decap_8 FILLER_197_832 ();
 sg13g2_fill_2 FILLER_197_839 ();
 sg13g2_decap_8 FILLER_197_879 ();
 sg13g2_fill_2 FILLER_197_886 ();
 sg13g2_fill_1 FILLER_197_888 ();
 sg13g2_decap_8 FILLER_197_901 ();
 sg13g2_fill_2 FILLER_197_908 ();
 sg13g2_fill_1 FILLER_197_910 ();
 sg13g2_decap_4 FILLER_197_915 ();
 sg13g2_decap_8 FILLER_197_948 ();
 sg13g2_decap_8 FILLER_197_955 ();
 sg13g2_decap_8 FILLER_197_962 ();
 sg13g2_decap_8 FILLER_197_969 ();
 sg13g2_decap_8 FILLER_197_976 ();
 sg13g2_decap_8 FILLER_197_983 ();
 sg13g2_decap_8 FILLER_197_990 ();
 sg13g2_decap_8 FILLER_197_997 ();
 sg13g2_decap_8 FILLER_197_1004 ();
 sg13g2_decap_8 FILLER_197_1011 ();
 sg13g2_decap_8 FILLER_197_1018 ();
 sg13g2_decap_8 FILLER_197_1025 ();
 sg13g2_decap_8 FILLER_197_1032 ();
 sg13g2_decap_8 FILLER_197_1039 ();
 sg13g2_decap_8 FILLER_197_1046 ();
 sg13g2_decap_8 FILLER_197_1053 ();
 sg13g2_decap_8 FILLER_197_1060 ();
 sg13g2_decap_8 FILLER_197_1067 ();
 sg13g2_decap_8 FILLER_197_1074 ();
 sg13g2_decap_8 FILLER_197_1081 ();
 sg13g2_decap_8 FILLER_197_1088 ();
 sg13g2_decap_8 FILLER_197_1095 ();
 sg13g2_decap_8 FILLER_197_1102 ();
 sg13g2_decap_8 FILLER_197_1109 ();
 sg13g2_decap_8 FILLER_197_1116 ();
 sg13g2_decap_8 FILLER_197_1123 ();
 sg13g2_decap_8 FILLER_197_1130 ();
 sg13g2_decap_8 FILLER_197_1137 ();
 sg13g2_decap_8 FILLER_197_1144 ();
 sg13g2_decap_8 FILLER_197_1151 ();
 sg13g2_decap_8 FILLER_197_1158 ();
 sg13g2_decap_8 FILLER_197_1165 ();
 sg13g2_decap_8 FILLER_197_1172 ();
 sg13g2_decap_8 FILLER_197_1179 ();
 sg13g2_decap_8 FILLER_197_1186 ();
 sg13g2_decap_8 FILLER_197_1193 ();
 sg13g2_decap_8 FILLER_197_1200 ();
 sg13g2_decap_8 FILLER_197_1207 ();
 sg13g2_decap_8 FILLER_197_1214 ();
 sg13g2_decap_8 FILLER_197_1221 ();
 sg13g2_decap_8 FILLER_197_1228 ();
 sg13g2_decap_8 FILLER_197_1235 ();
 sg13g2_decap_8 FILLER_197_1242 ();
 sg13g2_decap_8 FILLER_197_1249 ();
 sg13g2_decap_8 FILLER_197_1256 ();
 sg13g2_decap_8 FILLER_197_1263 ();
 sg13g2_decap_8 FILLER_197_1270 ();
 sg13g2_decap_8 FILLER_197_1277 ();
 sg13g2_decap_8 FILLER_197_1284 ();
 sg13g2_decap_8 FILLER_197_1291 ();
 sg13g2_decap_8 FILLER_197_1298 ();
 sg13g2_decap_8 FILLER_197_1305 ();
 sg13g2_decap_8 FILLER_197_1312 ();
 sg13g2_decap_8 FILLER_197_1319 ();
 sg13g2_decap_8 FILLER_197_1326 ();
 sg13g2_decap_8 FILLER_197_1333 ();
 sg13g2_decap_8 FILLER_197_1340 ();
 sg13g2_decap_8 FILLER_197_1347 ();
 sg13g2_decap_8 FILLER_197_1354 ();
 sg13g2_decap_8 FILLER_197_1361 ();
 sg13g2_decap_8 FILLER_197_1368 ();
 sg13g2_decap_8 FILLER_197_1375 ();
 sg13g2_decap_8 FILLER_197_1382 ();
 sg13g2_decap_8 FILLER_197_1389 ();
 sg13g2_decap_8 FILLER_197_1396 ();
 sg13g2_decap_8 FILLER_197_1403 ();
 sg13g2_decap_8 FILLER_197_1410 ();
 sg13g2_decap_8 FILLER_197_1417 ();
 sg13g2_decap_8 FILLER_197_1424 ();
 sg13g2_decap_8 FILLER_197_1431 ();
 sg13g2_decap_8 FILLER_197_1438 ();
 sg13g2_decap_8 FILLER_197_1445 ();
 sg13g2_decap_8 FILLER_197_1452 ();
 sg13g2_decap_8 FILLER_197_1459 ();
 sg13g2_decap_8 FILLER_197_1466 ();
 sg13g2_decap_8 FILLER_197_1473 ();
 sg13g2_decap_8 FILLER_197_1480 ();
 sg13g2_decap_8 FILLER_197_1487 ();
 sg13g2_decap_8 FILLER_197_1494 ();
 sg13g2_decap_8 FILLER_197_1501 ();
 sg13g2_decap_8 FILLER_197_1508 ();
 sg13g2_decap_8 FILLER_197_1515 ();
 sg13g2_decap_8 FILLER_197_1522 ();
 sg13g2_decap_8 FILLER_197_1529 ();
 sg13g2_decap_8 FILLER_197_1536 ();
 sg13g2_decap_8 FILLER_197_1543 ();
 sg13g2_decap_8 FILLER_197_1550 ();
 sg13g2_decap_8 FILLER_197_1557 ();
 sg13g2_decap_8 FILLER_197_1564 ();
 sg13g2_decap_8 FILLER_197_1571 ();
 sg13g2_decap_8 FILLER_197_1578 ();
 sg13g2_decap_8 FILLER_197_1585 ();
 sg13g2_decap_8 FILLER_197_1592 ();
 sg13g2_decap_8 FILLER_197_1599 ();
 sg13g2_decap_8 FILLER_197_1606 ();
 sg13g2_decap_8 FILLER_197_1613 ();
 sg13g2_decap_4 FILLER_197_1620 ();
 sg13g2_fill_1 FILLER_197_1624 ();
 sg13g2_decap_8 FILLER_198_0 ();
 sg13g2_decap_8 FILLER_198_7 ();
 sg13g2_decap_8 FILLER_198_14 ();
 sg13g2_decap_8 FILLER_198_21 ();
 sg13g2_decap_8 FILLER_198_28 ();
 sg13g2_decap_8 FILLER_198_35 ();
 sg13g2_decap_8 FILLER_198_42 ();
 sg13g2_decap_8 FILLER_198_49 ();
 sg13g2_decap_8 FILLER_198_56 ();
 sg13g2_decap_8 FILLER_198_63 ();
 sg13g2_decap_8 FILLER_198_70 ();
 sg13g2_decap_8 FILLER_198_77 ();
 sg13g2_decap_8 FILLER_198_84 ();
 sg13g2_decap_8 FILLER_198_91 ();
 sg13g2_decap_8 FILLER_198_98 ();
 sg13g2_decap_8 FILLER_198_105 ();
 sg13g2_decap_8 FILLER_198_112 ();
 sg13g2_decap_8 FILLER_198_119 ();
 sg13g2_decap_8 FILLER_198_126 ();
 sg13g2_decap_8 FILLER_198_133 ();
 sg13g2_decap_8 FILLER_198_140 ();
 sg13g2_decap_8 FILLER_198_147 ();
 sg13g2_decap_8 FILLER_198_154 ();
 sg13g2_decap_8 FILLER_198_161 ();
 sg13g2_decap_8 FILLER_198_168 ();
 sg13g2_decap_8 FILLER_198_175 ();
 sg13g2_decap_8 FILLER_198_182 ();
 sg13g2_decap_8 FILLER_198_189 ();
 sg13g2_decap_8 FILLER_198_196 ();
 sg13g2_decap_8 FILLER_198_203 ();
 sg13g2_decap_8 FILLER_198_210 ();
 sg13g2_decap_8 FILLER_198_217 ();
 sg13g2_decap_8 FILLER_198_224 ();
 sg13g2_decap_8 FILLER_198_231 ();
 sg13g2_decap_8 FILLER_198_238 ();
 sg13g2_decap_8 FILLER_198_245 ();
 sg13g2_decap_8 FILLER_198_252 ();
 sg13g2_decap_8 FILLER_198_259 ();
 sg13g2_decap_8 FILLER_198_266 ();
 sg13g2_decap_8 FILLER_198_273 ();
 sg13g2_decap_8 FILLER_198_280 ();
 sg13g2_decap_8 FILLER_198_287 ();
 sg13g2_decap_8 FILLER_198_294 ();
 sg13g2_decap_8 FILLER_198_301 ();
 sg13g2_decap_8 FILLER_198_308 ();
 sg13g2_decap_8 FILLER_198_315 ();
 sg13g2_fill_2 FILLER_198_322 ();
 sg13g2_fill_1 FILLER_198_324 ();
 sg13g2_decap_8 FILLER_198_351 ();
 sg13g2_decap_8 FILLER_198_362 ();
 sg13g2_decap_8 FILLER_198_369 ();
 sg13g2_fill_2 FILLER_198_376 ();
 sg13g2_fill_1 FILLER_198_378 ();
 sg13g2_decap_4 FILLER_198_391 ();
 sg13g2_decap_4 FILLER_198_400 ();
 sg13g2_fill_1 FILLER_198_404 ();
 sg13g2_decap_8 FILLER_198_460 ();
 sg13g2_decap_4 FILLER_198_467 ();
 sg13g2_fill_1 FILLER_198_471 ();
 sg13g2_decap_8 FILLER_198_481 ();
 sg13g2_decap_8 FILLER_198_491 ();
 sg13g2_decap_8 FILLER_198_506 ();
 sg13g2_decap_8 FILLER_198_513 ();
 sg13g2_decap_8 FILLER_198_520 ();
 sg13g2_decap_8 FILLER_198_527 ();
 sg13g2_decap_8 FILLER_198_534 ();
 sg13g2_decap_8 FILLER_198_541 ();
 sg13g2_decap_8 FILLER_198_548 ();
 sg13g2_decap_8 FILLER_198_555 ();
 sg13g2_decap_8 FILLER_198_575 ();
 sg13g2_decap_4 FILLER_198_582 ();
 sg13g2_decap_8 FILLER_198_590 ();
 sg13g2_decap_8 FILLER_198_597 ();
 sg13g2_decap_8 FILLER_198_604 ();
 sg13g2_decap_8 FILLER_198_611 ();
 sg13g2_decap_8 FILLER_198_618 ();
 sg13g2_decap_8 FILLER_198_625 ();
 sg13g2_fill_2 FILLER_198_632 ();
 sg13g2_fill_1 FILLER_198_634 ();
 sg13g2_decap_8 FILLER_198_648 ();
 sg13g2_fill_2 FILLER_198_655 ();
 sg13g2_fill_2 FILLER_198_665 ();
 sg13g2_decap_4 FILLER_198_676 ();
 sg13g2_fill_2 FILLER_198_680 ();
 sg13g2_fill_1 FILLER_198_686 ();
 sg13g2_fill_1 FILLER_198_692 ();
 sg13g2_decap_8 FILLER_198_719 ();
 sg13g2_decap_8 FILLER_198_726 ();
 sg13g2_decap_8 FILLER_198_733 ();
 sg13g2_decap_8 FILLER_198_740 ();
 sg13g2_decap_8 FILLER_198_747 ();
 sg13g2_decap_8 FILLER_198_754 ();
 sg13g2_decap_8 FILLER_198_761 ();
 sg13g2_decap_8 FILLER_198_768 ();
 sg13g2_decap_8 FILLER_198_775 ();
 sg13g2_decap_8 FILLER_198_782 ();
 sg13g2_decap_8 FILLER_198_789 ();
 sg13g2_decap_8 FILLER_198_796 ();
 sg13g2_decap_8 FILLER_198_803 ();
 sg13g2_decap_8 FILLER_198_810 ();
 sg13g2_decap_8 FILLER_198_817 ();
 sg13g2_decap_8 FILLER_198_824 ();
 sg13g2_decap_8 FILLER_198_831 ();
 sg13g2_decap_8 FILLER_198_838 ();
 sg13g2_decap_8 FILLER_198_845 ();
 sg13g2_decap_8 FILLER_198_852 ();
 sg13g2_decap_8 FILLER_198_859 ();
 sg13g2_decap_4 FILLER_198_866 ();
 sg13g2_fill_2 FILLER_198_870 ();
 sg13g2_decap_8 FILLER_198_940 ();
 sg13g2_decap_8 FILLER_198_947 ();
 sg13g2_decap_8 FILLER_198_954 ();
 sg13g2_decap_8 FILLER_198_961 ();
 sg13g2_decap_8 FILLER_198_968 ();
 sg13g2_decap_8 FILLER_198_975 ();
 sg13g2_decap_8 FILLER_198_982 ();
 sg13g2_decap_8 FILLER_198_989 ();
 sg13g2_decap_8 FILLER_198_996 ();
 sg13g2_decap_8 FILLER_198_1003 ();
 sg13g2_decap_8 FILLER_198_1010 ();
 sg13g2_decap_8 FILLER_198_1017 ();
 sg13g2_decap_8 FILLER_198_1024 ();
 sg13g2_decap_8 FILLER_198_1031 ();
 sg13g2_decap_8 FILLER_198_1038 ();
 sg13g2_decap_8 FILLER_198_1045 ();
 sg13g2_decap_8 FILLER_198_1052 ();
 sg13g2_decap_8 FILLER_198_1059 ();
 sg13g2_decap_8 FILLER_198_1066 ();
 sg13g2_decap_8 FILLER_198_1073 ();
 sg13g2_decap_8 FILLER_198_1080 ();
 sg13g2_decap_8 FILLER_198_1087 ();
 sg13g2_decap_8 FILLER_198_1094 ();
 sg13g2_decap_8 FILLER_198_1101 ();
 sg13g2_decap_8 FILLER_198_1108 ();
 sg13g2_decap_8 FILLER_198_1115 ();
 sg13g2_decap_8 FILLER_198_1122 ();
 sg13g2_decap_8 FILLER_198_1129 ();
 sg13g2_decap_8 FILLER_198_1136 ();
 sg13g2_decap_8 FILLER_198_1143 ();
 sg13g2_decap_8 FILLER_198_1150 ();
 sg13g2_decap_8 FILLER_198_1157 ();
 sg13g2_decap_8 FILLER_198_1164 ();
 sg13g2_decap_8 FILLER_198_1171 ();
 sg13g2_decap_8 FILLER_198_1178 ();
 sg13g2_decap_8 FILLER_198_1185 ();
 sg13g2_decap_8 FILLER_198_1192 ();
 sg13g2_decap_8 FILLER_198_1199 ();
 sg13g2_decap_8 FILLER_198_1206 ();
 sg13g2_decap_8 FILLER_198_1213 ();
 sg13g2_decap_8 FILLER_198_1220 ();
 sg13g2_decap_8 FILLER_198_1227 ();
 sg13g2_decap_8 FILLER_198_1234 ();
 sg13g2_decap_8 FILLER_198_1241 ();
 sg13g2_decap_8 FILLER_198_1248 ();
 sg13g2_decap_8 FILLER_198_1255 ();
 sg13g2_decap_8 FILLER_198_1262 ();
 sg13g2_decap_8 FILLER_198_1269 ();
 sg13g2_decap_8 FILLER_198_1276 ();
 sg13g2_decap_8 FILLER_198_1283 ();
 sg13g2_decap_8 FILLER_198_1290 ();
 sg13g2_decap_8 FILLER_198_1297 ();
 sg13g2_decap_8 FILLER_198_1304 ();
 sg13g2_decap_8 FILLER_198_1311 ();
 sg13g2_decap_8 FILLER_198_1318 ();
 sg13g2_decap_8 FILLER_198_1325 ();
 sg13g2_decap_8 FILLER_198_1332 ();
 sg13g2_decap_8 FILLER_198_1339 ();
 sg13g2_decap_8 FILLER_198_1346 ();
 sg13g2_decap_8 FILLER_198_1353 ();
 sg13g2_decap_8 FILLER_198_1360 ();
 sg13g2_decap_8 FILLER_198_1367 ();
 sg13g2_decap_8 FILLER_198_1374 ();
 sg13g2_decap_8 FILLER_198_1381 ();
 sg13g2_decap_8 FILLER_198_1388 ();
 sg13g2_decap_8 FILLER_198_1395 ();
 sg13g2_decap_8 FILLER_198_1402 ();
 sg13g2_decap_8 FILLER_198_1409 ();
 sg13g2_decap_8 FILLER_198_1416 ();
 sg13g2_decap_8 FILLER_198_1423 ();
 sg13g2_decap_8 FILLER_198_1430 ();
 sg13g2_decap_8 FILLER_198_1437 ();
 sg13g2_decap_8 FILLER_198_1444 ();
 sg13g2_decap_8 FILLER_198_1451 ();
 sg13g2_decap_8 FILLER_198_1458 ();
 sg13g2_decap_8 FILLER_198_1465 ();
 sg13g2_decap_8 FILLER_198_1472 ();
 sg13g2_decap_8 FILLER_198_1479 ();
 sg13g2_decap_8 FILLER_198_1486 ();
 sg13g2_decap_8 FILLER_198_1493 ();
 sg13g2_decap_8 FILLER_198_1500 ();
 sg13g2_decap_8 FILLER_198_1507 ();
 sg13g2_decap_8 FILLER_198_1514 ();
 sg13g2_decap_8 FILLER_198_1521 ();
 sg13g2_decap_8 FILLER_198_1528 ();
 sg13g2_decap_8 FILLER_198_1535 ();
 sg13g2_decap_8 FILLER_198_1542 ();
 sg13g2_decap_8 FILLER_198_1549 ();
 sg13g2_decap_8 FILLER_198_1556 ();
 sg13g2_decap_8 FILLER_198_1563 ();
 sg13g2_decap_8 FILLER_198_1570 ();
 sg13g2_decap_8 FILLER_198_1577 ();
 sg13g2_decap_8 FILLER_198_1584 ();
 sg13g2_decap_8 FILLER_198_1591 ();
 sg13g2_decap_8 FILLER_198_1598 ();
 sg13g2_decap_8 FILLER_198_1605 ();
 sg13g2_decap_8 FILLER_198_1612 ();
 sg13g2_decap_4 FILLER_198_1619 ();
 sg13g2_fill_2 FILLER_198_1623 ();
 sg13g2_decap_8 FILLER_199_0 ();
 sg13g2_decap_8 FILLER_199_7 ();
 sg13g2_decap_8 FILLER_199_14 ();
 sg13g2_decap_8 FILLER_199_21 ();
 sg13g2_decap_8 FILLER_199_28 ();
 sg13g2_decap_8 FILLER_199_35 ();
 sg13g2_decap_8 FILLER_199_42 ();
 sg13g2_decap_8 FILLER_199_49 ();
 sg13g2_decap_8 FILLER_199_56 ();
 sg13g2_decap_8 FILLER_199_63 ();
 sg13g2_decap_8 FILLER_199_70 ();
 sg13g2_decap_8 FILLER_199_77 ();
 sg13g2_decap_8 FILLER_199_84 ();
 sg13g2_decap_8 FILLER_199_91 ();
 sg13g2_decap_8 FILLER_199_98 ();
 sg13g2_decap_8 FILLER_199_105 ();
 sg13g2_decap_8 FILLER_199_112 ();
 sg13g2_decap_8 FILLER_199_119 ();
 sg13g2_decap_8 FILLER_199_126 ();
 sg13g2_decap_8 FILLER_199_133 ();
 sg13g2_decap_8 FILLER_199_140 ();
 sg13g2_decap_8 FILLER_199_147 ();
 sg13g2_decap_8 FILLER_199_154 ();
 sg13g2_decap_8 FILLER_199_161 ();
 sg13g2_decap_8 FILLER_199_168 ();
 sg13g2_decap_8 FILLER_199_175 ();
 sg13g2_decap_8 FILLER_199_182 ();
 sg13g2_decap_8 FILLER_199_189 ();
 sg13g2_decap_8 FILLER_199_196 ();
 sg13g2_decap_8 FILLER_199_203 ();
 sg13g2_decap_8 FILLER_199_210 ();
 sg13g2_decap_8 FILLER_199_217 ();
 sg13g2_decap_8 FILLER_199_224 ();
 sg13g2_decap_8 FILLER_199_231 ();
 sg13g2_decap_8 FILLER_199_238 ();
 sg13g2_decap_8 FILLER_199_245 ();
 sg13g2_decap_8 FILLER_199_252 ();
 sg13g2_decap_8 FILLER_199_259 ();
 sg13g2_decap_8 FILLER_199_266 ();
 sg13g2_decap_8 FILLER_199_273 ();
 sg13g2_decap_8 FILLER_199_280 ();
 sg13g2_decap_8 FILLER_199_287 ();
 sg13g2_decap_8 FILLER_199_294 ();
 sg13g2_decap_8 FILLER_199_301 ();
 sg13g2_decap_8 FILLER_199_308 ();
 sg13g2_decap_8 FILLER_199_315 ();
 sg13g2_decap_8 FILLER_199_322 ();
 sg13g2_decap_8 FILLER_199_329 ();
 sg13g2_decap_4 FILLER_199_336 ();
 sg13g2_fill_2 FILLER_199_340 ();
 sg13g2_decap_8 FILLER_199_367 ();
 sg13g2_decap_4 FILLER_199_374 ();
 sg13g2_fill_2 FILLER_199_378 ();
 sg13g2_decap_8 FILLER_199_406 ();
 sg13g2_decap_8 FILLER_199_413 ();
 sg13g2_decap_8 FILLER_199_420 ();
 sg13g2_fill_1 FILLER_199_427 ();
 sg13g2_decap_4 FILLER_199_431 ();
 sg13g2_decap_8 FILLER_199_441 ();
 sg13g2_decap_8 FILLER_199_448 ();
 sg13g2_fill_2 FILLER_199_467 ();
 sg13g2_decap_8 FILLER_199_474 ();
 sg13g2_fill_1 FILLER_199_481 ();
 sg13g2_decap_4 FILLER_199_492 ();
 sg13g2_fill_1 FILLER_199_496 ();
 sg13g2_fill_1 FILLER_199_510 ();
 sg13g2_fill_1 FILLER_199_519 ();
 sg13g2_decap_4 FILLER_199_524 ();
 sg13g2_decap_4 FILLER_199_533 ();
 sg13g2_decap_4 FILLER_199_542 ();
 sg13g2_fill_2 FILLER_199_546 ();
 sg13g2_decap_8 FILLER_199_556 ();
 sg13g2_fill_2 FILLER_199_567 ();
 sg13g2_fill_1 FILLER_199_569 ();
 sg13g2_decap_8 FILLER_199_604 ();
 sg13g2_decap_8 FILLER_199_611 ();
 sg13g2_decap_8 FILLER_199_618 ();
 sg13g2_decap_8 FILLER_199_625 ();
 sg13g2_decap_4 FILLER_199_632 ();
 sg13g2_decap_8 FILLER_199_645 ();
 sg13g2_decap_8 FILLER_199_652 ();
 sg13g2_fill_2 FILLER_199_659 ();
 sg13g2_decap_8 FILLER_199_691 ();
 sg13g2_decap_4 FILLER_199_698 ();
 sg13g2_decap_8 FILLER_199_706 ();
 sg13g2_decap_8 FILLER_199_713 ();
 sg13g2_decap_8 FILLER_199_720 ();
 sg13g2_decap_8 FILLER_199_727 ();
 sg13g2_decap_8 FILLER_199_734 ();
 sg13g2_decap_8 FILLER_199_741 ();
 sg13g2_decap_8 FILLER_199_748 ();
 sg13g2_decap_8 FILLER_199_755 ();
 sg13g2_decap_8 FILLER_199_762 ();
 sg13g2_decap_8 FILLER_199_769 ();
 sg13g2_decap_8 FILLER_199_776 ();
 sg13g2_decap_8 FILLER_199_783 ();
 sg13g2_decap_8 FILLER_199_790 ();
 sg13g2_decap_8 FILLER_199_797 ();
 sg13g2_decap_8 FILLER_199_804 ();
 sg13g2_decap_8 FILLER_199_811 ();
 sg13g2_decap_8 FILLER_199_818 ();
 sg13g2_decap_8 FILLER_199_825 ();
 sg13g2_decap_8 FILLER_199_832 ();
 sg13g2_decap_8 FILLER_199_839 ();
 sg13g2_decap_8 FILLER_199_846 ();
 sg13g2_decap_8 FILLER_199_853 ();
 sg13g2_decap_8 FILLER_199_860 ();
 sg13g2_decap_8 FILLER_199_867 ();
 sg13g2_decap_8 FILLER_199_874 ();
 sg13g2_fill_1 FILLER_199_885 ();
 sg13g2_decap_8 FILLER_199_911 ();
 sg13g2_decap_8 FILLER_199_918 ();
 sg13g2_decap_8 FILLER_199_925 ();
 sg13g2_decap_8 FILLER_199_932 ();
 sg13g2_decap_8 FILLER_199_939 ();
 sg13g2_decap_8 FILLER_199_946 ();
 sg13g2_decap_8 FILLER_199_953 ();
 sg13g2_decap_8 FILLER_199_960 ();
 sg13g2_decap_8 FILLER_199_967 ();
 sg13g2_decap_8 FILLER_199_974 ();
 sg13g2_decap_8 FILLER_199_981 ();
 sg13g2_decap_8 FILLER_199_988 ();
 sg13g2_decap_8 FILLER_199_995 ();
 sg13g2_decap_8 FILLER_199_1002 ();
 sg13g2_decap_8 FILLER_199_1009 ();
 sg13g2_decap_8 FILLER_199_1016 ();
 sg13g2_decap_8 FILLER_199_1023 ();
 sg13g2_decap_8 FILLER_199_1030 ();
 sg13g2_decap_8 FILLER_199_1037 ();
 sg13g2_decap_8 FILLER_199_1044 ();
 sg13g2_decap_8 FILLER_199_1051 ();
 sg13g2_decap_8 FILLER_199_1058 ();
 sg13g2_decap_8 FILLER_199_1065 ();
 sg13g2_decap_8 FILLER_199_1072 ();
 sg13g2_decap_8 FILLER_199_1079 ();
 sg13g2_decap_8 FILLER_199_1086 ();
 sg13g2_decap_8 FILLER_199_1093 ();
 sg13g2_decap_8 FILLER_199_1100 ();
 sg13g2_decap_8 FILLER_199_1107 ();
 sg13g2_decap_8 FILLER_199_1114 ();
 sg13g2_decap_8 FILLER_199_1121 ();
 sg13g2_decap_8 FILLER_199_1128 ();
 sg13g2_decap_8 FILLER_199_1135 ();
 sg13g2_decap_8 FILLER_199_1142 ();
 sg13g2_decap_8 FILLER_199_1149 ();
 sg13g2_decap_8 FILLER_199_1156 ();
 sg13g2_decap_8 FILLER_199_1163 ();
 sg13g2_decap_8 FILLER_199_1170 ();
 sg13g2_decap_8 FILLER_199_1177 ();
 sg13g2_decap_8 FILLER_199_1184 ();
 sg13g2_decap_8 FILLER_199_1191 ();
 sg13g2_decap_8 FILLER_199_1198 ();
 sg13g2_decap_8 FILLER_199_1205 ();
 sg13g2_decap_8 FILLER_199_1212 ();
 sg13g2_decap_8 FILLER_199_1219 ();
 sg13g2_decap_8 FILLER_199_1226 ();
 sg13g2_decap_8 FILLER_199_1233 ();
 sg13g2_decap_8 FILLER_199_1240 ();
 sg13g2_decap_8 FILLER_199_1247 ();
 sg13g2_decap_8 FILLER_199_1254 ();
 sg13g2_decap_8 FILLER_199_1261 ();
 sg13g2_decap_8 FILLER_199_1268 ();
 sg13g2_decap_8 FILLER_199_1275 ();
 sg13g2_decap_8 FILLER_199_1282 ();
 sg13g2_decap_8 FILLER_199_1289 ();
 sg13g2_decap_8 FILLER_199_1296 ();
 sg13g2_decap_8 FILLER_199_1303 ();
 sg13g2_decap_8 FILLER_199_1310 ();
 sg13g2_decap_8 FILLER_199_1317 ();
 sg13g2_decap_8 FILLER_199_1324 ();
 sg13g2_decap_8 FILLER_199_1331 ();
 sg13g2_decap_8 FILLER_199_1338 ();
 sg13g2_decap_8 FILLER_199_1345 ();
 sg13g2_decap_8 FILLER_199_1352 ();
 sg13g2_decap_8 FILLER_199_1359 ();
 sg13g2_decap_8 FILLER_199_1366 ();
 sg13g2_decap_8 FILLER_199_1373 ();
 sg13g2_decap_8 FILLER_199_1380 ();
 sg13g2_decap_8 FILLER_199_1387 ();
 sg13g2_decap_8 FILLER_199_1394 ();
 sg13g2_decap_8 FILLER_199_1401 ();
 sg13g2_decap_8 FILLER_199_1408 ();
 sg13g2_decap_8 FILLER_199_1415 ();
 sg13g2_decap_8 FILLER_199_1422 ();
 sg13g2_decap_8 FILLER_199_1429 ();
 sg13g2_decap_8 FILLER_199_1436 ();
 sg13g2_decap_8 FILLER_199_1443 ();
 sg13g2_decap_8 FILLER_199_1450 ();
 sg13g2_decap_8 FILLER_199_1457 ();
 sg13g2_decap_8 FILLER_199_1464 ();
 sg13g2_decap_8 FILLER_199_1471 ();
 sg13g2_decap_8 FILLER_199_1478 ();
 sg13g2_decap_8 FILLER_199_1485 ();
 sg13g2_decap_8 FILLER_199_1492 ();
 sg13g2_decap_8 FILLER_199_1499 ();
 sg13g2_decap_8 FILLER_199_1506 ();
 sg13g2_decap_8 FILLER_199_1513 ();
 sg13g2_decap_8 FILLER_199_1520 ();
 sg13g2_decap_8 FILLER_199_1527 ();
 sg13g2_decap_8 FILLER_199_1534 ();
 sg13g2_decap_8 FILLER_199_1541 ();
 sg13g2_decap_8 FILLER_199_1548 ();
 sg13g2_decap_8 FILLER_199_1555 ();
 sg13g2_decap_8 FILLER_199_1562 ();
 sg13g2_decap_8 FILLER_199_1569 ();
 sg13g2_decap_8 FILLER_199_1576 ();
 sg13g2_decap_8 FILLER_199_1583 ();
 sg13g2_decap_8 FILLER_199_1590 ();
 sg13g2_decap_8 FILLER_199_1597 ();
 sg13g2_decap_8 FILLER_199_1604 ();
 sg13g2_decap_8 FILLER_199_1611 ();
 sg13g2_decap_8 FILLER_199_1618 ();
 sg13g2_decap_8 FILLER_200_0 ();
 sg13g2_decap_8 FILLER_200_7 ();
 sg13g2_decap_8 FILLER_200_14 ();
 sg13g2_decap_8 FILLER_200_21 ();
 sg13g2_decap_8 FILLER_200_28 ();
 sg13g2_decap_8 FILLER_200_35 ();
 sg13g2_decap_8 FILLER_200_42 ();
 sg13g2_decap_8 FILLER_200_49 ();
 sg13g2_decap_8 FILLER_200_56 ();
 sg13g2_decap_8 FILLER_200_63 ();
 sg13g2_decap_8 FILLER_200_70 ();
 sg13g2_decap_8 FILLER_200_77 ();
 sg13g2_decap_8 FILLER_200_84 ();
 sg13g2_decap_8 FILLER_200_91 ();
 sg13g2_decap_8 FILLER_200_98 ();
 sg13g2_decap_8 FILLER_200_105 ();
 sg13g2_decap_8 FILLER_200_112 ();
 sg13g2_decap_8 FILLER_200_119 ();
 sg13g2_decap_8 FILLER_200_126 ();
 sg13g2_decap_8 FILLER_200_133 ();
 sg13g2_decap_8 FILLER_200_140 ();
 sg13g2_decap_8 FILLER_200_147 ();
 sg13g2_decap_8 FILLER_200_154 ();
 sg13g2_decap_8 FILLER_200_161 ();
 sg13g2_decap_8 FILLER_200_168 ();
 sg13g2_decap_8 FILLER_200_175 ();
 sg13g2_decap_8 FILLER_200_182 ();
 sg13g2_decap_8 FILLER_200_189 ();
 sg13g2_decap_8 FILLER_200_196 ();
 sg13g2_decap_8 FILLER_200_203 ();
 sg13g2_decap_8 FILLER_200_210 ();
 sg13g2_decap_8 FILLER_200_217 ();
 sg13g2_decap_8 FILLER_200_224 ();
 sg13g2_decap_8 FILLER_200_231 ();
 sg13g2_decap_8 FILLER_200_238 ();
 sg13g2_decap_8 FILLER_200_245 ();
 sg13g2_decap_8 FILLER_200_252 ();
 sg13g2_decap_8 FILLER_200_259 ();
 sg13g2_decap_8 FILLER_200_266 ();
 sg13g2_decap_8 FILLER_200_273 ();
 sg13g2_decap_8 FILLER_200_280 ();
 sg13g2_decap_8 FILLER_200_287 ();
 sg13g2_decap_8 FILLER_200_294 ();
 sg13g2_decap_8 FILLER_200_301 ();
 sg13g2_decap_8 FILLER_200_308 ();
 sg13g2_decap_8 FILLER_200_315 ();
 sg13g2_decap_8 FILLER_200_322 ();
 sg13g2_decap_8 FILLER_200_329 ();
 sg13g2_decap_8 FILLER_200_336 ();
 sg13g2_decap_8 FILLER_200_343 ();
 sg13g2_decap_8 FILLER_200_350 ();
 sg13g2_decap_8 FILLER_200_357 ();
 sg13g2_decap_8 FILLER_200_364 ();
 sg13g2_decap_8 FILLER_200_371 ();
 sg13g2_decap_8 FILLER_200_378 ();
 sg13g2_fill_1 FILLER_200_385 ();
 sg13g2_decap_8 FILLER_200_390 ();
 sg13g2_decap_8 FILLER_200_397 ();
 sg13g2_decap_8 FILLER_200_404 ();
 sg13g2_decap_8 FILLER_200_411 ();
 sg13g2_decap_8 FILLER_200_418 ();
 sg13g2_decap_8 FILLER_200_425 ();
 sg13g2_decap_8 FILLER_200_432 ();
 sg13g2_decap_8 FILLER_200_439 ();
 sg13g2_decap_4 FILLER_200_446 ();
 sg13g2_fill_1 FILLER_200_450 ();
 sg13g2_decap_8 FILLER_200_477 ();
 sg13g2_decap_8 FILLER_200_484 ();
 sg13g2_decap_8 FILLER_200_491 ();
 sg13g2_fill_2 FILLER_200_498 ();
 sg13g2_decap_4 FILLER_200_504 ();
 sg13g2_fill_1 FILLER_200_508 ();
 sg13g2_fill_2 FILLER_200_539 ();
 sg13g2_decap_4 FILLER_200_567 ();
 sg13g2_fill_2 FILLER_200_571 ();
 sg13g2_decap_8 FILLER_200_585 ();
 sg13g2_fill_1 FILLER_200_601 ();
 sg13g2_decap_8 FILLER_200_614 ();
 sg13g2_decap_8 FILLER_200_621 ();
 sg13g2_fill_2 FILLER_200_628 ();
 sg13g2_fill_1 FILLER_200_630 ();
 sg13g2_fill_2 FILLER_200_639 ();
 sg13g2_fill_1 FILLER_200_641 ();
 sg13g2_decap_4 FILLER_200_646 ();
 sg13g2_fill_2 FILLER_200_650 ();
 sg13g2_decap_8 FILLER_200_656 ();
 sg13g2_decap_8 FILLER_200_663 ();
 sg13g2_decap_8 FILLER_200_670 ();
 sg13g2_decap_8 FILLER_200_677 ();
 sg13g2_decap_4 FILLER_200_684 ();
 sg13g2_fill_2 FILLER_200_696 ();
 sg13g2_decap_8 FILLER_200_723 ();
 sg13g2_decap_8 FILLER_200_730 ();
 sg13g2_decap_8 FILLER_200_737 ();
 sg13g2_decap_8 FILLER_200_744 ();
 sg13g2_decap_8 FILLER_200_751 ();
 sg13g2_decap_8 FILLER_200_758 ();
 sg13g2_decap_8 FILLER_200_765 ();
 sg13g2_decap_8 FILLER_200_772 ();
 sg13g2_decap_8 FILLER_200_779 ();
 sg13g2_decap_8 FILLER_200_786 ();
 sg13g2_decap_8 FILLER_200_793 ();
 sg13g2_decap_8 FILLER_200_800 ();
 sg13g2_decap_8 FILLER_200_807 ();
 sg13g2_decap_8 FILLER_200_814 ();
 sg13g2_decap_8 FILLER_200_821 ();
 sg13g2_decap_8 FILLER_200_828 ();
 sg13g2_decap_8 FILLER_200_835 ();
 sg13g2_decap_8 FILLER_200_842 ();
 sg13g2_decap_8 FILLER_200_849 ();
 sg13g2_decap_8 FILLER_200_856 ();
 sg13g2_decap_8 FILLER_200_863 ();
 sg13g2_decap_4 FILLER_200_870 ();
 sg13g2_decap_8 FILLER_200_900 ();
 sg13g2_decap_8 FILLER_200_907 ();
 sg13g2_decap_8 FILLER_200_914 ();
 sg13g2_decap_8 FILLER_200_921 ();
 sg13g2_decap_8 FILLER_200_928 ();
 sg13g2_decap_8 FILLER_200_935 ();
 sg13g2_decap_8 FILLER_200_942 ();
 sg13g2_decap_8 FILLER_200_949 ();
 sg13g2_decap_8 FILLER_200_956 ();
 sg13g2_decap_8 FILLER_200_963 ();
 sg13g2_decap_8 FILLER_200_970 ();
 sg13g2_decap_8 FILLER_200_977 ();
 sg13g2_decap_8 FILLER_200_984 ();
 sg13g2_decap_8 FILLER_200_991 ();
 sg13g2_decap_8 FILLER_200_998 ();
 sg13g2_decap_8 FILLER_200_1005 ();
 sg13g2_decap_8 FILLER_200_1012 ();
 sg13g2_decap_8 FILLER_200_1019 ();
 sg13g2_decap_8 FILLER_200_1026 ();
 sg13g2_decap_8 FILLER_200_1033 ();
 sg13g2_decap_8 FILLER_200_1040 ();
 sg13g2_decap_8 FILLER_200_1047 ();
 sg13g2_decap_8 FILLER_200_1054 ();
 sg13g2_decap_8 FILLER_200_1061 ();
 sg13g2_decap_8 FILLER_200_1068 ();
 sg13g2_decap_8 FILLER_200_1075 ();
 sg13g2_decap_8 FILLER_200_1082 ();
 sg13g2_decap_8 FILLER_200_1089 ();
 sg13g2_decap_8 FILLER_200_1096 ();
 sg13g2_decap_8 FILLER_200_1103 ();
 sg13g2_decap_8 FILLER_200_1110 ();
 sg13g2_decap_8 FILLER_200_1117 ();
 sg13g2_decap_8 FILLER_200_1124 ();
 sg13g2_decap_8 FILLER_200_1131 ();
 sg13g2_decap_8 FILLER_200_1138 ();
 sg13g2_decap_8 FILLER_200_1145 ();
 sg13g2_decap_8 FILLER_200_1152 ();
 sg13g2_decap_8 FILLER_200_1159 ();
 sg13g2_decap_8 FILLER_200_1166 ();
 sg13g2_decap_8 FILLER_200_1173 ();
 sg13g2_decap_8 FILLER_200_1180 ();
 sg13g2_decap_8 FILLER_200_1187 ();
 sg13g2_decap_8 FILLER_200_1194 ();
 sg13g2_decap_8 FILLER_200_1201 ();
 sg13g2_decap_8 FILLER_200_1208 ();
 sg13g2_decap_8 FILLER_200_1215 ();
 sg13g2_decap_8 FILLER_200_1222 ();
 sg13g2_decap_8 FILLER_200_1229 ();
 sg13g2_decap_8 FILLER_200_1236 ();
 sg13g2_decap_8 FILLER_200_1243 ();
 sg13g2_decap_8 FILLER_200_1250 ();
 sg13g2_decap_8 FILLER_200_1257 ();
 sg13g2_decap_8 FILLER_200_1264 ();
 sg13g2_decap_8 FILLER_200_1271 ();
 sg13g2_decap_8 FILLER_200_1278 ();
 sg13g2_decap_8 FILLER_200_1285 ();
 sg13g2_decap_8 FILLER_200_1292 ();
 sg13g2_decap_8 FILLER_200_1299 ();
 sg13g2_decap_8 FILLER_200_1306 ();
 sg13g2_decap_8 FILLER_200_1313 ();
 sg13g2_decap_8 FILLER_200_1320 ();
 sg13g2_decap_8 FILLER_200_1327 ();
 sg13g2_decap_8 FILLER_200_1334 ();
 sg13g2_decap_8 FILLER_200_1341 ();
 sg13g2_decap_8 FILLER_200_1348 ();
 sg13g2_decap_8 FILLER_200_1355 ();
 sg13g2_decap_8 FILLER_200_1362 ();
 sg13g2_decap_8 FILLER_200_1369 ();
 sg13g2_decap_8 FILLER_200_1376 ();
 sg13g2_decap_8 FILLER_200_1383 ();
 sg13g2_decap_8 FILLER_200_1390 ();
 sg13g2_decap_8 FILLER_200_1397 ();
 sg13g2_decap_8 FILLER_200_1404 ();
 sg13g2_decap_8 FILLER_200_1411 ();
 sg13g2_decap_8 FILLER_200_1418 ();
 sg13g2_decap_8 FILLER_200_1425 ();
 sg13g2_decap_8 FILLER_200_1432 ();
 sg13g2_decap_8 FILLER_200_1439 ();
 sg13g2_decap_8 FILLER_200_1446 ();
 sg13g2_decap_8 FILLER_200_1453 ();
 sg13g2_decap_8 FILLER_200_1460 ();
 sg13g2_decap_8 FILLER_200_1467 ();
 sg13g2_decap_8 FILLER_200_1474 ();
 sg13g2_decap_8 FILLER_200_1481 ();
 sg13g2_decap_8 FILLER_200_1488 ();
 sg13g2_decap_8 FILLER_200_1495 ();
 sg13g2_decap_8 FILLER_200_1502 ();
 sg13g2_decap_8 FILLER_200_1509 ();
 sg13g2_decap_8 FILLER_200_1516 ();
 sg13g2_decap_8 FILLER_200_1523 ();
 sg13g2_decap_8 FILLER_200_1530 ();
 sg13g2_decap_8 FILLER_200_1537 ();
 sg13g2_decap_8 FILLER_200_1544 ();
 sg13g2_decap_8 FILLER_200_1551 ();
 sg13g2_decap_8 FILLER_200_1558 ();
 sg13g2_decap_8 FILLER_200_1565 ();
 sg13g2_decap_8 FILLER_200_1572 ();
 sg13g2_decap_8 FILLER_200_1579 ();
 sg13g2_decap_8 FILLER_200_1586 ();
 sg13g2_decap_8 FILLER_200_1593 ();
 sg13g2_decap_8 FILLER_200_1600 ();
 sg13g2_decap_8 FILLER_200_1607 ();
 sg13g2_decap_8 FILLER_200_1614 ();
 sg13g2_decap_4 FILLER_200_1621 ();
 sg13g2_decap_8 FILLER_201_0 ();
 sg13g2_decap_8 FILLER_201_7 ();
 sg13g2_decap_8 FILLER_201_14 ();
 sg13g2_decap_8 FILLER_201_21 ();
 sg13g2_decap_8 FILLER_201_28 ();
 sg13g2_decap_8 FILLER_201_35 ();
 sg13g2_decap_8 FILLER_201_42 ();
 sg13g2_decap_8 FILLER_201_49 ();
 sg13g2_decap_8 FILLER_201_56 ();
 sg13g2_decap_8 FILLER_201_63 ();
 sg13g2_decap_8 FILLER_201_70 ();
 sg13g2_decap_8 FILLER_201_77 ();
 sg13g2_decap_8 FILLER_201_84 ();
 sg13g2_decap_8 FILLER_201_91 ();
 sg13g2_decap_8 FILLER_201_98 ();
 sg13g2_decap_8 FILLER_201_105 ();
 sg13g2_decap_8 FILLER_201_112 ();
 sg13g2_decap_8 FILLER_201_119 ();
 sg13g2_decap_8 FILLER_201_126 ();
 sg13g2_decap_8 FILLER_201_133 ();
 sg13g2_decap_8 FILLER_201_140 ();
 sg13g2_decap_8 FILLER_201_147 ();
 sg13g2_decap_8 FILLER_201_154 ();
 sg13g2_decap_8 FILLER_201_161 ();
 sg13g2_decap_8 FILLER_201_168 ();
 sg13g2_decap_8 FILLER_201_175 ();
 sg13g2_decap_8 FILLER_201_182 ();
 sg13g2_decap_8 FILLER_201_189 ();
 sg13g2_decap_8 FILLER_201_196 ();
 sg13g2_decap_8 FILLER_201_203 ();
 sg13g2_decap_8 FILLER_201_210 ();
 sg13g2_decap_8 FILLER_201_217 ();
 sg13g2_decap_8 FILLER_201_224 ();
 sg13g2_decap_8 FILLER_201_231 ();
 sg13g2_decap_8 FILLER_201_238 ();
 sg13g2_decap_8 FILLER_201_245 ();
 sg13g2_decap_8 FILLER_201_252 ();
 sg13g2_decap_8 FILLER_201_259 ();
 sg13g2_decap_8 FILLER_201_266 ();
 sg13g2_decap_8 FILLER_201_273 ();
 sg13g2_decap_8 FILLER_201_280 ();
 sg13g2_decap_8 FILLER_201_287 ();
 sg13g2_decap_8 FILLER_201_294 ();
 sg13g2_decap_8 FILLER_201_301 ();
 sg13g2_decap_8 FILLER_201_308 ();
 sg13g2_decap_8 FILLER_201_315 ();
 sg13g2_decap_8 FILLER_201_322 ();
 sg13g2_decap_8 FILLER_201_329 ();
 sg13g2_decap_8 FILLER_201_336 ();
 sg13g2_decap_8 FILLER_201_343 ();
 sg13g2_decap_8 FILLER_201_350 ();
 sg13g2_decap_8 FILLER_201_357 ();
 sg13g2_decap_8 FILLER_201_364 ();
 sg13g2_decap_8 FILLER_201_371 ();
 sg13g2_decap_8 FILLER_201_378 ();
 sg13g2_decap_8 FILLER_201_385 ();
 sg13g2_decap_8 FILLER_201_392 ();
 sg13g2_decap_8 FILLER_201_399 ();
 sg13g2_decap_8 FILLER_201_406 ();
 sg13g2_decap_8 FILLER_201_413 ();
 sg13g2_decap_8 FILLER_201_420 ();
 sg13g2_decap_8 FILLER_201_427 ();
 sg13g2_decap_8 FILLER_201_434 ();
 sg13g2_decap_8 FILLER_201_441 ();
 sg13g2_decap_8 FILLER_201_448 ();
 sg13g2_fill_2 FILLER_201_455 ();
 sg13g2_fill_1 FILLER_201_457 ();
 sg13g2_decap_8 FILLER_201_462 ();
 sg13g2_decap_4 FILLER_201_469 ();
 sg13g2_fill_2 FILLER_201_473 ();
 sg13g2_decap_8 FILLER_201_491 ();
 sg13g2_decap_8 FILLER_201_498 ();
 sg13g2_decap_8 FILLER_201_505 ();
 sg13g2_decap_8 FILLER_201_512 ();
 sg13g2_fill_2 FILLER_201_519 ();
 sg13g2_fill_1 FILLER_201_521 ();
 sg13g2_fill_1 FILLER_201_539 ();
 sg13g2_decap_4 FILLER_201_544 ();
 sg13g2_fill_1 FILLER_201_548 ();
 sg13g2_decap_8 FILLER_201_553 ();
 sg13g2_decap_8 FILLER_201_560 ();
 sg13g2_fill_1 FILLER_201_567 ();
 sg13g2_fill_1 FILLER_201_635 ();
 sg13g2_decap_8 FILLER_201_670 ();
 sg13g2_decap_8 FILLER_201_677 ();
 sg13g2_decap_4 FILLER_201_684 ();
 sg13g2_fill_1 FILLER_201_688 ();
 sg13g2_decap_8 FILLER_201_719 ();
 sg13g2_decap_8 FILLER_201_726 ();
 sg13g2_decap_8 FILLER_201_733 ();
 sg13g2_decap_8 FILLER_201_740 ();
 sg13g2_decap_8 FILLER_201_747 ();
 sg13g2_decap_8 FILLER_201_754 ();
 sg13g2_decap_8 FILLER_201_761 ();
 sg13g2_decap_8 FILLER_201_768 ();
 sg13g2_decap_8 FILLER_201_775 ();
 sg13g2_decap_8 FILLER_201_782 ();
 sg13g2_decap_8 FILLER_201_789 ();
 sg13g2_decap_8 FILLER_201_796 ();
 sg13g2_decap_8 FILLER_201_803 ();
 sg13g2_decap_8 FILLER_201_810 ();
 sg13g2_decap_8 FILLER_201_817 ();
 sg13g2_decap_8 FILLER_201_824 ();
 sg13g2_decap_8 FILLER_201_831 ();
 sg13g2_decap_8 FILLER_201_838 ();
 sg13g2_decap_8 FILLER_201_845 ();
 sg13g2_decap_8 FILLER_201_852 ();
 sg13g2_decap_8 FILLER_201_859 ();
 sg13g2_decap_8 FILLER_201_866 ();
 sg13g2_decap_8 FILLER_201_873 ();
 sg13g2_decap_8 FILLER_201_880 ();
 sg13g2_decap_8 FILLER_201_887 ();
 sg13g2_decap_8 FILLER_201_894 ();
 sg13g2_decap_8 FILLER_201_901 ();
 sg13g2_decap_8 FILLER_201_908 ();
 sg13g2_decap_8 FILLER_201_915 ();
 sg13g2_decap_8 FILLER_201_922 ();
 sg13g2_decap_8 FILLER_201_929 ();
 sg13g2_decap_8 FILLER_201_936 ();
 sg13g2_decap_8 FILLER_201_943 ();
 sg13g2_decap_8 FILLER_201_950 ();
 sg13g2_decap_8 FILLER_201_957 ();
 sg13g2_decap_8 FILLER_201_964 ();
 sg13g2_decap_8 FILLER_201_971 ();
 sg13g2_decap_8 FILLER_201_978 ();
 sg13g2_decap_8 FILLER_201_985 ();
 sg13g2_decap_8 FILLER_201_992 ();
 sg13g2_decap_8 FILLER_201_999 ();
 sg13g2_decap_8 FILLER_201_1006 ();
 sg13g2_decap_8 FILLER_201_1013 ();
 sg13g2_decap_8 FILLER_201_1020 ();
 sg13g2_decap_8 FILLER_201_1027 ();
 sg13g2_decap_8 FILLER_201_1034 ();
 sg13g2_decap_8 FILLER_201_1041 ();
 sg13g2_decap_8 FILLER_201_1048 ();
 sg13g2_decap_8 FILLER_201_1055 ();
 sg13g2_decap_8 FILLER_201_1062 ();
 sg13g2_decap_8 FILLER_201_1069 ();
 sg13g2_decap_8 FILLER_201_1076 ();
 sg13g2_decap_8 FILLER_201_1083 ();
 sg13g2_decap_8 FILLER_201_1090 ();
 sg13g2_decap_8 FILLER_201_1097 ();
 sg13g2_decap_8 FILLER_201_1104 ();
 sg13g2_decap_8 FILLER_201_1111 ();
 sg13g2_decap_8 FILLER_201_1118 ();
 sg13g2_decap_8 FILLER_201_1125 ();
 sg13g2_decap_8 FILLER_201_1132 ();
 sg13g2_decap_8 FILLER_201_1139 ();
 sg13g2_decap_8 FILLER_201_1146 ();
 sg13g2_decap_8 FILLER_201_1153 ();
 sg13g2_decap_8 FILLER_201_1160 ();
 sg13g2_decap_8 FILLER_201_1167 ();
 sg13g2_decap_8 FILLER_201_1174 ();
 sg13g2_decap_8 FILLER_201_1181 ();
 sg13g2_decap_8 FILLER_201_1188 ();
 sg13g2_decap_8 FILLER_201_1195 ();
 sg13g2_decap_8 FILLER_201_1202 ();
 sg13g2_decap_8 FILLER_201_1209 ();
 sg13g2_decap_8 FILLER_201_1216 ();
 sg13g2_decap_8 FILLER_201_1223 ();
 sg13g2_decap_8 FILLER_201_1230 ();
 sg13g2_decap_8 FILLER_201_1237 ();
 sg13g2_decap_8 FILLER_201_1244 ();
 sg13g2_decap_8 FILLER_201_1251 ();
 sg13g2_decap_8 FILLER_201_1258 ();
 sg13g2_decap_8 FILLER_201_1265 ();
 sg13g2_decap_8 FILLER_201_1272 ();
 sg13g2_decap_8 FILLER_201_1279 ();
 sg13g2_decap_8 FILLER_201_1286 ();
 sg13g2_decap_8 FILLER_201_1293 ();
 sg13g2_decap_8 FILLER_201_1300 ();
 sg13g2_decap_8 FILLER_201_1307 ();
 sg13g2_decap_8 FILLER_201_1314 ();
 sg13g2_decap_8 FILLER_201_1321 ();
 sg13g2_decap_8 FILLER_201_1328 ();
 sg13g2_decap_8 FILLER_201_1335 ();
 sg13g2_decap_8 FILLER_201_1342 ();
 sg13g2_decap_8 FILLER_201_1349 ();
 sg13g2_decap_8 FILLER_201_1356 ();
 sg13g2_decap_8 FILLER_201_1363 ();
 sg13g2_decap_8 FILLER_201_1370 ();
 sg13g2_decap_8 FILLER_201_1377 ();
 sg13g2_decap_8 FILLER_201_1384 ();
 sg13g2_decap_8 FILLER_201_1391 ();
 sg13g2_decap_8 FILLER_201_1398 ();
 sg13g2_decap_8 FILLER_201_1405 ();
 sg13g2_decap_8 FILLER_201_1412 ();
 sg13g2_decap_8 FILLER_201_1419 ();
 sg13g2_decap_8 FILLER_201_1426 ();
 sg13g2_decap_8 FILLER_201_1433 ();
 sg13g2_decap_8 FILLER_201_1440 ();
 sg13g2_decap_8 FILLER_201_1447 ();
 sg13g2_decap_8 FILLER_201_1454 ();
 sg13g2_decap_8 FILLER_201_1461 ();
 sg13g2_decap_8 FILLER_201_1468 ();
 sg13g2_decap_8 FILLER_201_1475 ();
 sg13g2_decap_8 FILLER_201_1482 ();
 sg13g2_decap_8 FILLER_201_1489 ();
 sg13g2_decap_8 FILLER_201_1496 ();
 sg13g2_decap_8 FILLER_201_1503 ();
 sg13g2_decap_8 FILLER_201_1510 ();
 sg13g2_decap_8 FILLER_201_1517 ();
 sg13g2_decap_8 FILLER_201_1524 ();
 sg13g2_decap_8 FILLER_201_1531 ();
 sg13g2_decap_8 FILLER_201_1538 ();
 sg13g2_decap_8 FILLER_201_1545 ();
 sg13g2_decap_8 FILLER_201_1552 ();
 sg13g2_decap_8 FILLER_201_1559 ();
 sg13g2_decap_8 FILLER_201_1566 ();
 sg13g2_decap_8 FILLER_201_1573 ();
 sg13g2_decap_8 FILLER_201_1580 ();
 sg13g2_decap_8 FILLER_201_1587 ();
 sg13g2_decap_8 FILLER_201_1594 ();
 sg13g2_decap_8 FILLER_201_1601 ();
 sg13g2_decap_8 FILLER_201_1608 ();
 sg13g2_decap_8 FILLER_201_1615 ();
 sg13g2_fill_2 FILLER_201_1622 ();
 sg13g2_fill_1 FILLER_201_1624 ();
 sg13g2_decap_8 FILLER_202_0 ();
 sg13g2_decap_8 FILLER_202_7 ();
 sg13g2_decap_8 FILLER_202_14 ();
 sg13g2_decap_8 FILLER_202_21 ();
 sg13g2_decap_8 FILLER_202_28 ();
 sg13g2_decap_8 FILLER_202_35 ();
 sg13g2_decap_8 FILLER_202_42 ();
 sg13g2_decap_8 FILLER_202_49 ();
 sg13g2_decap_8 FILLER_202_56 ();
 sg13g2_decap_8 FILLER_202_63 ();
 sg13g2_decap_8 FILLER_202_70 ();
 sg13g2_decap_8 FILLER_202_77 ();
 sg13g2_decap_8 FILLER_202_84 ();
 sg13g2_decap_8 FILLER_202_91 ();
 sg13g2_decap_8 FILLER_202_98 ();
 sg13g2_decap_8 FILLER_202_105 ();
 sg13g2_decap_8 FILLER_202_112 ();
 sg13g2_decap_8 FILLER_202_119 ();
 sg13g2_decap_8 FILLER_202_126 ();
 sg13g2_decap_8 FILLER_202_133 ();
 sg13g2_decap_8 FILLER_202_140 ();
 sg13g2_decap_8 FILLER_202_147 ();
 sg13g2_decap_8 FILLER_202_154 ();
 sg13g2_decap_8 FILLER_202_161 ();
 sg13g2_decap_8 FILLER_202_168 ();
 sg13g2_decap_8 FILLER_202_175 ();
 sg13g2_decap_8 FILLER_202_182 ();
 sg13g2_decap_8 FILLER_202_189 ();
 sg13g2_decap_8 FILLER_202_196 ();
 sg13g2_decap_8 FILLER_202_203 ();
 sg13g2_decap_8 FILLER_202_210 ();
 sg13g2_decap_8 FILLER_202_217 ();
 sg13g2_decap_8 FILLER_202_224 ();
 sg13g2_decap_8 FILLER_202_231 ();
 sg13g2_decap_8 FILLER_202_238 ();
 sg13g2_decap_8 FILLER_202_245 ();
 sg13g2_decap_8 FILLER_202_252 ();
 sg13g2_decap_8 FILLER_202_259 ();
 sg13g2_decap_8 FILLER_202_266 ();
 sg13g2_decap_8 FILLER_202_273 ();
 sg13g2_decap_8 FILLER_202_280 ();
 sg13g2_decap_8 FILLER_202_287 ();
 sg13g2_decap_8 FILLER_202_294 ();
 sg13g2_decap_8 FILLER_202_301 ();
 sg13g2_decap_8 FILLER_202_308 ();
 sg13g2_decap_8 FILLER_202_315 ();
 sg13g2_decap_8 FILLER_202_322 ();
 sg13g2_decap_8 FILLER_202_329 ();
 sg13g2_decap_8 FILLER_202_336 ();
 sg13g2_decap_8 FILLER_202_343 ();
 sg13g2_decap_8 FILLER_202_350 ();
 sg13g2_decap_8 FILLER_202_357 ();
 sg13g2_decap_8 FILLER_202_364 ();
 sg13g2_decap_8 FILLER_202_371 ();
 sg13g2_decap_8 FILLER_202_378 ();
 sg13g2_decap_8 FILLER_202_385 ();
 sg13g2_decap_8 FILLER_202_392 ();
 sg13g2_decap_8 FILLER_202_399 ();
 sg13g2_decap_8 FILLER_202_406 ();
 sg13g2_decap_8 FILLER_202_413 ();
 sg13g2_decap_8 FILLER_202_420 ();
 sg13g2_decap_8 FILLER_202_427 ();
 sg13g2_decap_8 FILLER_202_434 ();
 sg13g2_decap_8 FILLER_202_441 ();
 sg13g2_fill_2 FILLER_202_448 ();
 sg13g2_fill_1 FILLER_202_450 ();
 sg13g2_decap_8 FILLER_202_487 ();
 sg13g2_decap_4 FILLER_202_494 ();
 sg13g2_fill_2 FILLER_202_498 ();
 sg13g2_decap_8 FILLER_202_512 ();
 sg13g2_decap_8 FILLER_202_544 ();
 sg13g2_decap_8 FILLER_202_551 ();
 sg13g2_decap_8 FILLER_202_558 ();
 sg13g2_decap_4 FILLER_202_565 ();
 sg13g2_decap_8 FILLER_202_599 ();
 sg13g2_decap_4 FILLER_202_606 ();
 sg13g2_fill_1 FILLER_202_610 ();
 sg13g2_fill_2 FILLER_202_640 ();
 sg13g2_decap_8 FILLER_202_671 ();
 sg13g2_decap_8 FILLER_202_678 ();
 sg13g2_decap_8 FILLER_202_685 ();
 sg13g2_decap_8 FILLER_202_692 ();
 sg13g2_decap_8 FILLER_202_699 ();
 sg13g2_decap_8 FILLER_202_706 ();
 sg13g2_decap_8 FILLER_202_713 ();
 sg13g2_decap_8 FILLER_202_720 ();
 sg13g2_decap_8 FILLER_202_727 ();
 sg13g2_decap_8 FILLER_202_734 ();
 sg13g2_decap_8 FILLER_202_741 ();
 sg13g2_decap_8 FILLER_202_748 ();
 sg13g2_decap_8 FILLER_202_755 ();
 sg13g2_decap_8 FILLER_202_762 ();
 sg13g2_decap_8 FILLER_202_769 ();
 sg13g2_decap_8 FILLER_202_776 ();
 sg13g2_decap_8 FILLER_202_783 ();
 sg13g2_decap_8 FILLER_202_790 ();
 sg13g2_decap_8 FILLER_202_797 ();
 sg13g2_decap_8 FILLER_202_804 ();
 sg13g2_decap_8 FILLER_202_811 ();
 sg13g2_decap_8 FILLER_202_818 ();
 sg13g2_decap_8 FILLER_202_825 ();
 sg13g2_decap_8 FILLER_202_832 ();
 sg13g2_decap_8 FILLER_202_839 ();
 sg13g2_decap_8 FILLER_202_846 ();
 sg13g2_decap_8 FILLER_202_853 ();
 sg13g2_decap_8 FILLER_202_860 ();
 sg13g2_decap_8 FILLER_202_867 ();
 sg13g2_decap_8 FILLER_202_874 ();
 sg13g2_decap_8 FILLER_202_881 ();
 sg13g2_decap_8 FILLER_202_888 ();
 sg13g2_decap_8 FILLER_202_895 ();
 sg13g2_decap_8 FILLER_202_902 ();
 sg13g2_decap_8 FILLER_202_909 ();
 sg13g2_decap_8 FILLER_202_916 ();
 sg13g2_decap_8 FILLER_202_923 ();
 sg13g2_decap_8 FILLER_202_930 ();
 sg13g2_decap_8 FILLER_202_937 ();
 sg13g2_decap_8 FILLER_202_944 ();
 sg13g2_decap_8 FILLER_202_951 ();
 sg13g2_decap_8 FILLER_202_958 ();
 sg13g2_decap_8 FILLER_202_965 ();
 sg13g2_decap_8 FILLER_202_972 ();
 sg13g2_decap_8 FILLER_202_979 ();
 sg13g2_decap_8 FILLER_202_986 ();
 sg13g2_decap_8 FILLER_202_993 ();
 sg13g2_decap_8 FILLER_202_1000 ();
 sg13g2_decap_8 FILLER_202_1007 ();
 sg13g2_decap_8 FILLER_202_1014 ();
 sg13g2_decap_8 FILLER_202_1021 ();
 sg13g2_decap_8 FILLER_202_1028 ();
 sg13g2_decap_8 FILLER_202_1035 ();
 sg13g2_decap_8 FILLER_202_1042 ();
 sg13g2_decap_8 FILLER_202_1049 ();
 sg13g2_decap_8 FILLER_202_1056 ();
 sg13g2_decap_8 FILLER_202_1063 ();
 sg13g2_decap_8 FILLER_202_1070 ();
 sg13g2_decap_8 FILLER_202_1077 ();
 sg13g2_decap_8 FILLER_202_1084 ();
 sg13g2_decap_8 FILLER_202_1091 ();
 sg13g2_decap_8 FILLER_202_1098 ();
 sg13g2_decap_8 FILLER_202_1105 ();
 sg13g2_decap_8 FILLER_202_1112 ();
 sg13g2_decap_8 FILLER_202_1119 ();
 sg13g2_decap_8 FILLER_202_1126 ();
 sg13g2_decap_8 FILLER_202_1133 ();
 sg13g2_decap_8 FILLER_202_1140 ();
 sg13g2_decap_8 FILLER_202_1147 ();
 sg13g2_decap_8 FILLER_202_1154 ();
 sg13g2_decap_8 FILLER_202_1161 ();
 sg13g2_decap_8 FILLER_202_1168 ();
 sg13g2_decap_8 FILLER_202_1175 ();
 sg13g2_decap_8 FILLER_202_1182 ();
 sg13g2_decap_8 FILLER_202_1189 ();
 sg13g2_decap_8 FILLER_202_1196 ();
 sg13g2_decap_8 FILLER_202_1203 ();
 sg13g2_decap_8 FILLER_202_1210 ();
 sg13g2_decap_8 FILLER_202_1217 ();
 sg13g2_decap_8 FILLER_202_1224 ();
 sg13g2_decap_8 FILLER_202_1231 ();
 sg13g2_decap_8 FILLER_202_1238 ();
 sg13g2_decap_8 FILLER_202_1245 ();
 sg13g2_decap_8 FILLER_202_1252 ();
 sg13g2_decap_8 FILLER_202_1259 ();
 sg13g2_decap_8 FILLER_202_1266 ();
 sg13g2_decap_8 FILLER_202_1273 ();
 sg13g2_decap_8 FILLER_202_1280 ();
 sg13g2_decap_8 FILLER_202_1287 ();
 sg13g2_decap_8 FILLER_202_1294 ();
 sg13g2_decap_8 FILLER_202_1301 ();
 sg13g2_decap_8 FILLER_202_1308 ();
 sg13g2_decap_8 FILLER_202_1315 ();
 sg13g2_decap_8 FILLER_202_1322 ();
 sg13g2_decap_8 FILLER_202_1329 ();
 sg13g2_decap_8 FILLER_202_1336 ();
 sg13g2_decap_8 FILLER_202_1343 ();
 sg13g2_decap_8 FILLER_202_1350 ();
 sg13g2_decap_8 FILLER_202_1357 ();
 sg13g2_decap_8 FILLER_202_1364 ();
 sg13g2_decap_8 FILLER_202_1371 ();
 sg13g2_decap_8 FILLER_202_1378 ();
 sg13g2_decap_8 FILLER_202_1385 ();
 sg13g2_decap_8 FILLER_202_1392 ();
 sg13g2_decap_8 FILLER_202_1399 ();
 sg13g2_decap_8 FILLER_202_1406 ();
 sg13g2_decap_8 FILLER_202_1413 ();
 sg13g2_decap_8 FILLER_202_1420 ();
 sg13g2_decap_8 FILLER_202_1427 ();
 sg13g2_decap_8 FILLER_202_1434 ();
 sg13g2_decap_8 FILLER_202_1441 ();
 sg13g2_decap_8 FILLER_202_1448 ();
 sg13g2_decap_8 FILLER_202_1455 ();
 sg13g2_decap_8 FILLER_202_1462 ();
 sg13g2_decap_8 FILLER_202_1469 ();
 sg13g2_decap_8 FILLER_202_1476 ();
 sg13g2_decap_8 FILLER_202_1483 ();
 sg13g2_decap_8 FILLER_202_1490 ();
 sg13g2_decap_8 FILLER_202_1497 ();
 sg13g2_decap_8 FILLER_202_1504 ();
 sg13g2_decap_8 FILLER_202_1511 ();
 sg13g2_decap_8 FILLER_202_1518 ();
 sg13g2_decap_8 FILLER_202_1525 ();
 sg13g2_decap_8 FILLER_202_1532 ();
 sg13g2_decap_8 FILLER_202_1539 ();
 sg13g2_decap_8 FILLER_202_1546 ();
 sg13g2_decap_8 FILLER_202_1553 ();
 sg13g2_decap_8 FILLER_202_1560 ();
 sg13g2_decap_8 FILLER_202_1567 ();
 sg13g2_decap_8 FILLER_202_1574 ();
 sg13g2_decap_8 FILLER_202_1581 ();
 sg13g2_decap_8 FILLER_202_1588 ();
 sg13g2_decap_8 FILLER_202_1595 ();
 sg13g2_decap_8 FILLER_202_1602 ();
 sg13g2_decap_8 FILLER_202_1609 ();
 sg13g2_decap_8 FILLER_202_1616 ();
 sg13g2_fill_2 FILLER_202_1623 ();
 sg13g2_decap_8 FILLER_203_0 ();
 sg13g2_decap_8 FILLER_203_7 ();
 sg13g2_decap_8 FILLER_203_14 ();
 sg13g2_decap_8 FILLER_203_21 ();
 sg13g2_decap_8 FILLER_203_28 ();
 sg13g2_decap_8 FILLER_203_35 ();
 sg13g2_decap_8 FILLER_203_42 ();
 sg13g2_decap_8 FILLER_203_49 ();
 sg13g2_decap_8 FILLER_203_56 ();
 sg13g2_decap_8 FILLER_203_63 ();
 sg13g2_decap_8 FILLER_203_70 ();
 sg13g2_decap_8 FILLER_203_77 ();
 sg13g2_decap_8 FILLER_203_84 ();
 sg13g2_decap_8 FILLER_203_91 ();
 sg13g2_decap_8 FILLER_203_98 ();
 sg13g2_decap_8 FILLER_203_105 ();
 sg13g2_decap_8 FILLER_203_112 ();
 sg13g2_decap_8 FILLER_203_119 ();
 sg13g2_decap_8 FILLER_203_126 ();
 sg13g2_decap_8 FILLER_203_133 ();
 sg13g2_decap_8 FILLER_203_140 ();
 sg13g2_decap_8 FILLER_203_147 ();
 sg13g2_decap_8 FILLER_203_154 ();
 sg13g2_decap_8 FILLER_203_161 ();
 sg13g2_decap_8 FILLER_203_168 ();
 sg13g2_decap_8 FILLER_203_175 ();
 sg13g2_decap_8 FILLER_203_182 ();
 sg13g2_decap_8 FILLER_203_189 ();
 sg13g2_decap_8 FILLER_203_196 ();
 sg13g2_decap_8 FILLER_203_203 ();
 sg13g2_decap_8 FILLER_203_210 ();
 sg13g2_decap_8 FILLER_203_217 ();
 sg13g2_decap_8 FILLER_203_224 ();
 sg13g2_decap_8 FILLER_203_231 ();
 sg13g2_decap_8 FILLER_203_238 ();
 sg13g2_decap_8 FILLER_203_245 ();
 sg13g2_decap_8 FILLER_203_252 ();
 sg13g2_decap_8 FILLER_203_259 ();
 sg13g2_decap_8 FILLER_203_266 ();
 sg13g2_decap_8 FILLER_203_273 ();
 sg13g2_decap_8 FILLER_203_280 ();
 sg13g2_decap_8 FILLER_203_287 ();
 sg13g2_decap_8 FILLER_203_294 ();
 sg13g2_decap_8 FILLER_203_301 ();
 sg13g2_decap_8 FILLER_203_308 ();
 sg13g2_decap_8 FILLER_203_315 ();
 sg13g2_decap_8 FILLER_203_322 ();
 sg13g2_decap_8 FILLER_203_329 ();
 sg13g2_decap_8 FILLER_203_336 ();
 sg13g2_decap_8 FILLER_203_343 ();
 sg13g2_decap_8 FILLER_203_350 ();
 sg13g2_decap_8 FILLER_203_357 ();
 sg13g2_decap_8 FILLER_203_364 ();
 sg13g2_decap_8 FILLER_203_371 ();
 sg13g2_decap_8 FILLER_203_378 ();
 sg13g2_decap_8 FILLER_203_385 ();
 sg13g2_decap_8 FILLER_203_392 ();
 sg13g2_decap_8 FILLER_203_399 ();
 sg13g2_decap_8 FILLER_203_406 ();
 sg13g2_decap_8 FILLER_203_413 ();
 sg13g2_decap_8 FILLER_203_420 ();
 sg13g2_decap_8 FILLER_203_427 ();
 sg13g2_decap_8 FILLER_203_434 ();
 sg13g2_decap_8 FILLER_203_441 ();
 sg13g2_fill_2 FILLER_203_526 ();
 sg13g2_decap_8 FILLER_203_554 ();
 sg13g2_decap_8 FILLER_203_561 ();
 sg13g2_decap_8 FILLER_203_568 ();
 sg13g2_decap_8 FILLER_203_575 ();
 sg13g2_decap_8 FILLER_203_582 ();
 sg13g2_decap_8 FILLER_203_589 ();
 sg13g2_decap_8 FILLER_203_596 ();
 sg13g2_decap_8 FILLER_203_603 ();
 sg13g2_fill_2 FILLER_203_610 ();
 sg13g2_decap_8 FILLER_203_664 ();
 sg13g2_decap_8 FILLER_203_671 ();
 sg13g2_decap_8 FILLER_203_678 ();
 sg13g2_decap_8 FILLER_203_685 ();
 sg13g2_decap_8 FILLER_203_692 ();
 sg13g2_decap_8 FILLER_203_699 ();
 sg13g2_decap_8 FILLER_203_706 ();
 sg13g2_decap_8 FILLER_203_713 ();
 sg13g2_decap_8 FILLER_203_720 ();
 sg13g2_decap_8 FILLER_203_727 ();
 sg13g2_decap_8 FILLER_203_734 ();
 sg13g2_decap_8 FILLER_203_741 ();
 sg13g2_decap_8 FILLER_203_748 ();
 sg13g2_decap_8 FILLER_203_755 ();
 sg13g2_decap_8 FILLER_203_762 ();
 sg13g2_decap_8 FILLER_203_769 ();
 sg13g2_decap_8 FILLER_203_776 ();
 sg13g2_decap_8 FILLER_203_783 ();
 sg13g2_decap_8 FILLER_203_790 ();
 sg13g2_decap_8 FILLER_203_797 ();
 sg13g2_decap_8 FILLER_203_804 ();
 sg13g2_decap_8 FILLER_203_811 ();
 sg13g2_decap_8 FILLER_203_818 ();
 sg13g2_decap_8 FILLER_203_825 ();
 sg13g2_decap_8 FILLER_203_832 ();
 sg13g2_decap_8 FILLER_203_839 ();
 sg13g2_decap_8 FILLER_203_846 ();
 sg13g2_decap_8 FILLER_203_853 ();
 sg13g2_decap_8 FILLER_203_860 ();
 sg13g2_decap_8 FILLER_203_867 ();
 sg13g2_decap_8 FILLER_203_874 ();
 sg13g2_decap_8 FILLER_203_881 ();
 sg13g2_decap_8 FILLER_203_888 ();
 sg13g2_decap_8 FILLER_203_895 ();
 sg13g2_decap_8 FILLER_203_902 ();
 sg13g2_decap_8 FILLER_203_909 ();
 sg13g2_decap_8 FILLER_203_916 ();
 sg13g2_decap_8 FILLER_203_923 ();
 sg13g2_decap_8 FILLER_203_930 ();
 sg13g2_decap_8 FILLER_203_937 ();
 sg13g2_decap_8 FILLER_203_944 ();
 sg13g2_decap_8 FILLER_203_951 ();
 sg13g2_decap_8 FILLER_203_958 ();
 sg13g2_decap_8 FILLER_203_965 ();
 sg13g2_decap_8 FILLER_203_972 ();
 sg13g2_decap_8 FILLER_203_979 ();
 sg13g2_decap_8 FILLER_203_986 ();
 sg13g2_decap_8 FILLER_203_993 ();
 sg13g2_decap_8 FILLER_203_1000 ();
 sg13g2_decap_8 FILLER_203_1007 ();
 sg13g2_decap_8 FILLER_203_1014 ();
 sg13g2_decap_8 FILLER_203_1021 ();
 sg13g2_decap_8 FILLER_203_1028 ();
 sg13g2_decap_8 FILLER_203_1035 ();
 sg13g2_decap_8 FILLER_203_1042 ();
 sg13g2_decap_8 FILLER_203_1049 ();
 sg13g2_decap_8 FILLER_203_1056 ();
 sg13g2_decap_8 FILLER_203_1063 ();
 sg13g2_decap_8 FILLER_203_1070 ();
 sg13g2_decap_8 FILLER_203_1077 ();
 sg13g2_decap_8 FILLER_203_1084 ();
 sg13g2_decap_8 FILLER_203_1091 ();
 sg13g2_decap_8 FILLER_203_1098 ();
 sg13g2_decap_8 FILLER_203_1105 ();
 sg13g2_decap_8 FILLER_203_1112 ();
 sg13g2_decap_8 FILLER_203_1119 ();
 sg13g2_decap_8 FILLER_203_1126 ();
 sg13g2_decap_8 FILLER_203_1133 ();
 sg13g2_decap_8 FILLER_203_1140 ();
 sg13g2_decap_8 FILLER_203_1147 ();
 sg13g2_decap_8 FILLER_203_1154 ();
 sg13g2_decap_8 FILLER_203_1161 ();
 sg13g2_decap_8 FILLER_203_1168 ();
 sg13g2_decap_8 FILLER_203_1175 ();
 sg13g2_decap_8 FILLER_203_1182 ();
 sg13g2_decap_8 FILLER_203_1189 ();
 sg13g2_decap_8 FILLER_203_1196 ();
 sg13g2_decap_8 FILLER_203_1203 ();
 sg13g2_decap_8 FILLER_203_1210 ();
 sg13g2_decap_8 FILLER_203_1217 ();
 sg13g2_decap_8 FILLER_203_1224 ();
 sg13g2_decap_8 FILLER_203_1231 ();
 sg13g2_decap_8 FILLER_203_1238 ();
 sg13g2_decap_8 FILLER_203_1245 ();
 sg13g2_decap_8 FILLER_203_1252 ();
 sg13g2_decap_8 FILLER_203_1259 ();
 sg13g2_decap_8 FILLER_203_1266 ();
 sg13g2_decap_8 FILLER_203_1273 ();
 sg13g2_decap_8 FILLER_203_1280 ();
 sg13g2_decap_8 FILLER_203_1287 ();
 sg13g2_decap_8 FILLER_203_1294 ();
 sg13g2_decap_8 FILLER_203_1301 ();
 sg13g2_decap_8 FILLER_203_1308 ();
 sg13g2_decap_8 FILLER_203_1315 ();
 sg13g2_decap_8 FILLER_203_1322 ();
 sg13g2_decap_8 FILLER_203_1329 ();
 sg13g2_decap_8 FILLER_203_1336 ();
 sg13g2_decap_8 FILLER_203_1343 ();
 sg13g2_decap_8 FILLER_203_1350 ();
 sg13g2_decap_8 FILLER_203_1357 ();
 sg13g2_decap_8 FILLER_203_1364 ();
 sg13g2_decap_8 FILLER_203_1371 ();
 sg13g2_decap_8 FILLER_203_1378 ();
 sg13g2_decap_8 FILLER_203_1385 ();
 sg13g2_decap_8 FILLER_203_1392 ();
 sg13g2_decap_8 FILLER_203_1399 ();
 sg13g2_decap_8 FILLER_203_1406 ();
 sg13g2_decap_8 FILLER_203_1413 ();
 sg13g2_decap_8 FILLER_203_1420 ();
 sg13g2_decap_8 FILLER_203_1427 ();
 sg13g2_decap_8 FILLER_203_1434 ();
 sg13g2_decap_8 FILLER_203_1441 ();
 sg13g2_decap_8 FILLER_203_1448 ();
 sg13g2_decap_8 FILLER_203_1455 ();
 sg13g2_decap_8 FILLER_203_1462 ();
 sg13g2_decap_8 FILLER_203_1469 ();
 sg13g2_decap_8 FILLER_203_1476 ();
 sg13g2_decap_8 FILLER_203_1483 ();
 sg13g2_decap_8 FILLER_203_1490 ();
 sg13g2_decap_8 FILLER_203_1497 ();
 sg13g2_decap_8 FILLER_203_1504 ();
 sg13g2_decap_8 FILLER_203_1511 ();
 sg13g2_decap_8 FILLER_203_1518 ();
 sg13g2_decap_8 FILLER_203_1525 ();
 sg13g2_decap_8 FILLER_203_1532 ();
 sg13g2_decap_8 FILLER_203_1539 ();
 sg13g2_decap_8 FILLER_203_1546 ();
 sg13g2_decap_8 FILLER_203_1553 ();
 sg13g2_decap_8 FILLER_203_1560 ();
 sg13g2_decap_8 FILLER_203_1567 ();
 sg13g2_decap_8 FILLER_203_1574 ();
 sg13g2_decap_8 FILLER_203_1581 ();
 sg13g2_decap_8 FILLER_203_1588 ();
 sg13g2_decap_8 FILLER_203_1595 ();
 sg13g2_decap_8 FILLER_203_1602 ();
 sg13g2_decap_8 FILLER_203_1609 ();
 sg13g2_decap_8 FILLER_203_1616 ();
 sg13g2_fill_2 FILLER_203_1623 ();
 sg13g2_decap_8 FILLER_204_0 ();
 sg13g2_decap_8 FILLER_204_7 ();
 sg13g2_decap_8 FILLER_204_14 ();
 sg13g2_decap_8 FILLER_204_21 ();
 sg13g2_decap_8 FILLER_204_28 ();
 sg13g2_decap_8 FILLER_204_35 ();
 sg13g2_decap_8 FILLER_204_42 ();
 sg13g2_decap_8 FILLER_204_49 ();
 sg13g2_decap_8 FILLER_204_56 ();
 sg13g2_decap_8 FILLER_204_63 ();
 sg13g2_decap_8 FILLER_204_70 ();
 sg13g2_decap_8 FILLER_204_77 ();
 sg13g2_decap_8 FILLER_204_84 ();
 sg13g2_decap_8 FILLER_204_91 ();
 sg13g2_decap_8 FILLER_204_98 ();
 sg13g2_decap_8 FILLER_204_105 ();
 sg13g2_decap_8 FILLER_204_112 ();
 sg13g2_decap_8 FILLER_204_119 ();
 sg13g2_decap_8 FILLER_204_126 ();
 sg13g2_decap_8 FILLER_204_133 ();
 sg13g2_decap_8 FILLER_204_140 ();
 sg13g2_decap_8 FILLER_204_147 ();
 sg13g2_decap_8 FILLER_204_154 ();
 sg13g2_decap_8 FILLER_204_161 ();
 sg13g2_decap_8 FILLER_204_168 ();
 sg13g2_decap_8 FILLER_204_175 ();
 sg13g2_decap_8 FILLER_204_182 ();
 sg13g2_decap_8 FILLER_204_189 ();
 sg13g2_decap_8 FILLER_204_196 ();
 sg13g2_decap_8 FILLER_204_203 ();
 sg13g2_decap_8 FILLER_204_210 ();
 sg13g2_decap_8 FILLER_204_217 ();
 sg13g2_decap_8 FILLER_204_224 ();
 sg13g2_decap_8 FILLER_204_231 ();
 sg13g2_decap_8 FILLER_204_238 ();
 sg13g2_decap_8 FILLER_204_245 ();
 sg13g2_decap_8 FILLER_204_252 ();
 sg13g2_decap_8 FILLER_204_259 ();
 sg13g2_decap_8 FILLER_204_266 ();
 sg13g2_decap_8 FILLER_204_273 ();
 sg13g2_decap_8 FILLER_204_280 ();
 sg13g2_decap_8 FILLER_204_287 ();
 sg13g2_decap_8 FILLER_204_294 ();
 sg13g2_decap_8 FILLER_204_301 ();
 sg13g2_decap_8 FILLER_204_308 ();
 sg13g2_decap_8 FILLER_204_315 ();
 sg13g2_decap_8 FILLER_204_322 ();
 sg13g2_decap_8 FILLER_204_329 ();
 sg13g2_decap_8 FILLER_204_336 ();
 sg13g2_decap_8 FILLER_204_343 ();
 sg13g2_decap_8 FILLER_204_350 ();
 sg13g2_decap_8 FILLER_204_357 ();
 sg13g2_decap_8 FILLER_204_364 ();
 sg13g2_decap_8 FILLER_204_371 ();
 sg13g2_decap_8 FILLER_204_378 ();
 sg13g2_decap_8 FILLER_204_385 ();
 sg13g2_decap_8 FILLER_204_392 ();
 sg13g2_decap_8 FILLER_204_399 ();
 sg13g2_decap_8 FILLER_204_406 ();
 sg13g2_decap_8 FILLER_204_413 ();
 sg13g2_decap_8 FILLER_204_420 ();
 sg13g2_decap_8 FILLER_204_427 ();
 sg13g2_decap_8 FILLER_204_434 ();
 sg13g2_decap_8 FILLER_204_441 ();
 sg13g2_decap_4 FILLER_204_448 ();
 sg13g2_fill_2 FILLER_204_452 ();
 sg13g2_decap_8 FILLER_204_458 ();
 sg13g2_decap_8 FILLER_204_465 ();
 sg13g2_decap_4 FILLER_204_472 ();
 sg13g2_fill_1 FILLER_204_476 ();
 sg13g2_decap_8 FILLER_204_485 ();
 sg13g2_decap_8 FILLER_204_492 ();
 sg13g2_fill_2 FILLER_204_499 ();
 sg13g2_decap_8 FILLER_204_505 ();
 sg13g2_decap_8 FILLER_204_512 ();
 sg13g2_decap_8 FILLER_204_519 ();
 sg13g2_fill_2 FILLER_204_526 ();
 sg13g2_fill_1 FILLER_204_528 ();
 sg13g2_fill_2 FILLER_204_533 ();
 sg13g2_decap_8 FILLER_204_539 ();
 sg13g2_decap_8 FILLER_204_546 ();
 sg13g2_decap_8 FILLER_204_553 ();
 sg13g2_decap_8 FILLER_204_560 ();
 sg13g2_decap_8 FILLER_204_567 ();
 sg13g2_decap_8 FILLER_204_574 ();
 sg13g2_decap_8 FILLER_204_581 ();
 sg13g2_decap_8 FILLER_204_588 ();
 sg13g2_decap_8 FILLER_204_595 ();
 sg13g2_decap_8 FILLER_204_602 ();
 sg13g2_decap_8 FILLER_204_609 ();
 sg13g2_decap_4 FILLER_204_616 ();
 sg13g2_fill_1 FILLER_204_620 ();
 sg13g2_decap_4 FILLER_204_625 ();
 sg13g2_decap_8 FILLER_204_633 ();
 sg13g2_decap_8 FILLER_204_640 ();
 sg13g2_decap_8 FILLER_204_647 ();
 sg13g2_decap_8 FILLER_204_654 ();
 sg13g2_decap_8 FILLER_204_661 ();
 sg13g2_decap_8 FILLER_204_668 ();
 sg13g2_decap_8 FILLER_204_675 ();
 sg13g2_decap_8 FILLER_204_682 ();
 sg13g2_decap_8 FILLER_204_689 ();
 sg13g2_decap_8 FILLER_204_696 ();
 sg13g2_decap_8 FILLER_204_703 ();
 sg13g2_decap_8 FILLER_204_710 ();
 sg13g2_decap_8 FILLER_204_717 ();
 sg13g2_decap_8 FILLER_204_724 ();
 sg13g2_decap_8 FILLER_204_731 ();
 sg13g2_decap_8 FILLER_204_738 ();
 sg13g2_decap_8 FILLER_204_745 ();
 sg13g2_decap_8 FILLER_204_752 ();
 sg13g2_decap_8 FILLER_204_759 ();
 sg13g2_decap_8 FILLER_204_766 ();
 sg13g2_decap_8 FILLER_204_773 ();
 sg13g2_decap_8 FILLER_204_780 ();
 sg13g2_decap_8 FILLER_204_787 ();
 sg13g2_decap_8 FILLER_204_794 ();
 sg13g2_decap_8 FILLER_204_801 ();
 sg13g2_decap_8 FILLER_204_808 ();
 sg13g2_decap_8 FILLER_204_815 ();
 sg13g2_decap_8 FILLER_204_822 ();
 sg13g2_decap_8 FILLER_204_829 ();
 sg13g2_decap_8 FILLER_204_836 ();
 sg13g2_decap_8 FILLER_204_843 ();
 sg13g2_decap_8 FILLER_204_850 ();
 sg13g2_decap_8 FILLER_204_857 ();
 sg13g2_decap_8 FILLER_204_864 ();
 sg13g2_decap_8 FILLER_204_871 ();
 sg13g2_decap_8 FILLER_204_878 ();
 sg13g2_decap_8 FILLER_204_885 ();
 sg13g2_decap_8 FILLER_204_892 ();
 sg13g2_decap_8 FILLER_204_899 ();
 sg13g2_decap_8 FILLER_204_906 ();
 sg13g2_decap_8 FILLER_204_913 ();
 sg13g2_decap_8 FILLER_204_920 ();
 sg13g2_decap_8 FILLER_204_927 ();
 sg13g2_decap_8 FILLER_204_934 ();
 sg13g2_decap_8 FILLER_204_941 ();
 sg13g2_decap_8 FILLER_204_948 ();
 sg13g2_decap_8 FILLER_204_955 ();
 sg13g2_decap_8 FILLER_204_962 ();
 sg13g2_decap_8 FILLER_204_969 ();
 sg13g2_decap_8 FILLER_204_976 ();
 sg13g2_decap_8 FILLER_204_983 ();
 sg13g2_decap_8 FILLER_204_990 ();
 sg13g2_decap_8 FILLER_204_997 ();
 sg13g2_decap_8 FILLER_204_1004 ();
 sg13g2_decap_8 FILLER_204_1011 ();
 sg13g2_decap_8 FILLER_204_1018 ();
 sg13g2_decap_8 FILLER_204_1025 ();
 sg13g2_decap_8 FILLER_204_1032 ();
 sg13g2_decap_8 FILLER_204_1039 ();
 sg13g2_decap_8 FILLER_204_1046 ();
 sg13g2_decap_8 FILLER_204_1053 ();
 sg13g2_decap_8 FILLER_204_1060 ();
 sg13g2_decap_8 FILLER_204_1067 ();
 sg13g2_decap_8 FILLER_204_1074 ();
 sg13g2_decap_8 FILLER_204_1081 ();
 sg13g2_decap_8 FILLER_204_1088 ();
 sg13g2_decap_8 FILLER_204_1095 ();
 sg13g2_decap_8 FILLER_204_1102 ();
 sg13g2_decap_8 FILLER_204_1109 ();
 sg13g2_decap_8 FILLER_204_1116 ();
 sg13g2_decap_8 FILLER_204_1123 ();
 sg13g2_decap_8 FILLER_204_1130 ();
 sg13g2_decap_8 FILLER_204_1137 ();
 sg13g2_decap_8 FILLER_204_1144 ();
 sg13g2_decap_8 FILLER_204_1151 ();
 sg13g2_decap_8 FILLER_204_1158 ();
 sg13g2_decap_8 FILLER_204_1165 ();
 sg13g2_decap_8 FILLER_204_1172 ();
 sg13g2_decap_8 FILLER_204_1179 ();
 sg13g2_decap_8 FILLER_204_1186 ();
 sg13g2_decap_8 FILLER_204_1193 ();
 sg13g2_decap_8 FILLER_204_1200 ();
 sg13g2_decap_8 FILLER_204_1207 ();
 sg13g2_decap_8 FILLER_204_1214 ();
 sg13g2_decap_8 FILLER_204_1221 ();
 sg13g2_decap_8 FILLER_204_1228 ();
 sg13g2_decap_8 FILLER_204_1235 ();
 sg13g2_decap_8 FILLER_204_1242 ();
 sg13g2_decap_8 FILLER_204_1249 ();
 sg13g2_decap_8 FILLER_204_1256 ();
 sg13g2_decap_8 FILLER_204_1263 ();
 sg13g2_decap_8 FILLER_204_1270 ();
 sg13g2_decap_8 FILLER_204_1277 ();
 sg13g2_decap_8 FILLER_204_1284 ();
 sg13g2_decap_8 FILLER_204_1291 ();
 sg13g2_decap_8 FILLER_204_1298 ();
 sg13g2_decap_8 FILLER_204_1305 ();
 sg13g2_decap_8 FILLER_204_1312 ();
 sg13g2_decap_8 FILLER_204_1319 ();
 sg13g2_decap_8 FILLER_204_1326 ();
 sg13g2_decap_8 FILLER_204_1333 ();
 sg13g2_decap_8 FILLER_204_1340 ();
 sg13g2_decap_8 FILLER_204_1347 ();
 sg13g2_decap_8 FILLER_204_1354 ();
 sg13g2_decap_8 FILLER_204_1361 ();
 sg13g2_decap_8 FILLER_204_1368 ();
 sg13g2_decap_8 FILLER_204_1375 ();
 sg13g2_decap_8 FILLER_204_1382 ();
 sg13g2_decap_8 FILLER_204_1389 ();
 sg13g2_decap_8 FILLER_204_1396 ();
 sg13g2_decap_8 FILLER_204_1403 ();
 sg13g2_decap_8 FILLER_204_1410 ();
 sg13g2_decap_8 FILLER_204_1417 ();
 sg13g2_decap_8 FILLER_204_1424 ();
 sg13g2_decap_8 FILLER_204_1431 ();
 sg13g2_decap_8 FILLER_204_1438 ();
 sg13g2_decap_8 FILLER_204_1445 ();
 sg13g2_decap_8 FILLER_204_1452 ();
 sg13g2_decap_8 FILLER_204_1459 ();
 sg13g2_decap_8 FILLER_204_1466 ();
 sg13g2_decap_8 FILLER_204_1473 ();
 sg13g2_decap_8 FILLER_204_1480 ();
 sg13g2_decap_8 FILLER_204_1487 ();
 sg13g2_decap_8 FILLER_204_1494 ();
 sg13g2_decap_8 FILLER_204_1501 ();
 sg13g2_decap_8 FILLER_204_1508 ();
 sg13g2_decap_8 FILLER_204_1515 ();
 sg13g2_decap_8 FILLER_204_1522 ();
 sg13g2_decap_8 FILLER_204_1529 ();
 sg13g2_decap_8 FILLER_204_1536 ();
 sg13g2_decap_8 FILLER_204_1543 ();
 sg13g2_decap_8 FILLER_204_1550 ();
 sg13g2_decap_8 FILLER_204_1557 ();
 sg13g2_decap_8 FILLER_204_1564 ();
 sg13g2_decap_8 FILLER_204_1571 ();
 sg13g2_decap_8 FILLER_204_1578 ();
 sg13g2_decap_8 FILLER_204_1585 ();
 sg13g2_decap_8 FILLER_204_1592 ();
 sg13g2_decap_8 FILLER_204_1599 ();
 sg13g2_decap_8 FILLER_204_1606 ();
 sg13g2_decap_8 FILLER_204_1613 ();
 sg13g2_decap_4 FILLER_204_1620 ();
 sg13g2_fill_1 FILLER_204_1624 ();
endmodule
