* Extracted by KLayout with SG13G2 LVS runset on : 12/09/2025 21:18

.SUBCKT asicone_202508 AVDD|anode|cathode|pad|vdd
+ anode|cathode|pad|pad_adc_rst_pad anode|cathode|pad|pad_adc_clk_pad
+ anode|cathode|pad|pad_adc_result_0_pad anode|cathode|pad|pad_adc_result_1_pad
+ anode|cathode|pad|pad_adc_result_2_pad anode|cathode|pad|pad_adc_result_3_pad
+ anode|cathode|pad|pad_adc_result_4_pad anode|cathode|pad|pad_adc_valid_pad
+ anode|cathode|pad|pad_adc_sample_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply VSSIO|anode|cathode|guard|iovss
+ gate|ngate|o gate|ngate|o$1 gate|ngate|o$2 gate|ngate|o$3 gate|ngate|o$4
+ gate|ngate|o$5 gate|ngate|o$6 gate|o|pgate gate|o|pgate$1 gate|o|pgate$2
+ gate|o|pgate$3 gate|o|pgate$4 gate|o|pgate$5 gate|o|pgate$6 core|padres core
+ core$1 VDD|pad|pin1|supply|vdd RESULT[0]|c2p|core|i|q RESULT[1]|c2p|core|i|q
+ RESULT[2]|c2p|core|i|q RESULT[3]|c2p|core|i|q RESULT[4]|c2p|core|i|q
+ VALID|a3|c2p|core|i|z SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|clk|vss
+ CLK|core|i|p2c anode|cathode|pad|pad_adc_go_pad i|z z zn z$1 z$2 i|z$1 z$3
+ z$4 i|z$2 z$5 GO|a2|core|p2c core$2 d|zn a2|zn a1|z b|zn z$6 zn$1 a1|z$1 d|z
+ b|zn$1 a1|z$2 a1|b|i|q a1|z$3 a2|z a2|a3|zn a1|b|i|q$1 a1|a2|a3|z d|zn$1
+ a2|zn$1 a1|z$4 d|z$1 cp|z a2 VIP|core|padres z$7 VIN|core|padres cp|z$1
+ anode|cathode|pad|pad_adc_vrefp_pad d|zn$2 VREFH|core|padres a2$1 z$8 z$9
+ a2|z$1 z$10 d|z$2 a2|z$2 a2|zn$2 a1|z$5 d|zn$3 b|zn$2 a1|z$6 a1|z$7
+ a1|b|i|q$2 d|zn$4 a1|z$8 d|zn$5 a1|z$9 a2|d|zn a2|zn$3 i|z$3 z$11 z$12 b|q
+ z$13 a2|i|q z$14 z$15 z$16 zn$2 d|z$3 z$17 z$18 z$19 a2|zn$4 z$20 d|zn$6
+ i|z$4 a1|b|i|q$3 a2|a3|z a1|z$10 b|zn$3 a2|z$3 a2|zn$5 in|pin2 a1|i|q
+ gate|out anode|cathode|pad|pad_adc_vrefn_pad i|zn i|z$5 i|z$6 i|z|zn i|z$7
+ z$21 i|z$8 cp|z$2 i|z$9 d|zn$7 i|z$10 i|z$11 i|z|zn$1 i|z$12 i|zn$1 i|z$13
+ i|z|zn$2 d|zn$8 i|z$14 i|z$15 VREFL|core|padres i|zn$2 i|z$16 i|z$17 i|z$18
+ i|z|zn$3 i|z$19 i|z$20 i|z$21 i|z$22 i|z|zn$4 i|z$23 a1|i|z|zn i|zn$3
+ i|z|zn$5 i|z$24 i|z|zn$6 i|z$25 i|z$26 i|z$27 i|z$28 i|z$29 i|zn$4 i|z$30
+ i|z$31 i|zn$5 i|z$32 a2|z$4 i|z$33 i|z$34 i|z$35 i|z$36 a1|z$11 i|zn$6 i|zn$7
+ i|z$37 i|z|zn$7 i|z$38 i|z|zn$8 i|z$39 i|z$40 i|z$41 a2|z$5 i|z$42 i|z$43
+ i|z$44 i|z$45 i|z$46 i|z$47 i|z$48 i|z$49 a1|i|q$1 i|z$50 i|z$51 a2|i|z
+ i|z$52 i|z$53 i|z$54 i|z$55 a1|c|i|zn z$22 z$23 i|z$56 i|zn$8 i|z$57 i|z$58
+ i|zn$9 i|zn$10 i|z$59 i|z$60 i|z$61 i|z$62 a2|b|z i|z$63 i|z$64 i|z$65 z$24
+ a1|c|i|zn$1 i|z$66 z$25 i|z$67 i|z$68 i|zn$11 i|z$69 i|z$70 i|z$71 i|z|zn$9
+ i|z$72 i|z$73 i|z$74 i|z$75 i|z$76 i|z$77 b|i|q i|z$78 i|z$79 b|i|q$1 i|z$80
+ i|z$81 i|z$82 i|z$83 i|z$84 i|z$85 i|z$86 a1|z$12 i|z$87 i|z$88 i|z$89 i|z$90
+ i|z$91 i|zn$12 i|z$92 i|z$93 i|z$94 i|z$95 b|i|q$2 i|z$96 i|z$97 i|zn$13
+ i|z$98 i|z$99 b|zn$4 cp|i|z zn$3 i|z$100 i|z$101 i|z$102 b|i|q$3 i|z$103
+ i|z$104 i|z$105 i|z$106 i|z$107 i|z$108 i|z$109 i|z$110 a2|zn$6 a1|z$13 zn$4
+ i|z$111 i|z$112 i|z$113 i|z$114 cp|z$3 d|zn$9 d|zn$10 a2|z$6
+ anode|cathode|pad|pad_adc_vin_pad b|zn$5 z$26 d|z$4 a2|z$7 b|zn$6 z$27 zn$5
+ gate|out$1 in|pin2$1 anode|cathode|pad|pad_adc_vip_pad
+ anode|cathode|pad|pad_miso_pad gate|o|pgate$7 DOUT_DAT|c2p|core|i|q
+ gate|ngate|o$7 s|zn s|z d|z$5 d|z$6 d|z$7 d|z$8 d|z$9 d|z$10 R[28]|i0|q
+ d|z$11 d|z$12 d|z$13 a1|a2|q a1|b|d|z d|z$14 a2|i|q$1 d|z$15 a1|a2|q$1 a2|q
+ a2|q$1 d|z$16 a1|a2|q$2 R[32]|i1|q i0|i1|q R[25]|i0|q cp|i|z$1 d|z$17 d|z$18
+ d|z$19 a3|zn R[27]|i0|q R[33]|i1|q i0|i1|q$1 a2|zn$7 d|z$20 d|z$21 d|z$22
+ a2|q$2 a1|a2|q$3 d|z$23 R[24]|i0|q R[34]|i1|q RST|a1|b|cdn|core|i|p2c
+ cp|i|z$2 d|z$24 a1|a2|q$4 a2|q$3 cp|i|z$3 R[26]|i0|q cp|i|z$4 d|z$25 d|z$26
+ d|z$27 d|z$28 a4|zn s|zn$1 z$28 d|z$29 a1|a2|q$5 a2|zn$8 a1|zn d|z$30 d|z$31
+ d|z$32 d|z$33 i0|i1|q$2 i|z$115 d|z$34 d|z$35 a2|zn$9 a2|q$4 a2|q$5
+ R[29]|i0|q R[36]|i1|q R[30]|i0|q i0|i1|q$3 a2|q$6 a2|zn$10 a1|i0|q
+ a1|i|i0|i1|q z$29 R[21]|i0|q d|z$36 z$30 R[20]|i0|q d|z$37 R[37]|i1|q
+ i0|i1|q$4 i0|i1|q$5 i0|i1|q$6 cp|z$4 d|z$38 a1|a2|q$6 a3|zn$1 a1|z$14 a4|zn$1
+ d|z$39 i0|i1|q$7 d|z$40 d|z$41 d|z$42 R[39]|i1|q d|z$43
+ anode|cathode|pad|pad_mosi_pad anode|cathode|pad|pad_RO_RST_B_pad d|s|zn z$31
+ a1|a2|q$7 d|s|z d|z$44 a2|i|s|zn a2|i|i0|i1|q R[18]|i0|q R[23]|i0|q d|z$45
+ R[53]|i1|q a1|i0|q$1 d|z$46 d|z$47 d|z$48 R[35]|i1|q d|z$49 d|z$50 a2|i|q$2
+ R[22]|i0|q d|z$51 s|zn$2 s|zn$3 a1|a2|q$8 d|z$52 a2|z$8 a1|zn$1 a1|a3|i|i1|q
+ R[50]|i1|q R[31]|i0|q R[17]|i0|q R[19]|i0|q R[38]|i1|q d|z$53 d|z$54 cp|i|z$5
+ a2|q$7 a4|zn$2 d|z$55 d|z$56 d|z$57 d|z$58 d|z$59 R[49]|i1|q d|z$60
+ R[51]|i1|q a1|a2|a4|z a1|a2|q$9 a1|a2|b|q|s R[54]|i1|q d|z$61 d|z$62
+ R[48]|i1|q R[55]|i1|q d|z$63 d|z$64 a2|zn$11 cp|i|z$6 d|z$65 a2|a3|zn$1
+ a2|z$9 R[52]|i1|q R[16]|i0|q d|z$66 d|z$67 s|z$1 s|zn$4 s|zn$5 s|zn$6 a3|zn$2
+ d|z$68 a1|zn$2 d|z$69 d|z$70 z$32 i1|z a2|zn$12 d|z$71 d|z$72 d|z$73 d|z$74
+ d|z$75 R[63]|i1|q R[47]|i0|q R[15]|i|i0|q R[12]|i|i0|q a2|a3|z$1 i0|z
+ CEB|a1|core|i|p2c R[7]|i|i0|q a1|z$15 CLK|core|i|p2c$1 cp|i|z$7 R[4]|i|i0|q
+ R[44]|i0|q i0|i1|q$8 i0|z$1 i1|z$1 d|z$76 z$33 a2|q$8 DOUT_EN|z R[43]|i0|q
+ R[46]|i0|q d|z$77 i0|i1|q$9 a2|d|z a2|z$10 d|z$78 d|z$79 R[60]|i1|q core$3
+ i0|i1|q$10 d|z$80 a2|zn$13 d|z$81 d|z$82 i1|z$2 RO_control|R[1]|i|i0|nclk|q
+ d|z$83 R[59]|i1|q DUT_Header|R[3]|Vup|i|i0|q R[14]|i|i0|q
+ R[0]|clk|i|i0|n_RO_control|q RESET_B|RSTB|core|p2c d|z$84 a2|zn$14 d|z$85
+ d|z$86 d|z$87 d|z$88 d|z$89 DATA|core|i0|i1|p2c core$4 d|z$90 i0|i1|q$11
+ i0|z$2 i0|z$3 d|z$91 R[58]|i1|q a1|zn$3 a1|zn$4 a2|zn$15 a1|zn$5 a2|z$11
+ a1|z$16 a2|zn$16 a2|zn$17 a3|zn$3 a1|z$17 a4|z d|z$92 d|z$93 d|z$94 d|z$95
+ i1|z$3 a1|i0|q$2 a2|zn$18 RD[39]|a2|z RD[28]|a2|z a2|zn$19 RD[33]|a2|z
+ RD[1]|a2|z a1|a3|z RD[29]|a2|zn RD[36]|a2|z RD[35]|a2|z R[6]|i|i0|q
+ R[40]|i0|q R[45]|i0|q R[57]|i1|q a3|zn$4 i0|i1|q$12 d|z$96 i0|z$4 R[61]|i1|q
+ a1|zn$6 a4|zn$3 a1|zn$7 a2|zn$20 a4|zn$4 a2|zn$21 i1|zn a1|zn$8 a1|zn$9
+ a4|z$1 a3|zn$5 a2|zn$22 a2|zn$23 a1|zn$10 a2|zn$24 z$34
+ DUT_Footer|R[2]|Vdn|i|i0|q R[41]|i0|q d|z$97 d|z$98 RD[7]|a2|zn i0|z$5
+ i0|i1|q$13 RD[25]|a2|zn a2|z$12 d|z$99 i1|zn$1 d|z$100 d|z$101 RD[4]|a2|z
+ RD[43]|a4|z RD[12]|a4|zn a4|zn$5 RD[19]|a4|z RD[17]|a4|z RD[23]|a4|z a2|zn$25
+ RD[9]|a4|z RD[46]|a4|z RD[38]|a2|z d|z$102 R[56]|i1|q d|z$103 R[62]|i1|q
+ i1|zn$2 a1|zn$11 a1|i1|q R[5]|i|i0|q a3|zn$6 a3|zn$7 a2|zn$26 a1|zn$12
+ a2|zn$27 a1|zn$13 a4|zn$6 a3|zn$8 R[13]|i|i0|q R[42]|i0|q d|z$104 d|z$105
+ d|z$106 RD[40]|a4|z RD[20]|a4|zn RD[16]|a4|zn RD[44]|a4|z RD[18]|a4|zn
+ a2|zn$28 a4|zn$7 RD[0]|a2|z RD[15]|a4|zn RD[22]|a4|zn RD[13]|a4|zn a4|zn$8
+ a2|z$13 RD[30]|a2|z RD[45]|a4|z d|z$107 d|z$108 DUT_Header|R[11]|Vup|i|i0|q
+ R[8]|clk|i|i0|n_RO_control|q RO_control|R[9]|i|i0|nclk|q b|z a2|zn$29
+ a1|zn$14 a2|zn$30 a1|zn$15 a3|zn$9 a2|zn$31 a1|zn$16 a2|zn$32 a1|zn$17
+ a1|zn$18 a1|zn$19 a3|zn$10 a2|zn$33 a2|zn$34 a3|zn$11 a1|zn$20 a2|zn$35
+ a1|zn$21 a1|zn$22 a1|zn$23 i0|z$6 RD[34]|a2|z RD[26]|a2|z RD[37]|a2|z
+ RD[31]|a2|zn RD[14]|a4|zn RD[32]|a2|z RD[2]|a2|z RD[10]|a4|zn RD[11]|a4|zn
+ RD[8]|a4|z RD[24]|a2|z RD[27]|a2|zn RD[21]|a4|z RD[47]|a4|z RD[3]|a2|z
+ RD[5]|a2|zn RD[6]|a2|zn Vin Vin|Vout|core|extra_load|padres
+ Drain_Sense|Vout|core|padres Drain_Force|Vout|core|padres Vout IN|Vout Vin$1
+ Vin$2 DUT_Footer|R[10]|Vdn|i|i0|q Vin|Vout D|Q_N Q D|Q_N$1 Q$1 D|Q_N$2 Q$2
+ D|Q_N$3 Q$3 D|Q_N$4 OUT|Q|c2p|core|i RO2VDD|VDD|anode|cathode|nclk|pad Vin$3
+ Vin$4 Vout$1 Vin$5 Vin$6 Vout$2 Vin$7 Vin$8 Vout$3 Vin$9 Vin$10 Vout$4 Vin$11
+ Vin$12 Vout$5 Vin$13 Vin$14 Vout$6 Vin$15 Vin$16 Vout$7 Vin$17 Vin$18 Vout$8
+ Vin$19 Vin$20 anode|cathode|pad|pad_sclk_pad
+ anode|cathode|pad|pad_RO_101_DUT_gate_pad RD[42]|a4|z RD[41]|a4|z i i$1 i$2
+ i$3 i$4 core$5 DUT_gate|core|p2c core$6 anode|cathode|pad|pad_cs_pad
+ anode|cathode|pad|pad_RO_13_DUT_gate_pad Vin|Vout|core|extra_load|padres$1
+ Vin$21 Vin$22 Vin$23 Vin$24 Vin$25 Vin$26 Vin$27 Vin$28 Vin$29 Vin$30 Vin$31
+ Vin$32 Vin$33 Vin$34 Vin$35 Vin$36 Vin$37 Vin$38 Vin$39 Vin$40 Vin$41 Vin$42
+ Vin$43 Vin$44 Vin$45 Vin$46 Vin$47 Vin$48 Vin$49 Vin$50 Vin$51 Vin$52 Vin$53
+ Vin$54 Vin$55 Vin$56 Vin$57 Vin$58 Vin$59 Vin$60 Vin$61 Vin$62 Vin$63 Vin$64
+ Vin$65 Vin$66 Vin$67 Vin$68 Vin$69 Vin$70 Vin$71 Vin$72 Vin$73 Vin$74 Vin$75
+ Vin$76 Vin$77 Vin$78 Vin$79 Vin$80 Vin$81 Vin$82 Vin$83 Vin$84 Vin$85 Vin$86
+ Vin$87 Vin$88 Vin$89 Vin$90 Vin$91 Vin$92 Vin$93 Vin$94 Vin$95 Vin$96 Vin$97
+ Vin$98 Vin$99 Vin$100 Vin$101 Vin$102 Vin$103 Vin$104 Vout$9 Vin$105 Vin$106
+ Vin$107 Drain_Sense|Vout|core|padres$1 Drain_Force|Vout|core|padres$1
+ IN|Vin|Vout Vin$108 Vin$109 Vin|Vout$1 Vin|Vout$2 Vin|Vout$3 Vin|Vout$4
+ Vin|Vout$5 Vin|Vout$6 Vin|Vout$7 Vin|Vout$8 Vin|Vout$9 Vin|Vout$10
+ Vin|Vout$11 Vin|Vout$12 Vin|Vout$13 Vin|Vout$14 Vin|Vout$15 Vin|Vout$16
+ Vin|Vout$17 Vin|Vout$18 Vin|Vout$19 Vin|Vout$20 Vin|Vout$21 Vin|Vout$22
+ Vin|Vout$23 Vin|Vout$24 Vin|Vout$25 Vin|Vout$26 Vin|Vout$27 Vin|Vout$28
+ Vin|Vout$29 Vin|Vout$30 Vin|Vout$31 Vin|Vout$32 Vin|Vout$33 Vin|Vout$34
+ Vin|Vout$35 Vin|Vout$36 Vin|Vout$37 Vin|Vout$38 Vin|Vout$39 Vin|Vout$40
+ Vin|Vout$41 Vin|Vout$42 Vin|Vout$43 Vin$110 ROVDD|VDD|anode|cathode|nclk|pad
+ Vin$111 Vin$112 Vin|Vout$44 Vin$113 Vin$114 Vin|Vout$45 Vin$115 Vin$116
+ Vin|Vout$46 Vin$117 Vin$118 Vin|Vout$47 Vin$119 Vin$120 Vin|Vout$48 Vin$121
+ Vin$122 Vin|Vout$49 Vin$123 Vin$124 Vin|Vout$50 Vin$125 Vin$126 Vin|Vout$51
+ Vin$127 Vin$128 Vin|Vout$52 Vin$129 Vin$130 Vin|Vout$53 Vin$131 Vin$132
+ Vin|Vout$54 Vin$133 Vin$134 Vin|Vout$55 Vin$135 Vin$136 Vin|Vout$56 Vin$137
+ Vin$138 Vin|Vout$57 Vin$139 Vin$140 Vin|Vout$58 Vin$141 Vin$142 Vin|Vout$59
+ Vin$143 Vin$144 Vin|Vout$60 Vin$145 Vin$146 Vin|Vout$61 Vin$147 Vin$148
+ Vin|Vout$62 Vin$149 Vin$150 Vin|Vout$63 Vin$151 Vin$152 Vin|Vout$64 Vin$153
+ Vin$154 Vin|Vout$65 Vin$155 Vin$156 Vin|Vout$66 Vin$157 Vin$158 Vin|Vout$67
+ Vin$159 Vin$160 Vin|Vout$68 Vin$161 Vin$162 Vin|Vout$69 Vin$163 Vin$164
+ Vin|Vout$70 Vin$165 Vin$166 Vin|Vout$71 Vin$167 Vin$168 Vin|Vout$72 Vin$169
+ Vin$170 Vin|Vout$73 Vin$171 Vin$172 Vin|Vout$74 Vin$173 Vin$174 Vin|Vout$75
+ Vin$175 Vin$176 Vin|Vout$76 Vin$177 Vin$178 Vin|Vout$77 Vin$179 Vin$180
+ Vin|Vout$78 Vin$181 Vin$182 Vin|Vout$79 Vin$183 Vin$184 Vin|Vout$80 Vin$185
+ Vin$186 Vin|Vout$81 Vin$187 Vin$188 Vin|Vout$82 Vin$189 Vin$190 Vin|Vout$83
+ Vin$191 Vin$192 Vin|Vout$84 Vin$193 Vin$194 Vin|Vout$85 Vin$195 Vin$196
+ Vin|Vout$86 Vin$197 Vin$198 Vin|Vout$87 Vin$199 Vin$200 Vin|Vout$88 Vin$201
+ Vin$202 Vin|Vout$89 Vin$203 Vin$204 Vin|Vout$90 Vin$205 Vin$206 Vin|Vout$91
+ Vin$207 Vin$208 Vin|Vout$92 Vin$209 Vin$210 Vin|Vout$93 Vin$211 Vin$212
+ Vin|Vout$94 Vin$213 Vin$214 Vin|Vout$95 Vin$215 Vin$216 Vin|Vout$96 Vin$217
+ Vin$218 core$7 OUT|Q|c2p|core|i$1 D|Q_N$5 D|Q_N$6 D|Q_N$7 D|Q_N$8 D|Q_N$9
+ DUT_gate|core|p2c$1 Q$4 Q$5 Q$6 Q$7 core$8
+ anode|cathode|pad|pad_RO_101_Drain_Force_pad
+ anode|cathode|pad|pad_RO_101_Drain_Sense_pad
+ anode|cathode|pad|pad_RO_101_extra_load_pad
+ anode|cathode|pad|pad_RO_13_Drain_Force_pad
+ anode|cathode|pad|pad_RO_13_Drain_Sense_pad
+ anode|cathode|pad|pad_RO_13_extra_load_pad core|padres$1 core|padres$2
+ gate|o|pgate$8 gate|ngate|o$8 gate|o|pgate$9 gate|ngate|o$9
+ anode|cathode|pad|pad_RO_101_Vout_pad anode|cathode|pad|pad_RO_13_Vout_pad
M$1 RST|a1|b|cdn|core|i|p2c \$64422 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$2 CLK|core|i|p2c \$64424 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$3 \$63550 RESULT[0]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$4 \$63551 RESULT[0]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$5 \$63553 RESULT[1]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$6 \$63554 RESULT[1]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$7 \$63556 RESULT[2]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$8 \$63557 RESULT[2]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$9 \$63559 RESULT[3]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$10 \$63560 RESULT[3]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$11 \$63562 RESULT[4]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$12 \$63563 RESULT[4]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$13 \$63565 VALID|a3|c2p|core|i|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$14 \$63566 VALID|a3|c2p|core|i|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$15 \$63568 SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$16 \$63569 SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$17 \$89657 \$89973 \$89657 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$53 \$89658 \$89974 \$89658 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$89 \$89659 \$89975 \$89659 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$125 \$89660 \$89976 \$89660 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$161 \$89661 \$89977 \$89661 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$197 \$89662 \$89978 \$89662 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$233 \$89663 \$89979 \$89663 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$269 \$89664 \$89980 \$89664 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$305 \$89665 \$89981 \$89665 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$341 \$89666 \$89982 \$89666 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$737 VSS|anode|cathode|clk|vss a2|zn \$92658 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$738 \$92658 a1|z d|zn VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$739 d|zn b|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$740 GO|a2|core|p2c \$90525 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$741 \$94761 \$95239 \$94761 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$753 \$92959 z$6 \$92959 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$754 \$89973 zn$1 \$92959 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$755 \$89973 z$6 \$89973 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$770 \$92960 zn$1 \$89973 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$771 \$92960 z$6 \$92960 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$786 \$92961 zn$1 \$89973 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$787 \$92961 z$6 \$92961 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$789 \$94762 \$95240 \$94762 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=829.44u AS=354.5856p AD=354.5856p PS=1883.52u PD=1883.52u
M$801 \$92962 z$6 \$92962 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$802 \$89974 zn$1 \$92962 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$803 \$89974 z$6 \$89974 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$818 \$92963 zn$1 \$89974 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$819 \$92963 z$6 \$92963 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$834 \$92964 zn$1 \$89974 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$835 \$92964 z$6 \$92964 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$849 \$92965 z$6 \$92965 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$850 \$89975 zn$1 \$92965 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$851 \$89975 z$6 \$89975 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$866 \$92966 zn$1 \$89975 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$867 \$92966 z$6 \$92966 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$882 \$92967 zn$1 \$89975 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$883 \$92967 z$6 \$92967 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$897 \$92968 z$6 \$92968 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$898 \$89976 zn$1 \$92968 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$899 \$89976 z$6 \$89976 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$914 \$92969 zn$1 \$89976 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$915 \$92969 z$6 \$92969 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$930 \$92970 zn$1 \$89976 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$931 \$92970 z$6 \$92970 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$945 \$92971 z$6 \$92971 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$946 \$89977 zn$1 \$92971 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$947 \$89977 z$6 \$89977 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$962 \$92972 zn$1 \$89977 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$963 \$92972 z$6 \$92972 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$978 \$92973 zn$1 \$89977 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$979 \$92973 z$6 \$92973 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$993 \$92974 z$6 \$92974 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$994 \$89978 zn$1 \$92974 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$995 \$89978 z$6 \$89978 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1010 \$92975 zn$1 \$89978 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1011 \$92975 z$6 \$92975 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1026 \$92976 zn$1 \$89978 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1027 \$92976 z$6 \$92976 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1041 \$92977 z$6 \$92977 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1042 \$89979 zn$1 \$92977 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1043 \$89979 z$6 \$89979 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1058 \$92978 zn$1 \$89979 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1059 \$92978 z$6 \$92978 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1074 \$92979 zn$1 \$89979 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1075 \$92979 z$6 \$92979 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1089 \$92980 z$6 \$92980 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1090 \$89980 zn$1 \$92980 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1091 \$89980 z$6 \$89980 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1106 \$92981 zn$1 \$89980 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1107 \$92981 z$6 \$92981 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1122 \$92982 zn$1 \$89980 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1123 \$92982 z$6 \$92982 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1137 \$92983 z$6 \$92983 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1138 \$89981 zn$1 \$92983 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1139 \$89981 z$6 \$89981 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1154 \$92984 zn$1 \$89981 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1155 \$92984 z$6 \$92984 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1170 \$92985 zn$1 \$89981 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1171 \$92985 z$6 \$92985 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1173 \$94763 \$95241 \$94763 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$1185 \$92986 z$6 \$92986 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1186 \$89982 zn$1 \$92986 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1187 \$89982 z$6 \$89982 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1202 \$92987 zn$1 \$89982 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1203 \$92987 z$6 \$92987 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1218 \$92988 zn$1 \$89982 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1219 \$92988 z$6 \$92988 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1581 \$94525 a1|z$3 \$95372 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$1582 VSS|anode|cathode|clk|vss a2|z \$95372 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.655u AS=0.2901875p AD=0.271825p PS=1.55u PD=1.485u
M$1583 VSS|anode|cathode|clk|vss \$94525 d|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2901875p AD=0.4068p PS=1.55u PD=2.57u
M$1584 b|zn$1 a1|a2|a3|z \$95374 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$1585 \$95374 GO|a2|core|p2c \$95375 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$1586 \$95375 a2|a3|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$1587 VSS|anode|cathode|clk|vss a2|zn$1 \$96161 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$1588 \$96161 a1|z$4 d|zn$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$1589 d|zn$1 b|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$1590 a1|z$1 a1|b|i|q$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$1591 a1|z$2 a1|b|i|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$1592 \$100188 \$100549 \$100188 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$1604 \$98170 z$6 \$98170 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1605 \$95239 zn$1 \$98170 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1606 \$95239 z$6 \$95239 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1621 \$98171 zn$1 \$95239 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1622 \$98171 z$6 \$98171 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1637 \$98172 zn$1 \$95239 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1638 \$98172 z$6 \$98172 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1652 a2 z$3 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1653 \$95240 z$1 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=11.52u
+ AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$1654 \$95240 z$3 \$95240 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1668 \$95240 z$7 \$95240 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1669 VIP|core|padres z$4 \$95240 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$1670 VIP|core|padres z$7 VIP|core|padres VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1684 \$95240 z$2 \$95240 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1685 VIN|core|padres zn \$95240 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$1686 VIN|core|padres z$2 VIN|core|padres VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1736 \$100189 \$100550 \$100189 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=414.72u AS=177.2928p AD=177.2928p PS=941.76u PD=941.76u
M$2024 \$100190 \$100551 \$100190 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$2036 \$98175 z$6 \$98175 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2037 \$95241 zn$1 \$98175 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2038 \$95241 z$6 \$95241 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$2053 \$98176 zn$1 \$95241 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2054 \$98176 z$6 \$98176 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2069 \$98177 zn$1 \$95241 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2070 \$98177 z$6 \$98177 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2072 \$97466 \$97411 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$2073 VSS|anode|cathode|clk|vss cp|z \$97411 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$2074 \$99070 \$98923 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$2075 VSS|anode|cathode|clk|vss cp|z$1 \$98923 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$2076 VSS|anode|cathode|clk|vss \$97411 \$98656 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$2077 \$98656 d|z$1 \$97412 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$2078 \$97412 \$97466 \$98657 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$2079 VSS|anode|cathode|clk|vss \$97467 \$98657 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$2080 VSS|anode|cathode|clk|vss \$97412 \$97467 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$2081 \$97467 \$97466 \$98590 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$2082 \$98590 \$97411 \$98658 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$2083 VSS|anode|cathode|clk|vss \$98130 \$98658 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$2084 VSS|anode|cathode|clk|vss \$98590 \$98130 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$2085 \$98924 \$99070 \$99259 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$2086 \$99259 \$98926 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$2087 \$98925 \$98923 \$99248 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$2088 \$99248 \$99071 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$2089 \$98926 \$99070 \$98925 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$2090 VSS|anode|cathode|clk|vss \$98923 \$99258 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$2091 \$99258 d|zn$1 \$98924 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$2092 VSS|anode|cathode|clk|vss \$98924 \$98926 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$2093 VSS|anode|cathode|clk|vss \$98925 \$99071 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$2094 b|i|q$1 \$98130 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$2095 RESULT[3]|c2p|core|i|q \$99071 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$2456 \$102321 \$102317 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$2457 VSS|anode|cathode|clk|vss cp|z$1 \$102317 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$2458 \$102318 \$102321 \$102586 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$2459 \$102586 \$102322 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$2460 \$102319 \$102317 \$102582 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$2461 \$102582 \$102599 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$2462 \$102322 \$102321 \$102319 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$2463 VSS|anode|cathode|clk|vss \$102317 \$102585 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$2464 \$102585 d|zn$2 \$102318 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$2465 VSS|anode|cathode|clk|vss \$102318 \$102322 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$2466 VSS|anode|cathode|clk|vss \$102319 \$102599 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$2467 RESULT[0]|c2p|core|i|q \$102599 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$2468 \$104013 z$6 \$104013 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2469 \$100549 zn$1 \$104013 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2470 \$100549 z$6 \$100549 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$2473 \$104014 zn$1 \$100549 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2474 \$104014 z$6 \$104014 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2477 \$104015 zn$1 \$100549 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2478 \$104015 z$6 \$104015 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2504 VREFH|core|padres z$7 VREFH|core|padres VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$2505 \$100550 z$4 VREFH|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$2506 \$100550 z$7 \$100550 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$2508 \$100550 z$9 \$100550 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$2509 a2 z \$100550 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$2510 a2 z$9 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$2512 \$100550 z$8 \$100550 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$2513 a2$1 z$5 \$100550 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$2514 a2$1 z$8 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$2576 \$104018 z$6 \$104018 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2577 \$100551 zn$1 \$104018 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2578 \$100551 z$6 \$100551 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$2581 \$104019 zn$1 \$100551 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2582 \$104019 z$6 \$104019 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2585 \$104020 zn$1 \$100551 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2586 \$104020 z$6 \$104020 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2588 VSS|anode|cathode|clk|vss a2|z$2 \$105732 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$2589 \$105732 a1|i|q b|zn VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$2590 b|zn RST|a1|b|cdn|core|i|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p
+ PS=1.55u PD=2.57u
M$2591 \$105439 a1|z$3 \$105735 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$2592 \$105735 a2|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.655u AS=0.271825p AD=0.2901875p PS=1.485u PD=1.55u
M$2593 VSS|anode|cathode|clk|vss \$105439 d|z$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2901875p AD=0.4068p PS=1.55u PD=2.57u
M$2594 VSS|anode|cathode|clk|vss a2|zn$2 \$105734 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$2595 \$105734 a1|z$5 d|zn$3 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$2596 d|zn$3 b|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$2597 \$105761 \$106210 \$105761 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$2705 \$105762 \$106211 \$105762 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=207.36u AS=88.6464p AD=88.6464p PS=470.88u PD=470.88u
M$2921 \$105763 \$106212 \$105763 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$3317 a1|z$5 RESULT[2]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$3318 b|zn$2 a1|z$7 \$108127 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$3319 \$108127 a2|i|q \$108128 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$3320 \$108128 a1|a2|a3|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$3321 \$107103 \$106574 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$3322 VSS|anode|cathode|clk|vss cp|z \$106574 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$3323 VSS|anode|cathode|clk|vss \$106574 \$108122 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$3324 \$108122 d|z \$106575 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$3325 \$106575 \$107103 \$108123 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$3326 VSS|anode|cathode|clk|vss \$107104 \$108123 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$3327 VSS|anode|cathode|clk|vss \$106575 \$107104 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$3328 \$107104 \$107103 \$107535 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$3329 \$107535 \$106574 \$108124 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$3330 VSS|anode|cathode|clk|vss \$107450 \$108124 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$3331 VSS|anode|cathode|clk|vss \$107535 \$107450 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$3332 b|i|q \$107450 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$3333 a1|z$6 a1|b|i|q$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$3334 \$110666 \$111316 \$110666 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$3346 \$108873 z$6 \$108873 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3347 \$106210 zn$1 \$108873 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3348 \$106210 z$6 \$106210 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$3363 \$108874 zn$1 \$106210 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3364 \$108874 z$6 \$108874 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3379 \$108875 zn$1 \$106210 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3380 \$108875 z$6 \$108875 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3478 \$110667 \$111317 \$110667 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=103.68u AS=44.3232p AD=44.3232p PS=235.44u PD=235.44u
M$3491 \$106211 z$4 VREFH|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$3492 \$106211 z$7 \$106211 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$3506 \$106211 z$12 \$106211 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$3507 a2 z$11 \$106211 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$3508 a2 z$12 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$3522 \$106211 z$10 \$106211 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$3523 a2$1 z$13 \$106211 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$3524 a2$1 z$10 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$3526 \$110668 \$111318 \$110668 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$3574 \$110669 \$111319 \$110669 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$3766 \$110670 \$111320 \$110670 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$3778 \$108876 z$6 \$108876 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3779 \$106212 zn$1 \$108876 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3780 \$106212 z$6 \$106212 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$3795 \$108877 zn$1 \$106212 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3796 \$108877 z$6 \$108877 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3811 \$108878 zn$1 \$106212 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3812 \$108878 z$6 \$108878 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3814 \$109960 \$109381 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$3815 VSS|anode|cathode|clk|vss cp|z \$109381 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$3816 VSS|anode|cathode|clk|vss \$109381 \$111115 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$3817 \$111115 d|z$2 \$109382 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$3818 \$109382 \$109960 \$111114 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$3819 VSS|anode|cathode|clk|vss \$109383 \$111114 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$3820 VSS|anode|cathode|clk|vss \$109382 \$109383 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$3821 \$109383 \$109960 \$110568 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$3822 \$110568 \$109381 \$111099 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$3823 VSS|anode|cathode|clk|vss \$109961 \$111099 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$3824 VSS|anode|cathode|clk|vss \$110568 \$109961 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$3825 a1|z$8 RESULT[1]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$3826 \$108454 a2|d|zn d|zn$4 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$3827 d|zn$4 a1|z$9 \$108454 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$3828 \$108454 b|zn$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$3829 \$108455 a2|zn$3 d|zn$5 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$3830 d|zn$5 a1|z$6 \$108455 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$3831 \$108455 b|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$3832 b|q \$109961 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$3833 \$108456 i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$3834 VSS|anode|cathode|clk|vss \$108456 cp|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$4195 a1|a2|a3|z RST|a1|b|cdn|core|i|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$4196 \$111321 i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$4197 VSS|anode|cathode|clk|vss \$111321 cp|z$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$4198 \$111624 \$111123 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$4199 VSS|anode|cathode|clk|vss cp|z$1 \$111123 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$4200 \$111124 \$111624 \$111538 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$4201 \$111538 \$111322 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$4202 \$111125 \$111123 \$111542 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$4203 \$111542 \$111626 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$4204 \$111322 \$111624 \$111125 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$4205 VSS|anode|cathode|clk|vss \$111123 \$111625 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$4206 \$111625 d|zn \$111124 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$4207 VSS|anode|cathode|clk|vss \$111124 \$111322 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$4208 VSS|anode|cathode|clk|vss \$111125 \$111626 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$4209 RESULT[4]|c2p|core|i|q \$111626 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$4210 \$114146 z$6 \$114146 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4211 \$111316 zn$1 \$114146 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4212 \$111316 z$6 \$111316 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$4215 \$114147 zn$1 \$111316 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4216 \$114147 z$6 \$114147 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4219 \$114148 zn$1 \$111316 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4220 \$114148 z$6 \$114148 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4247 \$111317 z$4 VREFH|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$4248 \$111317 z$7 \$111317 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4250 \$111317 z$14 \$111317 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4251 a2 z$15 \$111317 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$4252 a2 z$14 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4254 \$111317 z$18 \$111317 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4255 a2$1 z$19 \$111317 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$4256 a2$1 z$18 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4259 \$111318 z$4 VREFH|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4260 \$111318 z$7 \$111318 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4262 \$111318 z$16 \$111318 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4263 a2 z$25 \$111318 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4264 a2 z$16 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4266 \$111318 z$21 \$111318 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4267 a2$1 z$23 \$111318 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4268 a2$1 z$21 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4271 \$111319 z$4 VREFH|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4272 \$111319 z$7 \$111319 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4274 \$111319 z$17 \$111319 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4275 a2 zn$2 \$111319 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4276 a2 z$17 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4279 a2$1 zn$2 \$111319 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4280 a2$1 z$17 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4318 \$114150 z$6 \$114150 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4319 \$111320 zn$1 \$114150 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4320 \$111320 z$6 \$111320 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$4323 \$114151 zn$1 \$111320 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4324 \$114151 z$6 \$114151 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4327 \$114152 zn$1 \$111320 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4328 \$114152 z$6 \$114152 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4330 \$114426 \$114135 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$4331 VSS|anode|cathode|clk|vss cp|z \$114135 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$4332 \$114136 \$114426 \$114360 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$4333 \$114360 \$114153 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$4334 \$114137 \$114135 \$114354 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$4335 \$114354 \$114513 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$4336 \$114153 \$114426 \$114137 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$4337 VSS|anode|cathode|clk|vss \$114135 \$114464 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$4338 \$114464 d|z$3 \$114136 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$4339 VSS|anode|cathode|clk|vss \$114136 \$114153 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$4340 VSS|anode|cathode|clk|vss \$114137 \$114513 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$4341 \$112921 a1|z$7 \$113782 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$4342 VSS|anode|cathode|clk|vss a2|i|q \$113782 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.655u AS=0.2901875p AD=0.271825p PS=1.55u PD=1.485u
M$4343 VSS|anode|cathode|clk|vss \$112921 SAMPLE|a1|c2p|core|i|z
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2901875p
+ AD=0.4068p PS=1.55u PD=2.57u
M$4344 b|i|q$3 \$114513 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$4345 \$115923 \$116062 \$115923 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4381 \$115924 \$116063 \$115924 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4417 \$115925 \$116064 \$115925 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4453 \$115926 \$116065 \$115926 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4489 \$115927 \$116066 \$115927 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4525 \$115928 \$116067 \$115928 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4561 \$115929 \$116068 \$115929 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4597 \$115930 \$116069 \$115930 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4633 \$115931 \$116070 \$115931 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4669 \$115932 \$116071 \$115932 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$5065 \$119299 z$6 \$119299 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5066 \$116062 zn$1 \$119299 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5067 \$116062 z$6 \$116062 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5070 \$119300 zn$1 \$116062 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5071 \$119300 z$6 \$119300 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5074 \$119301 zn$1 \$116062 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5075 \$119301 z$6 \$119301 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5077 \$119302 z$6 \$119302 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5078 \$116063 zn$1 \$119302 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5079 \$116063 z$6 \$116063 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5082 \$119303 zn$1 \$116063 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5083 \$119303 z$6 \$119303 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5086 \$119304 zn$1 \$116063 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5087 \$119304 z$6 \$119304 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5089 \$119305 z$6 \$119305 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5090 \$116064 zn$1 \$119305 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5091 \$116064 z$6 \$116064 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5094 \$119306 zn$1 \$116064 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5095 \$119306 z$6 \$119306 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5098 \$119307 zn$1 \$116064 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5099 \$119307 z$6 \$119307 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5101 \$119308 z$6 \$119308 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5102 \$116065 zn$1 \$119308 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5103 \$116065 z$6 \$116065 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5106 \$119309 zn$1 \$116065 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5107 \$119309 z$6 \$119309 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5110 \$119310 zn$1 \$116065 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5111 \$119310 z$6 \$119310 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5113 \$119311 z$6 \$119311 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5114 \$116066 zn$1 \$119311 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5115 \$116066 z$6 \$116066 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5118 \$119312 zn$1 \$116066 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5119 \$119312 z$6 \$119312 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5122 \$119313 zn$1 \$116066 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5123 \$119313 z$6 \$119313 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5125 \$119314 z$6 \$119314 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5126 \$116067 zn$1 \$119314 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5127 \$116067 z$6 \$116067 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5130 \$119315 zn$1 \$116067 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5131 \$119315 z$6 \$119315 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5134 \$119316 zn$1 \$116067 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5135 \$119316 z$6 \$119316 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5137 \$119317 z$6 \$119317 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5138 \$116068 zn$1 \$119317 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5139 \$116068 z$6 \$116068 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5142 \$119318 zn$1 \$116068 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5143 \$119318 z$6 \$119318 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5146 \$119319 zn$1 \$116068 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5147 \$119319 z$6 \$119319 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5149 \$119320 z$6 \$119320 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5150 \$116069 zn$1 \$119320 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5151 \$116069 z$6 \$116069 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5154 \$119321 zn$1 \$116069 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5155 \$119321 z$6 \$119321 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5158 \$119322 zn$1 \$116069 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5159 \$119322 z$6 \$119322 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5161 \$119323 z$6 \$119323 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5162 \$116070 zn$1 \$119323 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5163 \$116070 z$6 \$116070 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5166 \$119324 zn$1 \$116070 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5167 \$119324 z$6 \$119324 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5170 \$119325 zn$1 \$116070 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5171 \$119325 z$6 \$119325 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5173 \$119326 z$6 \$119326 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5174 \$116071 zn$1 \$119326 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5175 \$116071 z$6 \$116071 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5178 \$119327 zn$1 \$116071 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5179 \$119327 z$6 \$119327 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5182 \$119328 zn$1 \$116071 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5183 \$119328 z$6 \$119328 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5185 \$120240 a1|i|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$5186 \$120241 a1|i|q \$120242 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2511p AD=0.1494p PS=1.55u PD=1.19u
M$5187 \$120242 \$120240 \$120243 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.36u AS=0.1494p AD=0.1494p PS=1.19u PD=1.19u
M$5188 \$120243 \$120241 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.1494p AD=0.2511p PS=1.19u PD=1.55u
M$5189 VSS|anode|cathode|clk|vss a2|i|q \$120241 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.2511p PS=1.55u PD=1.55u
M$5190 VSS|anode|cathode|clk|vss \$120242 a2|a3|zn VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$5191 VSS|anode|cathode|clk|vss i|z$4 \$118852 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2511p AD=0.2034p PS=1.55u PD=1.85u
M$5192 VSS|anode|cathode|clk|vss \$118852 i|z$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$5193 a2|zn$4 a1|b|i|q$3 \$120183 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5194 \$120183 a1|a2|a3|z \$120184 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5195 \$120184 a2|a3|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5196 a2|z$2 a2|i|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$5197 a2|z$3 \$120244 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5198 VSS|anode|cathode|clk|vss b|i|q$2 \$120244 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5199 \$120244 a1|b|i|q$1 \$120994 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5200 \$120994 a2|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5201 \$120097 a2|zn$3 d|zn$6 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5202 d|zn$6 a1|z$10 \$120097 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5203 \$120097 b|zn$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5204 z$20 i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$5205 \$120245 a1|i|q \$120932 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$5206 \$120932 a2|i|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.655u AS=0.271825p AD=0.2901875p PS=1.485u PD=1.55u
M$5207 VSS|anode|cathode|clk|vss \$120245 VALID|a3|c2p|core|i|z
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2901875p
+ AD=0.4068p PS=1.55u PD=2.57u
M$5208 VSS|anode|cathode|clk|vss i|zn \$123934 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5210 VSS|anode|cathode|clk|vss \$123934 i|z$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5214 \$123935 i|z|zn$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5215 VSS|anode|cathode|clk|vss \$123605 \$123936 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5216 \$123605 \$123935 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5217 VSS|anode|cathode|clk|vss \$123936 i|z$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5218 VSS|anode|cathode|clk|vss i|z$6 \$123938 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5224 VSS|anode|cathode|clk|vss \$123938 i|z|zn VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5240 VSS|anode|cathode|clk|vss i|z$7 \$123941 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5246 VSS|anode|cathode|clk|vss \$123941 z$21 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5262 VSS|anode|cathode|clk|vss \$124161 i|z$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5264 VSS|anode|cathode|clk|vss i|z$8 \$124161 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5265 \$123943 \$123606 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5266 VSS|anode|cathode|clk|vss cp|z$2 \$123606 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5267 \$123607 \$123943 \$124075 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$5268 \$124075 \$123944 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$5269 \$123608 \$123606 \$124076 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$5270 \$124076 \$124164 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$5271 \$123944 \$123943 \$123608 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$5272 VSS|anode|cathode|clk|vss \$123606 \$124072 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$5273 \$124072 d|zn$7 \$123607 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$5274 VSS|anode|cathode|clk|vss \$123607 \$123944 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$5275 VSS|anode|cathode|clk|vss \$123608 \$124164 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$5276 RESULT[1]|c2p|core|i|q \$124164 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$5277 VSS|anode|cathode|clk|vss i|z$2 \$125722 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5279 VSS|anode|cathode|clk|vss \$125722 i|z$10 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5283 \$125724 i|z$10 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5284 VSS|anode|cathode|clk|vss \$125725 \$125726 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5285 VSS|anode|cathode|clk|vss \$125724 \$125725 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5286 VSS|anode|cathode|clk|vss \$125726 i|z$11 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5287 VSS|anode|cathode|clk|vss \$126465 i|z$109 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5289 VSS|anode|cathode|clk|vss i|z$14 \$126465 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5290 \$125728 i|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5296 VSS|anode|cathode|clk|vss \$125728 z$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5312 \$125729 i|zn$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5318 VSS|anode|cathode|clk|vss \$125729 i|z|zn$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5334 \$125731 i|z$16 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5340 VSS|anode|cathode|clk|vss \$125731 z$15 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5356 \$125732 i|zn$8 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5357 VSS|anode|cathode|clk|vss \$125733 \$125734 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5358 VSS|anode|cathode|clk|vss \$125732 \$125733 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5359 VSS|anode|cathode|clk|vss \$125734 i|z$12 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5360 i|zn$1 i|z|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5368 \$125737 i|z$15 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5369 VSS|anode|cathode|clk|vss \$125738 \$125739 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5370 VSS|anode|cathode|clk|vss \$125737 \$125738 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5371 VSS|anode|cathode|clk|vss \$125739 i|z$13 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5372 \$125741 RESULT[1]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p
+ AD=1.65025p PS=9.3u PD=9.48u
M$5378 VSS|anode|cathode|clk|vss \$125741 i|z|zn$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5394 \$125743 i|z|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5395 VSS|anode|cathode|clk|vss \$125744 \$125745 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5396 VSS|anode|cathode|clk|vss \$125743 \$125744 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5397 VSS|anode|cathode|clk|vss \$125745 i|z$81 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5398 \$125747 \$125626 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5399 VSS|anode|cathode|clk|vss cp|z$2 \$125626 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5400 a1|b|i|q$3 \$126468 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$5401 VSS|anode|cathode|clk|vss \$127549 i|z$75 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5403 VSS|anode|cathode|clk|vss i|z \$127549 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5404 i|z|zn$1 i|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5412 VSS|anode|cathode|clk|vss i|z$67 \$127371 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5418 VSS|anode|cathode|clk|vss \$127371 z$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5434 \$127372 i|z$17 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5435 VSS|anode|cathode|clk|vss \$127110 \$127373 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5436 \$127110 \$127372 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5437 VSS|anode|cathode|clk|vss \$127373 i|z$19 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5438 VSS|anode|cathode|clk|vss \$127550 i|z$20 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5440 VSS|anode|cathode|clk|vss i|z$26 \$127550 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5441 VSS|anode|cathode|clk|vss \$127552 i|z$21 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5443 VSS|anode|cathode|clk|vss i|z$27 \$127552 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5444 VSS|anode|cathode|clk|vss i|z$22 \$127378 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5450 VSS|anode|cathode|clk|vss \$127378 z$12 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5466 VSS|anode|cathode|clk|vss RESULT[4]|c2p|core|i|q \$127379
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p
+ AD=1.730525p PS=9.48u PD=9.3u
M$5472 VSS|anode|cathode|clk|vss \$127379 i|z|zn$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5488 VSS|anode|cathode|clk|vss i|z$23 \$127382 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5494 VSS|anode|cathode|clk|vss \$127382 a1|i|z|zn VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5510 \$127384 i|z$18 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5511 VSS|anode|cathode|clk|vss \$127112 \$127385 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5512 \$127112 \$127384 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5513 VSS|anode|cathode|clk|vss \$127385 i|z$31 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5514 i|zn$3 i|z|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5522 VSS|anode|cathode|clk|vss RESULT[2]|c2p|core|i|q \$127387
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p
+ AD=1.730525p PS=9.48u PD=9.3u
M$5528 VSS|anode|cathode|clk|vss \$127387 i|z|zn$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5544 VSS|anode|cathode|clk|vss i|z$36 \$127389 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5550 VSS|anode|cathode|clk|vss \$127389 z$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5566 VSS|anode|cathode|clk|vss \$127554 i|z$106 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5568 VSS|anode|cathode|clk|vss i|z$28 \$127554 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5569 VSS|anode|cathode|clk|vss \$127556 i|z$24 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5571 VSS|anode|cathode|clk|vss i|z$12 \$127556 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5572 VSS|anode|cathode|clk|vss \$127557 i|z$15 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5574 VSS|anode|cathode|clk|vss i|z$29 \$127557 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5575 i|z|zn$6 i|zn$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5583 \$127392 i|zn$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5584 VSS|anode|cathode|clk|vss \$127114 \$127393 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5585 \$127114 \$127392 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5586 VSS|anode|cathode|clk|vss \$127393 i|z$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5587 i|z|zn$3 i|zn$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5595 \$127394 i|z$30 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$5596 VSS|anode|cathode|clk|vss \$127394 i|z$25 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$5597 \$127396 CLK|core|i|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p
+ PS=1.85u PD=1.55u
M$5598 VSS|anode|cathode|clk|vss \$127396 i|z$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$5599 VSS|anode|cathode|clk|vss \$125626 \$127014 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$5600 \$127014 d|zn$8 \$125627 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$5601 \$125627 \$125747 \$127016 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$5602 VSS|anode|cathode|clk|vss \$125748 \$127016 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$5603 VSS|anode|cathode|clk|vss \$125627 \$125748 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$5604 \$125748 \$125747 \$126892 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$5605 \$126892 \$125626 \$126997 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$5606 VSS|anode|cathode|clk|vss \$126468 \$126997 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$5607 VSS|anode|cathode|clk|vss \$126892 \$126468 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$5608 i|zn$4 i|z|zn$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5616 i|zn$5 i|z|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5624 VSS|anode|cathode|clk|vss a2|z$5 \$130091 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5625 \$130091 a1|z$12 \$128987 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5626 \$128987 a1|z$12 \$130090 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5627 \$130090 a2|z$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5628 VSS|anode|cathode|clk|vss \$128987 i|z$6 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5632 \$128988 i|z$38 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5633 VSS|anode|cathode|clk|vss \$128989 \$128990 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5634 VSS|anode|cathode|clk|vss \$128988 \$128989 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5635 VSS|anode|cathode|clk|vss \$128990 i|z$27 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5636 VSS|anode|cathode|clk|vss \$129730 i|z$32 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5638 VSS|anode|cathode|clk|vss i|z$42 \$129730 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5639 VSS|anode|cathode|clk|vss i|z$43 \$128992 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5641 VSS|anode|cathode|clk|vss \$128992 a2|z$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5645 \$128994 i|z|zn$8 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5646 VSS|anode|cathode|clk|vss \$128995 \$128996 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5647 VSS|anode|cathode|clk|vss \$128994 \$128995 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5648 VSS|anode|cathode|clk|vss \$128996 i|z$33 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5649 \$128998 i|z$39 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5650 VSS|anode|cathode|clk|vss \$128999 \$129000 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5651 VSS|anode|cathode|clk|vss \$128998 \$128999 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5652 VSS|anode|cathode|clk|vss \$129000 i|z$34 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5653 VSS|anode|cathode|clk|vss \$129733 i|z$35 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5655 VSS|anode|cathode|clk|vss i|z$44 \$129733 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5656 \$129003 i|z$45 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5662 VSS|anode|cathode|clk|vss \$129003 z$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5678 \$129004 i|z$46 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5684 VSS|anode|cathode|clk|vss \$129004 z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5700 \$129005 i|z|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.925u AS=0.942125p AD=0.834125p PS=5.67u PD=4.65u
M$5703 VSS|anode|cathode|clk|vss \$129005 i|z$36 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.3904p AD=2.4984p PS=12.4u PD=13.42u
M$5711 \$129007 i|z$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5717 VSS|anode|cathode|clk|vss \$129007 a1|z$11 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5733 \$129009 i|z$48 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5739 VSS|anode|cathode|clk|vss \$129009 z$13 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5755 \$129010 i|z$24 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5756 VSS|anode|cathode|clk|vss \$129011 \$129012 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5757 VSS|anode|cathode|clk|vss \$129010 \$129011 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5758 VSS|anode|cathode|clk|vss \$129012 i|z$29 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5759 i|z|zn$2 i|zn$8 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5767 \$129013 i|z$49 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5773 VSS|anode|cathode|clk|vss \$129013 z$14 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5789 \$129014 a2|i|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5790 VSS|anode|cathode|clk|vss \$129015 \$129016 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5791 VSS|anode|cathode|clk|vss \$129014 \$129015 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5792 VSS|anode|cathode|clk|vss \$129016 i|z$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5793 \$129017 i|z$113 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5794 VSS|anode|cathode|clk|vss \$129018 \$129019 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5795 VSS|anode|cathode|clk|vss \$129017 \$129018 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5796 VSS|anode|cathode|clk|vss \$129019 i|z$28 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5797 \$129970 \$129970 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$5798 i|zn$6 i|z|zn$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5806 i|z|zn$5 i|zn$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5814 i|zn$7 i|zn$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5822 \$129022 i|z$60 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5823 VSS|anode|cathode|clk|vss \$129023 \$129024 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5824 VSS|anode|cathode|clk|vss \$129022 \$129023 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5825 VSS|anode|cathode|clk|vss \$129024 i|z$37 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5826 VSS|anode|cathode|clk|vss \$129740 i|z$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5828 VSS|anode|cathode|clk|vss i|z$13 \$129740 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5829 \$129026 RESULT[3]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p
+ AD=1.65025p PS=9.3u PD=9.48u
M$5835 VSS|anode|cathode|clk|vss \$129026 i|z|zn$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5851 a2|zn a1|i|q$1 \$130187 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5852 \$130187 a1|a2|a3|z \$130188 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5853 \$130188 a2|a3|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5854 VSS|anode|cathode|clk|vss cp|i|z \$128890 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2511p AD=0.2034p PS=1.55u PD=1.85u
M$5855 VSS|anode|cathode|clk|vss \$128890 cp|z$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$5856 a2 z$7 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5857 a2$1 z$4 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.16u
+ AS=1.2204p AD=1.2204p PS=11.1u PD=11.1u
M$5858 a2$1 z$7 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5868 a1|c|i|zn a2$1 \$130271 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5872 a1|c|i|zn a1|z$11 \$130271 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5876 \$130333 a2|b|z \$130271 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5880 \$130333 a1|c|i|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5884 a1|c|i|zn a2$1 \$130272 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5888 a1|c|i|zn a1|z$11 \$130272 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5892 \$130334 a2|b|z \$130272 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5896 \$130334 a1|c|i|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5900 a1|c|i|zn a2$1 \$130273 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5904 a1|c|i|zn a1|z$11 \$130273 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5908 \$130335 a2|b|z \$130273 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5912 \$130335 a1|c|i|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5916 a1|c|i|zn a2$1 \$130274 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5920 a1|c|i|zn a1|z$11 \$130274 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5924 \$130336 a2|b|z \$130274 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5928 \$130336 a1|c|i|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5932 VSS|anode|cathode|clk|vss a2|b|z \$130598 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5933 \$130598 a1|c|i|zn a1|c|i|zn$1 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5934 a1|c|i|zn$1 a1|c|i|zn \$130599 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5935 \$130599 a2|b|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5936 \$130275 a1|c|i|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.154925p AD=0.1105875p PS=1.73u PD=1.13u
M$5937 VSS|anode|cathode|clk|vss \$130275 i|z$53 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1105875p AD=0.15625p PS=1.13u PD=1.73u
M$5938 VSS|anode|cathode|clk|vss \$130779 z$22 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5940 VSS|anode|cathode|clk|vss i|z$53 \$130779 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5941 \$130338 i|z$32 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5942 VSS|anode|cathode|clk|vss \$130277 \$130339 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5943 \$130277 \$130338 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5944 VSS|anode|cathode|clk|vss \$130339 i|z$26 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5945 VSS|anode|cathode|clk|vss i|z$40 \$130340 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5951 VSS|anode|cathode|clk|vss \$130340 z$23 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5967 \$130342 i|zn$11 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5968 VSS|anode|cathode|clk|vss \$130278 \$130343 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5969 \$130278 \$130342 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5970 VSS|anode|cathode|clk|vss \$130343 i|z$56 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5971 i|zn$8 i|z|zn$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5979 VSS|anode|cathode|clk|vss i|z$47 \$130346 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5985 VSS|anode|cathode|clk|vss \$130346 z$16 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6001 \$130347 i|z$52 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6002 VSS|anode|cathode|clk|vss \$130279 \$130348 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6003 \$130279 \$130347 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6004 VSS|anode|cathode|clk|vss \$130348 i|z$57 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6005 VSS|anode|cathode|clk|vss i|z$36 \$130350 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6011 VSS|anode|cathode|clk|vss \$130350 z$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6027 \$130351 i|z$35 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6028 VSS|anode|cathode|clk|vss \$130280 \$130352 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6029 \$130280 \$130351 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6030 VSS|anode|cathode|clk|vss \$130352 i|z$51 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6031 \$130353 i|z$54 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6032 VSS|anode|cathode|clk|vss \$130282 \$130354 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6033 \$130282 \$130353 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6034 VSS|anode|cathode|clk|vss \$130354 i|z$58 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6035 VSS|anode|cathode|clk|vss VALID|a3|c2p|core|i|z i|zn$9
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.88u AS=1.3032p AD=1.3032p
+ PS=7.22u PD=7.22u
M$6039 VSS|anode|cathode|clk|vss a2|i|z i|zn$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.3032p AD=1.3032p PS=7.22u PD=7.22u
M$6043 VSS|anode|cathode|clk|vss SAMPLE|a1|c2p|core|i|z i|zn$9
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.88u AS=1.3032p AD=1.3032p
+ PS=7.22u PD=7.22u
M$6047 a1|i|z|zn i|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=4.32u AS=1.9008p AD=1.9008p PS=10.32u PD=10.32u
M$6053 \$130283 \$130283 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6054 i|zn$10 i|z|zn$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6062 \$130358 i|z|zn$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6063 VSS|anode|cathode|clk|vss \$130284 \$130359 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6064 \$130284 \$130358 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6065 VSS|anode|cathode|clk|vss \$130359 i|z$42 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6066 VSS|anode|cathode|clk|vss \$130780 i|z$59 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6068 VSS|anode|cathode|clk|vss i|z$34 \$130780 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6069 VSS|anode|cathode|clk|vss \$130781 i|z$60 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6071 VSS|anode|cathode|clk|vss i|z$1 \$130781 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6072 VSS|anode|cathode|clk|vss \$130782 i|z$49 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6074 VSS|anode|cathode|clk|vss i|z$58 \$130782 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6075 \$130362 i|z|zn$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6076 VSS|anode|cathode|clk|vss \$130285 \$130363 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6077 \$130285 \$130362 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6078 VSS|anode|cathode|clk|vss \$130363 i|z$114 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6079 \$130364 i|z$55 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6080 VSS|anode|cathode|clk|vss \$130287 \$130365 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6081 \$130287 \$130364 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6082 VSS|anode|cathode|clk|vss \$130365 i|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6083 zn$5 \$130824 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6084 \$130366 i|z$41 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6085 VSS|anode|cathode|clk|vss \$130288 \$130367 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6086 \$130288 \$130366 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6087 VSS|anode|cathode|clk|vss \$130367 i|z$61 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6088 VSS|anode|cathode|clk|vss i|zn$9 \$130369 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.925u AS=0.942125p AD=0.834125p PS=5.67u PD=4.65u
M$6091 VSS|anode|cathode|clk|vss \$130369 i|z$23 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.3904p AD=2.4984p PS=12.4u PD=13.42u
M$6099 VSS|anode|cathode|clk|vss \$130783 i|z$55 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6101 VSS|anode|cathode|clk|vss i|z$37 \$130783 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6102 i|zn$2 SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p
+ PS=13.42u PD=13.42u
M$6110 VSS|anode|cathode|clk|vss i|z$11 \$130370 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6112 VSS|anode|cathode|clk|vss \$130370 i|z$18 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6116 VSS|anode|cathode|clk|vss i|z$25 \$130371 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6122 VSS|anode|cathode|clk|vss \$130371 a2|i|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6138 \$130289 CLK|core|i|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p
+ PS=1.85u PD=1.55u
M$6139 VSS|anode|cathode|clk|vss \$130289 i|z$62 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$6140 \$130290 i|z$62 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$6141 VSS|anode|cathode|clk|vss \$130290 i|z$30 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$6142 a2|z$1 \$130373 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6143 VSS|anode|cathode|clk|vss b|q \$130373 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6144 \$130373 a1|b|i|q$2 \$130753 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6145 \$130753 a2|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6146 \$130374 \$130291 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6147 VSS|anode|cathode|clk|vss cp|z$2 \$130291 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6148 \$130292 \$130374 \$130747 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$6149 \$130747 \$130293 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$6150 \$130294 \$130291 \$130749 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$6151 \$130749 \$130375 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$6152 \$130293 \$130374 \$130294 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$6153 VSS|anode|cathode|clk|vss \$130291 \$130744 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$6154 \$130744 d|zn$3 \$130292 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$6155 VSS|anode|cathode|clk|vss \$130292 \$130293 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$6156 VSS|anode|cathode|clk|vss \$130294 \$130375 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$6157 RESULT[2]|c2p|core|i|q \$130375 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$6158 a1|c|i|zn$1 a2 \$132940 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6162 a1|c|i|zn$1 a1|z$11 \$132940 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6166 \$132709 a2|b|z \$132940 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6170 \$132709 a1|c|i|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6174 a1|c|i|zn$1 a2 \$132941 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6178 a1|c|i|zn$1 a1|z$11 \$132941 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6182 \$132710 a2|b|z \$132941 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6186 \$132710 a1|c|i|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6190 a1|c|i|zn$1 a2 \$132942 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6194 a1|c|i|zn$1 a1|z$11 \$132942 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6198 \$132711 a2|b|z \$132942 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6202 \$132711 a1|c|i|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6206 a1|c|i|zn$1 a2 \$132943 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6210 a1|c|i|zn$1 a1|z$11 \$132943 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6214 \$132712 a2|b|z \$132943 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6218 \$132712 a1|c|i|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6222 VSS|anode|cathode|clk|vss a2|b|z \$133171 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6223 \$133171 a1|c|i|zn$1 a1|c|i|zn VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6224 a1|c|i|zn a1|c|i|zn$1 \$133169 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6225 \$133169 a2|b|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6226 VSS|anode|cathode|clk|vss \$132660 a2|a3|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6228 VSS|anode|cathode|clk|vss i|z$65 \$132660 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6229 VSS|anode|cathode|clk|vss a2|z$4 \$133174 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6230 \$133174 a1|i|z|zn \$131972 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6231 \$131972 a1|i|z|zn \$133172 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6232 \$133172 a2|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6233 VSS|anode|cathode|clk|vss \$131972 i|z$66 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6237 \$131974 i|z$74 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6243 VSS|anode|cathode|clk|vss \$131974 z$11 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6259 \$132944 \$132944 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6260 i|z|zn$7 i|zn$10 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6268 \$131975 i|z$75 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6274 VSS|anode|cathode|clk|vss \$131975 z$25 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6290 \$131977 i|z|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.925u AS=0.942125p AD=0.834125p PS=5.67u PD=4.65u
M$6293 VSS|anode|cathode|clk|vss \$131977 i|z$67 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.3904p AD=2.4984p PS=12.4u PD=13.42u
M$6301 \$131979 i|z|zn$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6302 VSS|anode|cathode|clk|vss \$131980 \$131981 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6303 VSS|anode|cathode|clk|vss \$131979 \$131980 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6304 VSS|anode|cathode|clk|vss \$131981 i|z$63 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6305 \$131982 i|z$76 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6311 VSS|anode|cathode|clk|vss \$131982 z$10 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6327 \$131983 i|z$59 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6333 VSS|anode|cathode|clk|vss \$131983 z$19 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6349 VSS|anode|cathode|clk|vss \$132664 i|z$74 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6351 VSS|anode|cathode|clk|vss i|z$101 \$132664 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6352 \$131984 i|zn$10 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6353 VSS|anode|cathode|clk|vss \$131985 \$131986 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6354 VSS|anode|cathode|clk|vss \$131984 \$131985 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6355 VSS|anode|cathode|clk|vss \$131986 i|z$68 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6356 i|zn$11 i|z|zn$8 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6364 \$132946 \$132946 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6365 \$131989 b|i|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6371 VSS|anode|cathode|clk|vss \$131989 i|z|zn$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6387 VSS|anode|cathode|clk|vss \$132668 i|z$69 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6389 VSS|anode|cathode|clk|vss i|z$77 \$132668 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6390 \$131991 i|z$72 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6391 VSS|anode|cathode|clk|vss \$131992 \$131993 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6392 VSS|anode|cathode|clk|vss \$131991 \$131992 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6393 VSS|anode|cathode|clk|vss \$131993 i|z$64 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6394 \$131994 i|z$69 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6395 VSS|anode|cathode|clk|vss \$131995 \$131996 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6396 VSS|anode|cathode|clk|vss \$131994 \$131995 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6397 VSS|anode|cathode|clk|vss \$131996 i|z$70 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6398 VSS|anode|cathode|clk|vss \$132670 i|z$46 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6400 VSS|anode|cathode|clk|vss i|z$79 \$132670 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6401 \$131998 i|z$103 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6402 VSS|anode|cathode|clk|vss \$131999 \$132000 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6403 VSS|anode|cathode|clk|vss \$131998 \$131999 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6404 VSS|anode|cathode|clk|vss \$132000 i|z$111 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6405 \$132001 i|z$73 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6406 VSS|anode|cathode|clk|vss \$132002 \$132003 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6407 VSS|anode|cathode|clk|vss \$132001 \$132002 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6408 VSS|anode|cathode|clk|vss \$132003 i|z$71 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6409 VSS|anode|cathode|clk|vss \$132671 i|z$16 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6411 VSS|anode|cathode|clk|vss i|z$80 \$132671 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6412 \$132005 b|i|q$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6418 VSS|anode|cathode|clk|vss \$132005 i|z|zn$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6434 \$132007 \$131965 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6435 VSS|anode|cathode|clk|vss cp|z$1 \$131965 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6436 a1|i|q$1 \$132009 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6437 \$133281 \$133281 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6438 zn$3 \$133696 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6439 i|z|zn i|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6447 VSS|anode|cathode|clk|vss i|z$66 \$133345 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6453 VSS|anode|cathode|clk|vss \$133345 a2|b|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6469 zn \$133697 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6470 \$133346 i|z$83 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6471 VSS|anode|cathode|clk|vss \$133283 \$133347 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6472 \$133283 \$133346 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6473 VSS|anode|cathode|clk|vss \$133347 i|z$86 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6474 VSS|anode|cathode|clk|vss i|zn$7 \$133349 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.925u AS=0.942125p AD=0.834125p PS=5.67u PD=4.65u
M$6477 VSS|anode|cathode|clk|vss \$133349 a1|z$12 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.3904p AD=2.4984p PS=12.4u PD=13.42u
M$6485 VSS|anode|cathode|clk|vss \$133351 i|z$83 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6487 VSS|anode|cathode|clk|vss i|z$87 \$133351 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6488 VSS|anode|cathode|clk|vss \$133353 i|z$88 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6490 VSS|anode|cathode|clk|vss i|z$102 \$133353 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6491 \$133355 a1|i|z|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6492 VSS|anode|cathode|clk|vss \$133284 \$133356 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6493 \$133284 \$133355 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6494 VSS|anode|cathode|clk|vss \$133356 i|z$43 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6495 \$131962 a1|c|i|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.154925p AD=0.1105875p PS=1.73u PD=1.13u
M$6496 VSS|anode|cathode|clk|vss \$131962 i|z$65 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1105875p AD=0.15625p PS=1.13u PD=1.73u
M$6497 VSS|anode|cathode|clk|vss i|z$89 \$133358 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6503 VSS|anode|cathode|clk|vss \$133358 z$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6519 \$133359 i|z$84 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6520 VSS|anode|cathode|clk|vss \$133286 \$133360 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6521 \$133286 \$133359 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6522 VSS|anode|cathode|clk|vss \$133360 i|z$80 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6523 \$133361 i|zn$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6524 VSS|anode|cathode|clk|vss \$133287 \$133362 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6525 \$133287 \$133361 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6526 VSS|anode|cathode|clk|vss \$133362 i|z$90 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6527 VSS|anode|cathode|clk|vss \$133364 i|z$82 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6529 VSS|anode|cathode|clk|vss i|z$91 \$133364 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6530 i|zn$12 i|z|zn$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6538 VSS|anode|cathode|clk|vss i|z$31 \$133367 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6540 VSS|anode|cathode|clk|vss \$133367 a2|z$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6544 i|zn a1|i|z|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=4.32u AS=1.9008p AD=1.9008p PS=10.32u PD=10.32u
M$6550 VSS|anode|cathode|clk|vss \$133368 i|z$17 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6552 VSS|anode|cathode|clk|vss i|z$81 \$133368 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6553 \$133369 i|z$50 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6554 VSS|anode|cathode|clk|vss \$133288 \$133370 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6555 \$133288 \$133369 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6556 VSS|anode|cathode|clk|vss \$133370 i|z$79 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6557 VSS|anode|cathode|clk|vss i|z$88 \$133371 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6563 VSS|anode|cathode|clk|vss \$133371 z$18 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6579 VSS|anode|cathode|clk|vss \$133372 i|z$39 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6581 VSS|anode|cathode|clk|vss i|z$19 \$133372 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6582 VSS|anode|cathode|clk|vss \$133373 i|z$41 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6584 VSS|anode|cathode|clk|vss i|z$33 \$133373 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6585 VSS|anode|cathode|clk|vss i|z$78 \$133374 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6591 VSS|anode|cathode|clk|vss \$133374 z$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6607 VSS|anode|cathode|clk|vss \$133376 i|z$45 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6609 VSS|anode|cathode|clk|vss i|z$93 \$133376 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6610 VSS|anode|cathode|clk|vss \$133378 i|z$94 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6612 VSS|anode|cathode|clk|vss i|z$95 \$133378 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6613 VSS|anode|cathode|clk|vss \$133381 i|z$89 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6615 VSS|anode|cathode|clk|vss i|z$92 \$133381 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6616 VSS|anode|cathode|clk|vss b|i|q$2 \$133383 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6622 VSS|anode|cathode|clk|vss \$133383 i|z|zn$6 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6638 \$133384 i|z|zn$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6639 VSS|anode|cathode|clk|vss \$133289 \$133385 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6640 \$133289 \$133384 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6641 VSS|anode|cathode|clk|vss \$133385 i|z$91 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6642 \$133386 i|z$85 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6643 VSS|anode|cathode|clk|vss \$133291 \$133387 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6644 \$133291 \$133386 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6645 VSS|anode|cathode|clk|vss \$133387 i|z$96 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6646 VSS|anode|cathode|clk|vss \$133389 i|z$47 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6648 VSS|anode|cathode|clk|vss i|z$70 \$133389 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6649 \$133390 i|z$82 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6650 VSS|anode|cathode|clk|vss \$133292 \$133391 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6651 \$133292 \$133390 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6652 VSS|anode|cathode|clk|vss \$133391 i|z$97 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6653 VSS|anode|cathode|clk|vss \$133393 i|z$85 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6655 VSS|anode|cathode|clk|vss i|z$71 \$133393 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6656 i|z|zn$9 i|zn$13 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6664 \$133395 i|z$107 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6665 VSS|anode|cathode|clk|vss \$133293 \$133396 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6666 \$133293 \$133395 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6667 VSS|anode|cathode|clk|vss \$133396 i|z$100 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6668 \$133397 i|zn$12 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6669 VSS|anode|cathode|clk|vss \$133294 \$133398 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6670 \$133294 \$133397 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6671 VSS|anode|cathode|clk|vss \$133398 i|z$98 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6672 VSS|anode|cathode|clk|vss \$133401 i|z$52 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6674 VSS|anode|cathode|clk|vss i|z$99 \$133401 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6675 VSS|anode|cathode|clk|vss \$133402 i|z$72 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6677 VSS|anode|cathode|clk|vss i|z$98 \$133402 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6678 VSS|anode|cathode|clk|vss \$131965 \$133229 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$6679 \$133229 d|zn$4 \$131966 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$6680 \$131966 \$132007 \$133230 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$6681 VSS|anode|cathode|clk|vss \$132008 \$133230 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$6682 VSS|anode|cathode|clk|vss \$131966 \$132008 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$6683 \$132008 \$132007 \$132948 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$6684 \$132948 \$131965 \$133220 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$6685 VSS|anode|cathode|clk|vss \$132009 \$133220 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$6686 VSS|anode|cathode|clk|vss \$132948 \$132009 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$6687 \$133304 a2|a3|zn b|zn$4 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6688 b|zn$4 RST|a1|b|cdn|core|i|p2c \$133304 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6689 \$133304 a1|b|i|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6690 \$133305 i|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$6691 VSS|anode|cathode|clk|vss \$133305 cp|i|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$6692 \$134936 i|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6698 VSS|anode|cathode|clk|vss \$134936 z$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6714 \$134937 i|z$9 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6715 VSS|anode|cathode|clk|vss \$134938 \$134875 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6716 VSS|anode|cathode|clk|vss \$134937 \$134938 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6717 VSS|anode|cathode|clk|vss \$134875 i|z$87 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6718 VSS|anode|cathode|clk|vss \$135839 i|z$50 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6720 VSS|anode|cathode|clk|vss i|z$57 \$135839 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6721 zn$4 \$134939 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6722 \$134940 i|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6728 VSS|anode|cathode|clk|vss \$134940 z$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6744 VSS|anode|cathode|clk|vss \$135840 i|z$22 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6746 VSS|anode|cathode|clk|vss i|z$86 \$135840 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6747 \$134941 i|z|zn$9 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6748 VSS|anode|cathode|clk|vss \$134942 \$134876 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6749 VSS|anode|cathode|clk|vss \$134941 \$134942 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6750 VSS|anode|cathode|clk|vss \$134876 i|z$99 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6751 \$134943 b|i|q$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6757 VSS|anode|cathode|clk|vss \$134943 i|z|zn$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6773 \$134944 i|z$20 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6774 VSS|anode|cathode|clk|vss \$134945 \$134877 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6775 VSS|anode|cathode|clk|vss \$134944 \$134945 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6776 VSS|anode|cathode|clk|vss \$134877 i|z$105 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6777 \$134947 i|z$106 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6778 VSS|anode|cathode|clk|vss \$134949 \$134878 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6779 VSS|anode|cathode|clk|vss \$134947 \$134949 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6780 VSS|anode|cathode|clk|vss \$134878 i|z$101 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6781 VSS|anode|cathode|clk|vss \$135841 i|z$103 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6783 VSS|anode|cathode|clk|vss i|z$56 \$135841 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6784 \$136067 \$136067 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6785 VSS|anode|cathode|clk|vss \$135842 i|z$38 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6787 VSS|anode|cathode|clk|vss i|z$90 \$135842 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6788 i|zn$13 i|z|zn$9 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6796 VSS|anode|cathode|clk|vss \$135843 i|z$107 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6798 VSS|anode|cathode|clk|vss i|z$97 \$135843 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6799 zn$2 \$134951 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6800 \$134952 i|z$108 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6801 VSS|anode|cathode|clk|vss \$134954 \$134879 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6802 VSS|anode|cathode|clk|vss \$134952 \$134954 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6803 VSS|anode|cathode|clk|vss \$134879 i|z$92 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6804 \$134955 i|z$109 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6805 VSS|anode|cathode|clk|vss \$134957 \$134880 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6806 VSS|anode|cathode|clk|vss \$134955 \$134957 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6807 VSS|anode|cathode|clk|vss \$134880 i|z$77 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6808 i|z|zn$4 i|zn$12 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6816 VSS|anode|cathode|clk|vss \$135844 i|z$110 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6818 VSS|anode|cathode|clk|vss i|z$104 \$135844 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6819 i|z|zn$8 i|zn$11 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6827 VSS|anode|cathode|clk|vss \$135845 i|z$73 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6829 VSS|anode|cathode|clk|vss i|z$68 \$135845 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6830 VSS|anode|cathode|clk|vss \$135846 i|z$108 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6832 VSS|anode|cathode|clk|vss i|z$64 \$135846 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6833 \$134959 i|z$110 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6834 VSS|anode|cathode|clk|vss \$134960 \$134881 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6835 VSS|anode|cathode|clk|vss \$134959 \$134960 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6836 VSS|anode|cathode|clk|vss \$134881 i|z$95 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6837 \$134961 i|z$94 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6838 VSS|anode|cathode|clk|vss \$134962 \$134882 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6839 VSS|anode|cathode|clk|vss \$134961 \$134962 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6840 VSS|anode|cathode|clk|vss \$134882 i|z$93 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6841 VSS|anode|cathode|clk|vss \$135847 i|z$84 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6843 VSS|anode|cathode|clk|vss i|z$61 \$135847 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6844 VSS|anode|cathode|clk|vss \$135848 i|z$40 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6846 VSS|anode|cathode|clk|vss i|z$105 \$135848 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6847 VSS|anode|cathode|clk|vss \$135849 i|z$76 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6849 VSS|anode|cathode|clk|vss i|z$96 \$135849 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6850 \$134963 i|z$21 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6851 VSS|anode|cathode|clk|vss \$134964 \$134883 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6852 VSS|anode|cathode|clk|vss \$134963 \$134964 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6853 VSS|anode|cathode|clk|vss \$134883 i|z$102 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6854 \$134965 i|z$112 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6855 VSS|anode|cathode|clk|vss \$134966 \$134884 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6856 VSS|anode|cathode|clk|vss \$134965 \$134966 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6857 VSS|anode|cathode|clk|vss \$134884 i|z$44 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6858 VSS|anode|cathode|clk|vss \$135850 i|z$48 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6860 VSS|anode|cathode|clk|vss i|z$100 \$135850 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6861 \$134967 i|zn$13 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6862 VSS|anode|cathode|clk|vss \$134968 \$134885 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6863 VSS|anode|cathode|clk|vss \$134967 \$134968 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6864 VSS|anode|cathode|clk|vss \$134885 i|z$104 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6865 VSS|anode|cathode|clk|vss \$135851 i|z$78 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6867 VSS|anode|cathode|clk|vss i|z$51 \$135851 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6868 \$134969 \$134735 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6869 VSS|anode|cathode|clk|vss cp|z$2 \$134735 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6870 a1|b|i|q$2 \$134970 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6871 VSS|anode|cathode|clk|vss a2|zn$6 \$136317 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6872 \$136317 a1|z$13 d|zn$2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6873 d|zn$2 b|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6874 zn$1 \$137099 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6875 \$136386 i|zn$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6876 VSS|anode|cathode|clk|vss \$136342 \$136387 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6877 \$136342 \$136386 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6878 VSS|anode|cathode|clk|vss \$136387 i|z$14 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6879 VSS|anode|cathode|clk|vss i|zn$5 \$136388 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6885 VSS|anode|cathode|clk|vss \$136388 z$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6901 VSS|anode|cathode|clk|vss i|z$67 \$136389 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6907 VSS|anode|cathode|clk|vss \$136389 z$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6923 VSS|anode|cathode|clk|vss \$136706 i|z$113 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6925 VSS|anode|cathode|clk|vss i|z$114 \$136706 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6926 VSS|anode|cathode|clk|vss \$136708 i|z$54 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6928 VSS|anode|cathode|clk|vss i|z$111 \$136708 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6929 VSS|anode|cathode|clk|vss \$136709 i|z$112 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6931 VSS|anode|cathode|clk|vss i|z$63 \$136709 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6932 \$136391 \$136343 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6933 VSS|anode|cathode|clk|vss cp|i|z \$136343 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6934 \$136344 \$136391 \$136685 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$6935 \$136685 \$136392 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$6936 \$136345 \$136343 \$136680 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$6937 \$136680 \$136393 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$6938 \$136392 \$136391 \$136345 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$6939 VSS|anode|cathode|clk|vss \$136343 \$136683 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$6940 \$136683 d|zn$9 \$136344 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$6941 VSS|anode|cathode|clk|vss \$136344 \$136392 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$6942 VSS|anode|cathode|clk|vss \$136345 \$136393 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$6943 VSS|anode|cathode|clk|vss \$134735 \$136321 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$6944 \$136321 d|zn$6 \$134736 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$6945 \$134736 \$134969 \$136323 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$6946 VSS|anode|cathode|clk|vss \$134886 \$136323 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$6947 VSS|anode|cathode|clk|vss \$134736 \$134886 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$6948 \$134886 \$134969 \$136070 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$6949 \$136070 \$134735 \$136311 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$6950 VSS|anode|cathode|clk|vss \$134970 \$136311 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$6951 VSS|anode|cathode|clk|vss \$136070 \$134970 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$6952 a1|b|i|q$1 \$136393 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6953 \$136394 \$136346 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6954 VSS|anode|cathode|clk|vss cp|z$3 \$136346 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6955 \$136347 \$136394 \$136676 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$6956 \$136676 \$136395 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$6957 \$136348 \$136346 \$136678 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$6958 \$136678 \$136396 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$6959 \$136395 \$136394 \$136348 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$6960 VSS|anode|cathode|clk|vss \$136346 \$136674 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$6961 \$136674 d|zn$10 \$136347 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$6962 VSS|anode|cathode|clk|vss \$136347 \$136395 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$6963 VSS|anode|cathode|clk|vss \$136348 \$136396 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$6964 a1|b|i|q \$136396 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6965 \$139964 \$140018 \$139964 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7001 \$139965 \$140019 \$139965 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7037 \$139966 \$140020 \$139966 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7073 \$139967 \$140021 \$139967 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7109 \$139968 \$140022 \$139968 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7145 \$139969 \$140023 \$139969 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7181 \$139970 \$140024 \$139970 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7217 \$139971 \$140025 \$139971 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7253 \$139972 \$140026 \$139972 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7289 \$139973 \$140027 \$139973 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7325 \$140028 a1|z$3 \$140390 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$7326 \$140390 a2|z$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.655u AS=0.271825p AD=0.2901875p PS=1.485u PD=1.55u
M$7327 VSS|anode|cathode|clk|vss \$140028 d|z$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2901875p AD=0.4068p PS=1.55u PD=2.57u
M$7328 a2|zn$6 a1|b|i|q$2 \$139778 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$7329 \$139778 a1|a2|a3|z \$139781 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$7330 \$139781 a2|a3|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$7691 \$141594 \$141285 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$7692 VSS|anode|cathode|clk|vss cp|z$3 \$141285 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$7693 a2|i|q \$141596 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$7694 a2|z \$141598 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$7695 VSS|anode|cathode|clk|vss b|i|q \$141598 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$7696 \$141598 a1|b|i|q \$142915 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$7697 \$142915 a2|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$7698 \$145293 \$145605 \$145293 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7710 \$143069 z$26 \$143069 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7711 \$140018 zn$3 \$143069 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7712 \$140018 z$26 \$140018 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7727 \$143070 zn$3 \$140018 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7728 \$143070 z$26 \$143070 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7743 \$143071 zn$3 \$140018 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7744 \$143071 z$26 \$143071 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7746 \$145294 \$145606 \$145294 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=829.44u AS=354.5856p AD=354.5856p PS=1883.52u PD=1883.52u
M$7758 \$143072 z$26 \$143072 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7759 \$140019 zn$3 \$143072 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7760 \$140019 z$26 \$140019 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7775 \$143073 zn$3 \$140019 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7776 \$143073 z$26 \$143073 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7791 \$143074 zn$3 \$140019 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7792 \$143074 z$26 \$143074 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7794 \$145295 \$145607 \$145295 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=414.72u AS=177.2928p AD=177.2928p PS=941.76u PD=941.76u
M$7806 \$143075 z$26 \$143075 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7807 \$140020 zn$3 \$143075 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7808 \$140020 z$26 \$140020 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7823 \$143076 zn$3 \$140020 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7824 \$143076 z$26 \$143076 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7839 \$143077 zn$3 \$140020 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7840 \$143077 z$26 \$143077 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7842 \$145296 \$145608 \$145296 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=103.68u AS=44.3232p AD=44.3232p PS=235.44u PD=235.44u
M$7854 \$143078 z$26 \$143078 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7855 \$140021 zn$3 \$143078 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7856 \$140021 z$26 \$140021 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7871 \$143079 zn$3 \$140021 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7872 \$143079 z$26 \$143079 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7887 \$143080 zn$3 \$140021 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7888 \$143080 z$26 \$143080 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7890 \$145297 \$145609 \$145297 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7902 \$143081 z$26 \$143081 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7903 \$140022 zn$3 \$143081 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7904 \$140022 z$26 \$140022 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7919 \$143082 zn$3 \$140022 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7920 \$143082 z$26 \$143082 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7935 \$143083 zn$3 \$140022 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7936 \$143083 z$26 \$143083 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7938 \$145298 \$145610 \$145298 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7950 \$143084 z$26 \$143084 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7951 \$140023 zn$3 \$143084 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7952 \$140023 z$26 \$140023 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7967 \$143085 zn$3 \$140023 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7968 \$143085 z$26 \$143085 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7983 \$143086 zn$3 \$140023 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7984 \$143086 z$26 \$143086 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7998 \$143087 z$26 \$143087 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7999 \$140024 zn$3 \$143087 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8000 \$140024 z$26 \$140024 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$8015 \$143088 zn$3 \$140024 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8016 \$143088 z$26 \$143088 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8031 \$143089 zn$3 \$140024 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8032 \$143089 z$26 \$143089 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8046 \$143090 z$26 \$143090 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8047 \$140025 zn$3 \$143090 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8048 \$140025 z$26 \$140025 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$8063 \$143091 zn$3 \$140025 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8064 \$143091 z$26 \$143091 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8079 \$143092 zn$3 \$140025 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8080 \$143092 z$26 \$143092 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8094 \$143093 z$26 \$143093 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8095 \$140026 zn$3 \$143093 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8096 \$140026 z$26 \$140026 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$8111 \$143094 zn$3 \$140026 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8112 \$143094 z$26 \$143094 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8127 \$143095 zn$3 \$140026 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8128 \$143095 z$26 \$143095 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8130 \$145299 \$145611 \$145299 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$8142 \$143096 z$26 \$143096 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8143 \$140027 zn$3 \$143096 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8144 \$140027 z$26 \$140027 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$8159 \$143097 zn$3 \$140027 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8160 \$143097 z$26 \$143097 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8175 \$143098 zn$3 \$140027 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8176 \$143098 z$26 \$143098 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8178 VSS|anode|cathode|clk|vss \$141285 \$142911 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$8179 \$142911 d|zn$5 \$141286 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$8180 \$141286 \$141594 \$142909 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$8181 VSS|anode|cathode|clk|vss \$141595 \$142909 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$8182 VSS|anode|cathode|clk|vss \$141286 \$141595 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$8183 \$141595 \$141594 \$142757 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$8184 \$142757 \$141285 \$142907 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$8185 VSS|anode|cathode|clk|vss \$141596 \$142907 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$8186 VSS|anode|cathode|clk|vss \$142757 \$141596 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$8187 \$143030 a2|a3|zn b|zn$5 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$8188 b|zn$5 RST|a1|b|cdn|core|i|p2c \$143030 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$8189 \$143030 a1|b|i|q$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$8550 \$145049 \$144246 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$8551 VSS|anode|cathode|clk|vss cp|z$3 \$144246 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$8552 VSS|anode|cathode|clk|vss \$144246 \$146158 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$8553 \$146158 d|z$4 \$144248 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$8554 \$144248 \$145049 \$146157 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$8555 VSS|anode|cathode|clk|vss \$144249 \$146157 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$8556 VSS|anode|cathode|clk|vss \$144248 \$144249 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$8557 \$144249 \$145049 \$145612 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$8558 \$145612 \$144246 \$146160 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$8559 VSS|anode|cathode|clk|vss \$145050 \$146160 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$8560 VSS|anode|cathode|clk|vss \$145612 \$145050 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$8561 a1|z$3 \$146514 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$8562 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$146514
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p
+ PS=1.55u PD=1.55u
M$8563 \$146514 a1|i|q \$146908 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$8564 \$146908 a2|z$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$8565 \$146314 a1|z$3 \$146913 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$8566 \$146913 a2|z$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.655u AS=0.271825p AD=0.2901875p PS=1.485u PD=1.55u
M$8567 VSS|anode|cathode|clk|vss \$146314 d|z$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2901875p AD=0.4068p PS=1.55u PD=2.57u
M$8568 b|i|q$2 \$145050 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$8569 \$146315 cp|i|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$8570 VSS|anode|cathode|clk|vss \$146315 cp|z$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$8571 \$150121 \$150578 \$150121 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$8583 \$148728 z$26 \$148728 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8584 \$145605 zn$3 \$148728 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8585 \$145605 z$26 \$145605 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$8600 \$148729 zn$3 \$145605 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8601 \$148729 z$26 \$148729 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8616 \$148730 zn$3 \$145605 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8617 \$148730 z$26 \$148730 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8631 a2$1 z$3 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8632 \$145606 z$1 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=11.52u AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$8633 \$145606 z$3 \$145606 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8647 \$145606 z$7 \$145606 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8648 VIN|core|padres z$4 \$145606 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$8649 VIN|core|padres z$7 VIN|core|padres VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8663 \$145606 z$27 \$145606 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8664 VIP|core|padres zn$5 \$145606 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$8665 VIP|core|padres z$27 VIP|core|padres VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8679 VREFL|core|padres z$7 VREFL|core|padres VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8680 \$145607 z$4 VREFL|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8681 \$145607 z$7 \$145607 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$8695 \$145607 z$9 \$145607 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$8696 a2$1 z \$145607 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8697 a2$1 z$9 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$8711 \$145607 z$8 \$145607 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$8712 a2 z$5 \$145607 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8713 a2 z$8 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$8715 \$150122 \$150579 \$150122 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=207.36u AS=88.6464p AD=88.6464p PS=470.88u PD=470.88u
M$8728 \$145608 z$4 VREFL|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$8729 \$145608 z$7 \$145608 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8743 \$145608 z$14 \$145608 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8744 a2$1 z$15 \$145608 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$8745 a2$1 z$14 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8759 \$145608 z$18 \$145608 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8760 a2 z$19 \$145608 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$8761 a2 z$18 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8776 \$145609 z$4 VREFL|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8777 \$145609 z$7 \$145609 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8791 \$145609 z$16 \$145609 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8792 a2$1 z$25 \$145609 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8793 a2$1 z$16 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8807 \$145609 z$21 \$145609 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8808 a2 z$23 \$145609 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8809 a2 z$21 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8824 \$145610 z$4 VREFL|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8825 \$145610 z$7 \$145610 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8839 \$145610 z$24 \$145610 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8840 a2$1 zn$4 \$145610 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8841 a2$1 z$24 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8856 a2 zn$4 \$145610 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8857 a2 z$24 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9003 \$150123 \$150580 \$150123 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$9015 \$148731 z$26 \$148731 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9016 \$145611 zn$3 \$148731 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9017 \$145611 z$26 \$145611 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$9032 \$148732 zn$3 \$145611 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9033 \$148732 z$26 \$148732 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9048 \$148733 zn$3 \$145611 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9049 \$148733 z$26 \$148733 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9051 a2|z$6 \$149324 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$9052 VSS|anode|cathode|clk|vss b|i|q$1 \$149324 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9053 \$149324 a1|i|q$1 \$149357 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9054 \$149357 a2|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$9055 \$148957 a2|zn$3 d|zn$9 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$9056 d|zn$9 a1|z$9 \$148957 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9057 \$148957 b|zn$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$9418 \$150581 a1|z$3 \$151835 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$9419 VSS|anode|cathode|clk|vss a2|z$3 \$151835 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.655u AS=0.2901875p AD=0.271825p PS=1.55u PD=1.485u
M$9420 VSS|anode|cathode|clk|vss \$150581 d|z$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2901875p AD=0.4068p PS=1.55u PD=2.57u
M$9421 \$152106 a2|a3|zn b|zn$6 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$9422 b|zn$6 RST|a1|b|cdn|core|i|p2c \$152106 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9423 \$152106 a1|b|i|q$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$9424 \$153380 z$26 \$153380 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9425 \$150578 zn$3 \$153380 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9426 \$150578 z$26 \$150578 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$9429 \$153381 zn$3 \$150578 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9430 \$153381 z$26 \$153381 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9433 \$153382 zn$3 \$150578 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9434 \$153382 z$26 \$153382 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9461 \$150579 z$4 VREFL|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$9462 \$150579 z$7 \$150579 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$9464 \$150579 z$12 \$150579 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$9465 a2$1 z$11 \$150579 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$9466 a2$1 z$12 a2$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$9468 \$150579 z$10 \$150579 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$9469 a2 z$13 \$150579 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$9470 a2 z$10 a2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$9532 \$153383 z$26 \$153383 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9533 \$150580 zn$3 \$153383 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9534 \$150580 z$26 \$150580 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$9537 \$153384 zn$3 \$150580 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9538 \$153384 z$26 \$153384 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9541 \$153385 zn$3 \$150580 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9542 \$153385 z$26 \$153385 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9544 a1|z$13 RESULT[0]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$9545 a2|z$7 \$155174 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$9546 VSS|anode|cathode|clk|vss b|i|q$3 \$155174 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9547 \$155174 a1|b|i|q$3 \$155223 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9548 \$155223 a2|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$9549 \$154584 a2|zn$3 d|zn$10 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$9550 d|zn$10 a1|z$1 \$154584 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9551 \$154584 b|zn$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$9552 a1|z RESULT[4]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$9553 \$155172 \$155875 \$155172 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$9877 \$155173 \$155876 \$155173 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$10273 a2|zn$1 a1|b|i|q$1 \$157750 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$10274 \$157750 a1|a2|a3|z \$157749 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$10275 \$157749 a2|a3|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$10276 \$159177 z$26 \$159177 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10277 \$155875 zn$3 \$159177 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10278 \$155875 z$26 \$155875 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$10281 \$159178 zn$3 \$155875 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10282 \$159178 z$26 \$159178 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10285 \$159179 zn$3 \$155875 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10286 \$159179 z$26 \$159179 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10384 \$159180 z$26 \$159180 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10385 \$155876 zn$3 \$159180 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10386 \$155876 z$26 \$155876 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$10389 \$159181 zn$3 \$155876 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10390 \$159181 z$26 \$159181 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10393 \$159182 zn$3 \$155876 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10394 \$159182 z$26 \$159182 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10396 \$158510 \$157993 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$10397 VSS|anode|cathode|clk|vss cp|z$3 \$157993 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$10398 \$157994 \$158510 \$158513 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$10399 \$158513 \$158244 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$10400 \$157995 \$157993 \$158514 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$10401 \$158514 \$158511 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$10402 \$158244 \$158510 \$157995 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$10403 VSS|anode|cathode|clk|vss \$157993 \$158512 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$10404 \$158512 a2|d|zn \$157994 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$10405 VSS|anode|cathode|clk|vss \$157994 \$158244 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$10406 VSS|anode|cathode|clk|vss \$157995 \$158511 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$10407 a2|zn$2 a1|b|i|q \$160947 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$10408 \$160947 a1|a2|a3|z \$160948 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$10409 \$160948 a2|a3|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$10410 a1|i|q \$158511 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$10411 \$160833 \$161529 \$160833 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$10735 \$160834 \$161530 \$160834 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11131 VSS|anode|cathode|clk|vss a2|zn$4 \$161652 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$11132 \$161652 a1|z$8 d|zn$7 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$11133 d|zn$7 b|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$11134 VSS|anode|cathode|clk|vss a2|a3|zn a2|d|zn VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$11135 a2|d|zn RST|a1|b|cdn|core|i|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p
+ PS=1.55u PD=2.57u
M$11136 \$164854 z$26 \$164854 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11137 \$161529 zn$3 \$164854 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11138 \$161529 z$26 \$161529 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$11141 \$164855 zn$3 \$161529 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11142 \$164855 z$26 \$164855 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11145 \$164856 zn$3 \$161529 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11146 \$164856 z$26 \$164856 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11244 \$164857 z$26 \$164857 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11245 \$161530 zn$3 \$164857 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11246 \$161530 z$26 \$161530 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$11249 \$164858 zn$3 \$161530 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11250 \$164858 z$26 \$164858 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11253 \$164859 zn$3 \$161530 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11254 \$164859 z$26 \$164859 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11256 \$164152 a2|zn$3 d|zn$8 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$11257 d|zn$8 a1|z$2 \$164152 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$11258 \$164152 b|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$11259 \$164860 a2|a3|zn b|zn$3 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$11260 b|zn$3 RST|a1|b|cdn|core|i|p2c \$164860 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$11261 \$164860 a1|b|i|q$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$11262 a2|zn$3 a1|i|q \$164315 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$11263 \$164315 a2|z$2 \$164316 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$11264 \$164316 a1|a2|a3|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$11265 a1|z$7 a1|i|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$11266 \$166600 \$167242 \$166600 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11302 \$166601 \$167243 \$166601 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11338 \$166602 \$167244 \$166602 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11374 \$166603 \$167245 \$166603 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11410 \$166604 \$167246 \$166604 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11446 \$166605 \$167247 \$166605 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11482 \$166606 \$167248 \$166606 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11518 \$166607 \$167249 \$166607 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11554 \$166608 \$167250 \$166608 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11590 \$166609 \$167251 \$166609 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11986 \$169906 z$26 \$169906 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11987 \$167242 zn$3 \$169906 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11988 \$167242 z$26 \$167242 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$11991 \$169907 zn$3 \$167242 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11992 \$169907 z$26 \$169907 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11995 \$169908 zn$3 \$167242 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11996 \$169908 z$26 \$169908 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11998 \$169909 z$26 \$169909 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11999 \$167243 zn$3 \$169909 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12000 \$167243 z$26 \$167243 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12003 \$169910 zn$3 \$167243 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12004 \$169910 z$26 \$169910 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12007 \$169911 zn$3 \$167243 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12008 \$169911 z$26 \$169911 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12010 \$169912 z$26 \$169912 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12011 \$167244 zn$3 \$169912 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12012 \$167244 z$26 \$167244 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12015 \$169913 zn$3 \$167244 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12016 \$169913 z$26 \$169913 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12019 \$169914 zn$3 \$167244 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12020 \$169914 z$26 \$169914 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12022 \$169915 z$26 \$169915 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12023 \$167245 zn$3 \$169915 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12024 \$167245 z$26 \$167245 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12027 \$169916 zn$3 \$167245 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12028 \$169916 z$26 \$169916 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12031 \$169917 zn$3 \$167245 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12032 \$169917 z$26 \$169917 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12034 \$169918 z$26 \$169918 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12035 \$167246 zn$3 \$169918 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12036 \$167246 z$26 \$167246 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12039 \$169919 zn$3 \$167246 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12040 \$169919 z$26 \$169919 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12043 \$169920 zn$3 \$167246 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12044 \$169920 z$26 \$169920 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12046 \$169921 z$26 \$169921 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12047 \$167247 zn$3 \$169921 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12048 \$167247 z$26 \$167247 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12051 \$169922 zn$3 \$167247 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12052 \$169922 z$26 \$169922 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12055 \$169923 zn$3 \$167247 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12056 \$169923 z$26 \$169923 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12058 \$169924 z$26 \$169924 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12059 \$167248 zn$3 \$169924 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12060 \$167248 z$26 \$167248 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12063 \$169925 zn$3 \$167248 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12064 \$169925 z$26 \$169925 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12067 \$169926 zn$3 \$167248 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12068 \$169926 z$26 \$169926 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12070 \$169927 z$26 \$169927 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12071 \$167249 zn$3 \$169927 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12072 \$167249 z$26 \$167249 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12075 \$169928 zn$3 \$167249 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12076 \$169928 z$26 \$169928 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12079 \$169929 zn$3 \$167249 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12080 \$169929 z$26 \$169929 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12082 \$169930 z$26 \$169930 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12083 \$167250 zn$3 \$169930 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12084 \$167250 z$26 \$167250 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12087 \$169931 zn$3 \$167250 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12088 \$169931 z$26 \$169931 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12091 \$169932 zn$3 \$167250 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12092 \$169932 z$26 \$169932 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12094 \$169933 z$26 \$169933 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12095 \$167251 zn$3 \$169933 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12096 \$167251 z$26 \$167251 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12099 \$169934 zn$3 \$167251 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12100 \$169934 z$26 \$169934 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12103 \$169935 zn$3 \$167251 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12104 \$169935 z$26 \$169935 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12106 a1|z$9 a1|i|q$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$12107 a1|z$10 a1|b|i|q$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$12108 VSS|anode|cathode|clk|vss a2|a3|z a2|zn$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$12109 a2|zn$5 RST|a1|b|cdn|core|i|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p
+ PS=1.55u PD=2.57u
M$12110 a1|z$4 RESULT[3]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$12111 RD[8]|a4|z \$181364 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12112 VSS|anode|cathode|clk|vss VALID|a3|c2p|core|i|z \$181364
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$12113 RD[9]|a4|z \$181365 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12114 VSS|anode|cathode|clk|vss SAMPLE|a1|c2p|core|i|z \$181365
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$12115 \$198889 DOUT_DAT|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$12116 \$200224 DOUT_DAT|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$12117 VSS|anode|cathode|clk|vss a1|a2|q \$207820 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12118 \$207820 a1|b|d|z \$207273 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12119 VSS|anode|cathode|clk|vss \$207273 d|z$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12120 VSS|anode|cathode|clk|vss cp|i|z$2 \$207275 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12121 VSS|anode|cathode|clk|vss \$207275 \$207253 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12122 \$207276 \$207253 \$207543 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12123 \$207543 \$207277 \$207541 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12124 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207541
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12125 \$207254 \$207275 \$207278 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12126 VSS|anode|cathode|clk|vss \$207275 \$207544 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12127 \$207544 d|z$14 \$207276 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12128 VSS|anode|cathode|clk|vss \$207276 \$207277 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12129 \$207277 \$207253 \$207254 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12130 VSS|anode|cathode|clk|vss \$207279 \$207278 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12131 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207828
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12132 \$207828 \$207254 \$207279 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12133 VSS|anode|cathode|clk|vss \$207279 a2|q$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12134 VSS|anode|cathode|clk|vss a2|i|q$1 \$207832 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12135 \$207832 a1|b|d|z \$207280 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12136 VSS|anode|cathode|clk|vss \$207280 d|z$6 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12137 VSS|anode|cathode|clk|vss cp|i|z$2 \$207282 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12138 VSS|anode|cathode|clk|vss \$207282 \$207255 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12139 \$207283 \$207255 \$207554 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12140 \$207554 \$207284 \$207565 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12141 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207565
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12142 \$207256 \$207282 \$207285 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12143 VSS|anode|cathode|clk|vss \$207282 \$207555 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12144 \$207555 d|z$15 \$207283 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12145 VSS|anode|cathode|clk|vss \$207283 \$207284 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12146 \$207284 \$207255 \$207256 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12147 VSS|anode|cathode|clk|vss \$207286 \$207285 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12148 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207835
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12149 \$207835 \$207256 \$207286 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12150 VSS|anode|cathode|clk|vss \$207286 a2|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12151 VSS|anode|cathode|clk|vss a1|a2|q$1 a3|zn VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12152 a3|zn a2|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12153 VSS|anode|cathode|clk|vss a2|q$2 \$207837 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12154 \$207837 a1|b|d|z \$207287 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12155 VSS|anode|cathode|clk|vss \$207287 d|z$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12156 VSS|anode|cathode|clk|vss a2|q$1 \$207838 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12157 \$207838 a1|b|d|z \$207289 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12158 VSS|anode|cathode|clk|vss \$207289 d|z$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12159 VSS|anode|cathode|clk|vss cp|i|z$3 \$207291 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12160 VSS|anode|cathode|clk|vss \$207291 \$207257 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12161 \$207292 \$207257 \$207569 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12162 \$207569 \$207293 \$207576 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12163 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207576
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12164 \$207258 \$207291 \$207294 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12165 VSS|anode|cathode|clk|vss \$207291 \$207570 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12166 \$207570 d|z$16 \$207292 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12167 VSS|anode|cathode|clk|vss \$207292 \$207293 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12168 \$207293 \$207257 \$207258 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12169 VSS|anode|cathode|clk|vss \$207295 \$207294 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12170 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207841
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12171 \$207841 \$207258 \$207295 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12172 VSS|anode|cathode|clk|vss \$207295 a1|a2|q$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12173 VSS|anode|cathode|clk|vss a1|a2|q$2 \$207840 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12174 \$207840 a1|b|d|z \$207296 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12175 VSS|anode|cathode|clk|vss \$207296 d|z$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12176 \$207298 s|zn \$207299 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12177 \$207300 \$207260 \$207298 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12178 VSS|anode|cathode|clk|vss i0|i1|q \$207300 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12179 VSS|anode|cathode|clk|vss R[32]|i1|q \$207299 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12180 VSS|anode|cathode|clk|vss s|zn \$207260 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12181 VSS|anode|cathode|clk|vss \$207298 d|z$10 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12182 \$207302 s|z \$207303 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12183 \$207305 \$207262 \$207302 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12184 VSS|anode|cathode|clk|vss R[28]|i0|q \$207305 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12185 VSS|anode|cathode|clk|vss i0|i1|q$5 \$207303 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12186 VSS|anode|cathode|clk|vss s|z \$207262 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12187 VSS|anode|cathode|clk|vss \$207302 d|z$11 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12188 VSS|anode|cathode|clk|vss cp|i|z$4 \$207307 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12189 VSS|anode|cathode|clk|vss \$207307 \$207263 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12190 \$207308 \$207263 \$207559 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12191 \$207559 \$207309 \$207560 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12192 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207560
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12193 \$207264 \$207307 \$207310 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12194 VSS|anode|cathode|clk|vss \$207307 \$207568 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12195 \$207568 d|z$11 \$207308 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12196 VSS|anode|cathode|clk|vss \$207308 \$207309 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12197 \$207309 \$207263 \$207264 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12198 VSS|anode|cathode|clk|vss \$207311 \$207310 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12199 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207869
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12200 \$207869 \$207264 \$207311 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12201 VSS|anode|cathode|clk|vss \$207311 R[28]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12202 \$207312 s|z \$207313 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12203 \$207314 \$207265 \$207312 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12204 VSS|anode|cathode|clk|vss R[25]|i0|q \$207314 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12205 VSS|anode|cathode|clk|vss i0|i1|q$6 \$207313 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12206 VSS|anode|cathode|clk|vss s|z \$207265 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12207 VSS|anode|cathode|clk|vss \$207312 d|z$12 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12208 VSS|anode|cathode|clk|vss cp|i|z$1 \$207316 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12209 VSS|anode|cathode|clk|vss \$207316 \$207266 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12210 \$207317 \$207266 \$207547 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12211 \$207547 \$207318 \$207549 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12212 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207549
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12213 \$207267 \$207316 \$207319 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12214 VSS|anode|cathode|clk|vss \$207316 \$207556 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12215 \$207556 d|z$17 \$207317 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12216 VSS|anode|cathode|clk|vss \$207317 \$207318 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12217 \$207318 \$207266 \$207267 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12218 VSS|anode|cathode|clk|vss \$207320 \$207319 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12219 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207924
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12220 \$207924 \$207267 \$207320 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12221 VSS|anode|cathode|clk|vss \$207320 R[27]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12222 VSS|anode|cathode|clk|vss cp|i|z$1 \$207321 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12223 VSS|anode|cathode|clk|vss \$207321 \$207268 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12224 \$207322 \$207268 \$207546 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12225 \$207546 \$207323 \$207536 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12226 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207536
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12227 \$207269 \$207321 \$207324 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12228 VSS|anode|cathode|clk|vss \$207321 \$207545 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12229 \$207545 d|z$18 \$207322 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12230 VSS|anode|cathode|clk|vss \$207322 \$207323 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12231 \$207323 \$207268 \$207269 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12232 VSS|anode|cathode|clk|vss \$207325 \$207324 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12233 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207970
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12234 \$207970 \$207269 \$207325 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12235 VSS|anode|cathode|clk|vss \$207325 R[33]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12236 VSS|anode|cathode|clk|vss cp|i|z$1 \$207326 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12237 VSS|anode|cathode|clk|vss \$207326 \$207270 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12238 \$207327 \$207270 \$207535 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12239 \$207535 \$207328 \$207524 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12240 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$207524
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12241 \$207271 \$207326 \$207329 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12242 VSS|anode|cathode|clk|vss \$207326 \$207534 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12243 \$207534 d|z$19 \$207327 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12244 VSS|anode|cathode|clk|vss \$207327 \$207328 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12245 \$207328 \$207270 \$207271 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12246 VSS|anode|cathode|clk|vss \$207330 \$207329 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12247 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$208011
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12248 \$208011 \$207271 \$207330 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12249 VSS|anode|cathode|clk|vss \$207330 i0|i1|q$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12250 \$207331 s|zn$1 \$207332 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12251 \$207333 \$207272 \$207331 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12252 VSS|anode|cathode|clk|vss i0|i1|q$5 \$207333 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12253 VSS|anode|cathode|clk|vss i0|i1|q$7 \$207332 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12254 VSS|anode|cathode|clk|vss s|zn$1 \$207272 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12255 VSS|anode|cathode|clk|vss \$207331 d|z$13 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12256 VSS|anode|cathode|clk|vss \$210072 \$211083 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12257 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211146
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12258 \$211146 \$209540 \$210072 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12259 VSS|anode|cathode|clk|vss \$210072 a1|a2|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12260 VSS|anode|cathode|clk|vss a1|a2|q$4 a2|zn$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12261 a2|zn$7 a2|q$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12262 d|z$20 \$209542 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12263 VSS|anode|cathode|clk|vss \$210075 \$211084 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12264 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211150
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12265 \$211150 \$209549 \$210075 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12266 VSS|anode|cathode|clk|vss \$210075 a2|i|q$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12267 d|z$21 \$209550 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12268 d|z$22 \$209552 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12269 VSS|anode|cathode|clk|vss \$210077 \$211085 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12270 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211162
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12271 \$211162 \$209559 \$210077 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12272 VSS|anode|cathode|clk|vss \$210077 a2|q$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12273 VSS|anode|cathode|clk|vss \$210078 \$211086 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12274 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211171
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12275 \$211171 \$209566 \$210078 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12276 VSS|anode|cathode|clk|vss \$210078 a1|a2|q$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12277 VSS|anode|cathode|clk|vss \$210079 \$211087 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12278 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211179
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12279 \$211179 \$209573 \$210079 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12280 VSS|anode|cathode|clk|vss \$210079 a2|q$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12281 VSS|anode|cathode|clk|vss \$210080 \$211088 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12282 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211181
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12283 \$211181 \$209579 \$210080 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12284 VSS|anode|cathode|clk|vss \$210080 R[32]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12285 \$209581 s|z \$209580 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12286 \$209581 i0|i1|q$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12287 VSS|anode|cathode|clk|vss R[26]|i0|q \$209582 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12288 \$209582 \$209149 \$209580 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12289 VSS|anode|cathode|clk|vss s|z \$209149 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12290 VSS|anode|cathode|clk|vss \$209580 d|z$23 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12291 VSS|anode|cathode|clk|vss \$210083 \$211089 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12292 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211173
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12293 \$211173 \$209589 \$210083 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12294 VSS|anode|cathode|clk|vss \$210083 R[26]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12295 VSS|anode|cathode|clk|vss \$210084 \$211090 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12296 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211172
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12297 \$211172 \$209595 \$210084 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12298 VSS|anode|cathode|clk|vss \$210084 R[25]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12299 VSS|anode|cathode|clk|vss \$210086 \$211091 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12300 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211158
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12301 \$211158 \$209601 \$210086 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12302 VSS|anode|cathode|clk|vss \$210086 R[24]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12303 VSS|anode|cathode|clk|vss \$210088 \$211092 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12304 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211145
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12305 \$211145 \$209608 \$210088 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12306 VSS|anode|cathode|clk|vss \$210088 R[34]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12307 VSS|anode|cathode|clk|vss \$210090 \$211093 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12308 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211144
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12309 \$211144 \$209615 \$210090 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12310 VSS|anode|cathode|clk|vss \$210090 i0|i1|q$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12311 VSS|anode|cathode|clk|vss \$210092 \$211094 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12312 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211134
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12313 \$211134 \$209621 \$210092 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12314 VSS|anode|cathode|clk|vss \$210092 i0|i1|q$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12315 VSS|anode|cathode|clk|vss \$210093 \$211095 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12316 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211130
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12317 \$211130 \$209627 \$210093 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12318 VSS|anode|cathode|clk|vss \$210093 i0|i1|q$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12319 \$209535 cp|i|z$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12320 VSS|anode|cathode|clk|vss \$209535 \$209536 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12321 VSS|anode|cathode|clk|vss \$209535 \$211143 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12322 \$211143 d|z$24 \$209537 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12323 \$209537 \$209536 \$211142 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12324 \$211142 \$209539 \$211141 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12325 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211141
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12326 \$209539 \$209537 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12327 \$209539 \$209536 \$209540 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12328 \$209540 \$209535 \$211083 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12329 VSS|anode|cathode|clk|vss a2|q$3 \$211148 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12330 \$211148 a1|b|d|z \$209542 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12331 \$209544 cp|i|z$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12332 VSS|anode|cathode|clk|vss \$209544 \$209545 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12333 VSS|anode|cathode|clk|vss \$209544 \$211147 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12334 \$211147 d|z$20 \$209546 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12335 \$209546 \$209545 \$211154 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12336 \$211154 \$209548 \$211153 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12337 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211153
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12338 \$209548 \$209546 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12339 \$209548 \$209545 \$209549 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12340 \$209549 \$209544 \$211084 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12341 VSS|anode|cathode|clk|vss a1|a2|q$5 \$211157 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12342 \$211157 a1|b|d|z \$209550 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12343 VSS|anode|cathode|clk|vss a2|q \$211156 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12344 \$211156 a1|b|d|z \$209552 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12345 \$209554 cp|i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12346 VSS|anode|cathode|clk|vss \$209554 \$209555 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12347 VSS|anode|cathode|clk|vss \$209554 \$211161 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12348 \$211161 d|z$22 \$209556 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12349 \$209556 \$209555 \$211160 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12350 \$211160 \$209558 \$211159 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12351 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211159
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12352 \$209558 \$209556 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12353 \$209558 \$209555 \$209559 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12354 \$209559 \$209554 \$211085 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12355 \$209561 cp|i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12356 VSS|anode|cathode|clk|vss \$209561 \$209562 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12357 VSS|anode|cathode|clk|vss \$209561 \$211168 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12358 \$211168 d|z$7 \$209563 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12359 \$209563 \$209562 \$211167 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12360 \$211167 \$209565 \$211166 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12361 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211166
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12362 \$209565 \$209563 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12363 \$209565 \$209562 \$209566 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12364 \$209566 \$209561 \$211086 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12365 \$209568 cp|i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12366 VSS|anode|cathode|clk|vss \$209568 \$209569 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12367 VSS|anode|cathode|clk|vss \$209568 \$211176 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12368 \$211176 d|z$9 \$209570 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12369 \$209570 \$209569 \$211175 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12370 \$211175 \$209572 \$211174 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12371 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211174
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12372 \$209572 \$209570 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12373 \$209572 \$209569 \$209573 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12374 \$209573 \$209568 \$211087 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12375 \$209574 cp|i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12376 VSS|anode|cathode|clk|vss \$209574 \$209575 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12377 VSS|anode|cathode|clk|vss \$209574 \$211177 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12378 \$211177 d|z$10 \$209576 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12379 \$209576 \$209575 \$211185 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12380 \$211185 \$209578 \$211184 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12381 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211184
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12382 \$209578 \$209576 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12383 \$209578 \$209575 \$209579 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12384 \$209579 \$209574 \$211088 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12385 \$209584 cp|i|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12386 VSS|anode|cathode|clk|vss \$209584 \$209585 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12387 VSS|anode|cathode|clk|vss \$209584 \$211180 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12388 \$211180 d|z$23 \$209586 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12389 \$209586 \$209585 \$211182 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12390 \$211182 \$209588 \$211183 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12391 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211183
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12392 \$209588 \$209586 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12393 \$209588 \$209585 \$209589 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12394 \$209589 \$209584 \$211089 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12395 \$209590 cp|i|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12396 VSS|anode|cathode|clk|vss \$209590 \$209591 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12397 VSS|anode|cathode|clk|vss \$209590 \$211178 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12398 \$211178 d|z$12 \$209592 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12399 \$209592 \$209591 \$211169 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12400 \$211169 \$209594 \$211170 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12401 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211170
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12402 \$209594 \$209592 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12403 \$209594 \$209591 \$209595 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12404 \$209595 \$209590 \$211090 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12405 \$209596 cp|i|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12406 VSS|anode|cathode|clk|vss \$209596 \$209597 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12407 VSS|anode|cathode|clk|vss \$209596 \$211163 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12408 \$211163 d|z$25 \$209598 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12409 \$209598 \$209597 \$211164 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12410 \$211164 \$209600 \$211165 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12411 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211165
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12412 \$209600 \$209598 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12413 \$209600 \$209597 \$209601 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12414 \$209601 \$209596 \$211091 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12415 \$209603 cp|i|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12416 VSS|anode|cathode|clk|vss \$209603 \$209604 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12417 VSS|anode|cathode|clk|vss \$209603 \$211151 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12418 \$211151 d|z$26 \$209605 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12419 \$209605 \$209604 \$211152 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12420 \$211152 \$209607 \$211155 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12421 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211155
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12422 \$209607 \$209605 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12423 \$209607 \$209604 \$209608 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12424 \$209608 \$209603 \$211092 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12425 \$209610 cp|i|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12426 VSS|anode|cathode|clk|vss \$209610 \$209611 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12427 VSS|anode|cathode|clk|vss \$209610 \$211149 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12428 \$211149 d|z$27 \$209612 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12429 \$209612 \$209611 \$211139 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12430 \$211139 \$209614 \$211140 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12431 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211140
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12432 \$209614 \$209612 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12433 \$209614 \$209611 \$209615 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12434 \$209615 \$209610 \$211093 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12435 \$209616 cp|i|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12436 VSS|anode|cathode|clk|vss \$209616 \$209617 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12437 VSS|anode|cathode|clk|vss \$209616 \$211136 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12438 \$211136 d|z$28 \$209618 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12439 \$209618 \$209617 \$211137 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12440 \$211137 \$209620 \$211138 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12441 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211138
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12442 \$209620 \$209618 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12443 \$209620 \$209617 \$209621 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12444 \$209621 \$209616 \$211094 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12445 \$209622 cp|i|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12446 VSS|anode|cathode|clk|vss \$209622 \$209623 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12447 VSS|anode|cathode|clk|vss \$209622 \$211131 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12448 \$211131 d|z$13 \$209624 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12449 \$209624 \$209623 \$211132 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12450 \$211132 \$209626 \$211133 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12451 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211133
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12452 \$209626 \$209624 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12453 \$209626 \$209623 \$209627 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12454 \$209627 \$209622 \$211095 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12455 VSS|anode|cathode|clk|vss cp|i|z$2 \$211694 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12456 VSS|anode|cathode|clk|vss \$211694 \$211695 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12457 \$211696 \$211695 \$211840 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12458 \$211840 \$211697 \$211839 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12459 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211839
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12460 \$211698 \$211694 \$211699 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12461 VSS|anode|cathode|clk|vss \$211694 \$211841 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12462 \$211841 d|z$5 \$211696 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12463 VSS|anode|cathode|clk|vss \$211696 \$211697 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12464 \$211697 \$211695 \$211698 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12465 VSS|anode|cathode|clk|vss \$211700 \$211699 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12466 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212102
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12467 \$212102 \$211698 \$211700 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12468 VSS|anode|cathode|clk|vss \$211700 a2|q$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12469 VSS|anode|cathode|clk|vss cp|i|z$2 \$211701 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12470 VSS|anode|cathode|clk|vss \$211701 \$211702 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12471 \$211703 \$211702 \$211846 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12472 \$211846 \$211704 \$211845 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12473 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211845
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12474 \$211705 \$211701 \$211706 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12475 VSS|anode|cathode|clk|vss \$211701 \$211847 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12476 \$211847 d|z$29 \$211703 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12477 VSS|anode|cathode|clk|vss \$211703 \$211704 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12478 \$211704 \$211702 \$211705 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12479 VSS|anode|cathode|clk|vss \$211707 \$211706 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12480 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212147
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12481 \$212147 \$211705 \$211707 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12482 VSS|anode|cathode|clk|vss \$211707 a1|a2|q$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12483 VSS|anode|cathode|clk|vss i|z$115 \$211708 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12484 VSS|anode|cathode|clk|vss \$211708 cp|i|z$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12485 VSS|anode|cathode|clk|vss cp|i|z$2 \$211709 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12486 VSS|anode|cathode|clk|vss \$211709 \$211710 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12487 \$211711 \$211710 \$211853 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12488 \$211853 \$211712 \$211851 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12489 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211851
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12490 \$211713 \$211709 \$211714 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12491 VSS|anode|cathode|clk|vss \$211709 \$211856 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12492 \$211856 d|z$6 \$211711 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12493 VSS|anode|cathode|clk|vss \$211711 \$211712 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12494 \$211712 \$211710 \$211713 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12495 VSS|anode|cathode|clk|vss \$211715 \$211714 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12496 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212214
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12497 \$212214 \$211713 \$211715 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12498 VSS|anode|cathode|clk|vss \$211715 a1|a2|q$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12499 VSS|anode|cathode|clk|vss cp|i|z$2 \$211716 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12500 VSS|anode|cathode|clk|vss \$211716 \$211717 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12501 \$211718 \$211717 \$211861 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12502 \$211861 \$211719 \$211860 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12503 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211860
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12504 \$211720 \$211716 \$211721 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12505 VSS|anode|cathode|clk|vss \$211716 \$211862 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12506 \$211862 d|z$21 \$211718 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12507 VSS|anode|cathode|clk|vss \$211718 \$211719 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12508 \$211719 \$211717 \$211720 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12509 VSS|anode|cathode|clk|vss \$211722 \$211721 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12510 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212256
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12511 \$212256 \$211720 \$211722 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12512 VSS|anode|cathode|clk|vss \$211722 a1|a2|q$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12513 VSS|anode|cathode|clk|vss a1|a2|q$5 a4|zn VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12514 a4|zn a2|q$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12515 \$211724 a3|zn \$212265 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12516 \$212265 a2|zn$8 \$212305 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12517 \$212305 a1|zn a2|zn$9 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12518 VSS|anode|cathode|clk|vss a4|zn \$211724 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12519 VSS|anode|cathode|clk|vss a1|a2|q$3 \$212283 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12520 \$212283 a1|b|d|z \$211725 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12521 VSS|anode|cathode|clk|vss \$211725 d|z$16 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12522 VSS|anode|cathode|clk|vss cp|i|z$3 \$211726 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12523 VSS|anode|cathode|clk|vss \$211726 \$211727 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12524 \$211728 \$211727 \$211864 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12525 \$211864 \$211729 \$211865 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12526 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211865
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12527 \$211730 \$211726 \$211731 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12528 VSS|anode|cathode|clk|vss \$211726 \$211863 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12529 \$211863 d|z$8 \$211728 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12530 VSS|anode|cathode|clk|vss \$211728 \$211729 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12531 \$211729 \$211727 \$211730 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12532 VSS|anode|cathode|clk|vss \$211732 \$211731 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12533 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212370
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12534 \$212370 \$211730 \$211732 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12535 VSS|anode|cathode|clk|vss \$211732 a2|q$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12536 VSS|anode|cathode|clk|vss cp|i|z$3 \$211733 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12537 VSS|anode|cathode|clk|vss \$211733 \$211734 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12538 \$211735 \$211734 \$211858 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12539 \$211858 \$211736 \$211859 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12540 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211859
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12541 \$211737 \$211733 \$211738 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12542 VSS|anode|cathode|clk|vss \$211733 \$211857 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12543 \$211857 d|z$30 \$211735 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12544 VSS|anode|cathode|clk|vss \$211735 \$211736 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12545 \$211736 \$211734 \$211737 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12546 VSS|anode|cathode|clk|vss \$211739 \$211738 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12547 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212405
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12548 \$212405 \$211737 \$211739 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12549 VSS|anode|cathode|clk|vss \$211739 i0|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12550 VSS|anode|cathode|clk|vss cp|i|z$4 \$211740 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12551 VSS|anode|cathode|clk|vss \$211740 \$211741 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12552 \$211742 \$211741 \$211854 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12553 \$211854 \$211743 \$211855 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12554 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211855
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12555 \$211744 \$211740 \$211745 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12556 VSS|anode|cathode|clk|vss \$211740 \$211852 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12557 \$211852 d|z$31 \$211742 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12558 VSS|anode|cathode|clk|vss \$211742 \$211743 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12559 \$211743 \$211741 \$211744 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12560 VSS|anode|cathode|clk|vss \$211746 \$211745 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12561 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212446
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12562 \$212446 \$211744 \$211746 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12563 VSS|anode|cathode|clk|vss \$211746 R[29]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12564 VSS|anode|cathode|clk|vss cp|i|z$4 \$211747 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12565 VSS|anode|cathode|clk|vss \$211747 \$211748 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12566 \$211749 \$211748 \$211849 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12567 \$211849 \$211750 \$211850 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12568 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211850
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12569 \$211751 \$211747 \$211752 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12570 VSS|anode|cathode|clk|vss \$211747 \$211848 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12571 \$211848 d|z$32 \$211749 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12572 VSS|anode|cathode|clk|vss \$211749 \$211750 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12573 \$211750 \$211748 \$211751 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12574 VSS|anode|cathode|clk|vss \$211753 \$211752 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12575 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212465
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12576 \$212465 \$211751 \$211753 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12577 VSS|anode|cathode|clk|vss \$211753 R[36]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12578 \$211754 s|z \$211755 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12579 \$211756 \$211757 \$211754 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12580 VSS|anode|cathode|clk|vss R[24]|i0|q \$211756 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12581 VSS|anode|cathode|clk|vss i0|i1|q \$211755 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12582 VSS|anode|cathode|clk|vss s|z \$211757 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12583 VSS|anode|cathode|clk|vss \$211754 d|z$25 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12584 VSS|anode|cathode|clk|vss cp|i|z$4 \$211758 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12585 VSS|anode|cathode|clk|vss \$211758 \$211759 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12586 \$211760 \$211759 \$211843 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12587 \$211843 \$211761 \$211844 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12588 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211844
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12589 \$211762 \$211758 \$211763 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12590 VSS|anode|cathode|clk|vss \$211758 \$211842 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12591 \$211842 d|z$33 \$211760 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12592 VSS|anode|cathode|clk|vss \$211760 \$211761 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12593 \$211761 \$211759 \$211762 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12594 VSS|anode|cathode|clk|vss \$211764 \$211763 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12595 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212485
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12596 \$212485 \$211762 \$211764 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12597 VSS|anode|cathode|clk|vss \$211764 R[30]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12598 \$211765 s|z \$211766 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12599 \$211767 \$211768 \$211765 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12600 VSS|anode|cathode|clk|vss R[27]|i0|q \$211767 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12601 VSS|anode|cathode|clk|vss i0|i1|q$1 \$211766 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12602 VSS|anode|cathode|clk|vss s|z \$211768 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12603 VSS|anode|cathode|clk|vss \$211765 d|z$17 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12604 \$211769 s|zn \$211770 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12605 \$211771 \$211772 \$211769 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12606 VSS|anode|cathode|clk|vss i0|i1|q$2 \$211771 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12607 VSS|anode|cathode|clk|vss R[34]|i1|q \$211770 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12608 VSS|anode|cathode|clk|vss s|zn \$211772 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12609 VSS|anode|cathode|clk|vss \$211769 d|z$26 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12610 \$211773 s|zn$1 \$211775 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12611 \$211776 \$211777 \$211773 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12612 VSS|anode|cathode|clk|vss i0|i1|q$6 \$211776 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12613 VSS|anode|cathode|clk|vss i0|i1|q$2 \$211775 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12614 VSS|anode|cathode|clk|vss s|zn$1 \$211777 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12615 VSS|anode|cathode|clk|vss \$211773 d|z$27 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12616 \$211778 s|zn$1 \$211779 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12617 \$211780 \$211781 \$211778 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12618 VSS|anode|cathode|clk|vss i0|i1|q$2 \$211780 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12619 VSS|anode|cathode|clk|vss i0|i1|q$1 \$211779 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12620 VSS|anode|cathode|clk|vss s|zn$1 \$211781 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12621 VSS|anode|cathode|clk|vss \$211778 d|z$19 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12622 VSS|anode|cathode|clk|vss i|z$115 \$211782 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12623 VSS|anode|cathode|clk|vss \$211782 cp|i|z$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12624 z$28 cp|i|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12625 VSS|anode|cathode|clk|vss cp|i|z$1 \$211784 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12626 VSS|anode|cathode|clk|vss \$211784 \$211785 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12627 \$211786 \$211785 \$211834 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12628 \$211834 \$211787 \$211835 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12629 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211835
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12630 \$211788 \$211784 \$211789 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12631 VSS|anode|cathode|clk|vss \$211784 \$211836 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12632 \$211836 d|z$34 \$211786 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12633 VSS|anode|cathode|clk|vss \$211786 \$211787 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12634 \$211787 \$211785 \$211788 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12635 VSS|anode|cathode|clk|vss \$211790 \$211789 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12636 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212478
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12637 \$212478 \$211788 \$211790 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12638 VSS|anode|cathode|clk|vss \$211790 i0|i1|q$6 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12639 VSS|anode|cathode|clk|vss cp|i|z$1 \$211791 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12640 VSS|anode|cathode|clk|vss \$211791 \$211792 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12641 \$211793 \$211792 \$211830 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12642 \$211830 \$211794 \$211831 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12643 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$211831
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12644 \$211795 \$211791 \$211796 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12645 VSS|anode|cathode|clk|vss \$211791 \$211833 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12646 \$211833 d|z$35 \$211793 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12647 VSS|anode|cathode|clk|vss \$211793 \$211794 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12648 \$211794 \$211792 \$211795 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12649 VSS|anode|cathode|clk|vss \$211797 \$211796 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12650 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$212447
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12651 \$212447 \$211795 \$211797 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12652 VSS|anode|cathode|clk|vss \$211797 i0|i1|q$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12653 VSS|anode|cathode|clk|vss a2|q$6 \$215449 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12654 \$215449 a1|b|d|z \$213634 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12655 d|z$24 \$213634 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12656 VSS|anode|cathode|clk|vss \$214361 \$215224 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12657 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215454
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12658 \$215454 \$213640 \$214361 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12659 VSS|anode|cathode|clk|vss \$214361 a2|q$6 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12660 VSS|anode|cathode|clk|vss a1|a2|q$6 \$215471 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12661 \$215471 a1|b|d|z \$213642 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12662 d|z$38 \$213642 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12663 VSS|anode|cathode|clk|vss a1|a2|q$4 \$215469 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12664 \$215469 a1|b|d|z \$213643 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12665 d|z$14 \$213643 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12666 \$215225 a3|zn$1 \$215466 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12667 \$215466 a2|zn$7 \$215465 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12668 \$215465 a1|z$14 a2|zn$10 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12669 \$215225 a4|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12670 a1|z$14 a2|i|q$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12671 VSS|anode|cathode|clk|vss a1|b|d|z \$215226 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12672 \$215226 a1|zn$1 s|zn$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12673 s|zn$1 a2|zn$10 \$215226 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12674 VSS|anode|cathode|clk|vss \$214362 \$215227 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12675 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215482
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12676 \$215482 \$213650 \$214362 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12677 VSS|anode|cathode|clk|vss \$214362 a1|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12678 VSS|anode|cathode|clk|vss a1|a2|q$1 \$215479 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12679 \$215479 a1|b|d|z \$213652 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12680 d|z$15 \$213652 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12681 VSS|anode|cathode|clk|vss \$214363 \$215228 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12682 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215483
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12683 \$215483 \$213658 \$214363 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12684 VSS|anode|cathode|clk|vss \$214363 a1|i|i0|i1|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$12685 z$29 cp|i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12686 VSS|anode|cathode|clk|vss a1|a2|q$3 a2|zn$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12687 a2|zn$8 a2|q$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12688 cp|i|z$3 \$213661 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12689 VSS|anode|cathode|clk|vss i|z$115 \$213661 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12690 \$213663 s|zn$1 \$213662 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12691 \$213663 i0|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12692 VSS|anode|cathode|clk|vss DATA|core|i0|i1|p2c \$213664
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$12693 \$213664 \$213585 \$213662 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12694 VSS|anode|cathode|clk|vss s|zn$1 \$213585 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12695 VSS|anode|cathode|clk|vss \$213662 d|z$30 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12696 VSS|anode|cathode|clk|vss \$214364 \$215229 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12697 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215498
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12698 \$215498 \$213670 \$214364 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12699 VSS|anode|cathode|clk|vss \$214364 R[21]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12700 \$213673 s|z \$213672 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12701 \$213673 i0|i1|q$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12702 VSS|anode|cathode|clk|vss R[29]|i0|q \$213674 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12703 \$213674 \$213586 \$213672 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12704 VSS|anode|cathode|clk|vss s|z \$213586 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12705 VSS|anode|cathode|clk|vss \$213672 d|z$31 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12706 \$213676 s|zn \$213675 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12707 \$213676 R[39]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12708 VSS|anode|cathode|clk|vss i0|i1|q$4 \$213677 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12709 \$213677 \$213587 \$213675 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12710 VSS|anode|cathode|clk|vss s|zn \$213587 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12711 VSS|anode|cathode|clk|vss \$213675 d|z$36 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12712 \$213680 s|zn \$213679 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12713 \$213680 R[36]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12714 VSS|anode|cathode|clk|vss i0|i1|q$5 \$213681 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12715 \$213681 \$213588 \$213679 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12716 VSS|anode|cathode|clk|vss s|zn \$213588 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12717 VSS|anode|cathode|clk|vss \$213679 d|z$32 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12718 z$30 cp|i|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12719 cp|i|z$4 \$213683 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12720 VSS|anode|cathode|clk|vss i|z$115 \$213683 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12721 \$213685 s|z \$213684 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12722 \$213685 i0|i1|q$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12723 VSS|anode|cathode|clk|vss R[30]|i0|q \$213686 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12724 \$213686 \$213589 \$213684 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12725 VSS|anode|cathode|clk|vss s|z \$213589 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12726 VSS|anode|cathode|clk|vss \$213684 d|z$33 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12727 VSS|anode|cathode|clk|vss \$214367 \$215230 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12728 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215485
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12729 \$215485 \$213692 \$214367 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12730 VSS|anode|cathode|clk|vss \$214367 R[20]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12731 \$213695 s|zn \$213694 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12732 \$213695 R[33]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12733 VSS|anode|cathode|clk|vss i0|i1|q$6 \$213696 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12734 \$213696 \$213590 \$213694 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12735 VSS|anode|cathode|clk|vss s|zn \$213590 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12736 VSS|anode|cathode|clk|vss \$213694 d|z$18 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12737 \$213698 s|zn \$213697 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12738 \$213698 R[37]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12739 VSS|anode|cathode|clk|vss i0|i1|q$7 \$213699 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12740 \$213699 \$213591 \$213697 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12741 VSS|anode|cathode|clk|vss s|zn \$213591 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12742 VSS|anode|cathode|clk|vss \$213697 d|z$37 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12743 VSS|anode|cathode|clk|vss \$214369 \$215231 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12744 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215478
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12745 \$215478 \$213706 \$214369 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12746 VSS|anode|cathode|clk|vss \$214369 R[37]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12747 \$213709 s|zn$1 \$213708 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12748 \$213709 i0|i1|q$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12749 VSS|anode|cathode|clk|vss i0|i1|q$1 \$213710 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12750 \$213710 \$213592 \$213708 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12751 VSS|anode|cathode|clk|vss s|zn$1 \$213592 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12752 VSS|anode|cathode|clk|vss \$213708 d|z$28 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12753 \$213712 s|zn$1 \$213711 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12754 \$213712 i0|i1|q$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12755 VSS|anode|cathode|clk|vss i0|i1|q \$213713 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12756 \$213713 \$213593 \$213711 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12757 VSS|anode|cathode|clk|vss s|zn$1 \$213593 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12758 VSS|anode|cathode|clk|vss \$213711 d|z$34 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12759 VSS|anode|cathode|clk|vss \$214371 \$215232 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12760 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215458
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12761 \$215458 \$213719 \$214371 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12762 VSS|anode|cathode|clk|vss \$214371 i0|i1|q$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12763 \$213635 cp|i|z$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12764 VSS|anode|cathode|clk|vss \$213635 \$213636 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12765 VSS|anode|cathode|clk|vss \$213635 \$215463 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12766 \$215463 d|z$38 \$213637 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12767 \$213637 \$213636 \$215461 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12768 \$215461 \$213639 \$215460 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12769 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215460
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12770 \$213639 \$213637 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12771 \$213639 \$213636 \$213640 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12772 \$213640 \$213635 \$215224 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12773 \$213645 cp|i|z$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12774 VSS|anode|cathode|clk|vss \$213645 \$213646 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12775 VSS|anode|cathode|clk|vss \$213645 \$215474 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12776 \$215474 d|z$41 \$213647 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12777 \$213647 \$213646 \$215473 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12778 \$215473 \$213649 \$215472 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12779 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215472
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12780 \$213649 \$213647 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12781 \$213649 \$213646 \$213650 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12782 \$213650 \$213645 \$215227 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12783 \$213653 cp|i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12784 VSS|anode|cathode|clk|vss \$213653 \$213654 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12785 VSS|anode|cathode|clk|vss \$213653 \$215488 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12786 \$215488 d|z$42 \$213655 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12787 \$213655 \$213654 \$215487 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12788 \$215487 \$213657 \$215486 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12789 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215486
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12790 \$213657 \$213655 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12791 \$213657 \$213654 \$213658 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12792 \$213658 \$213653 \$215228 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12793 \$213665 cp|i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12794 VSS|anode|cathode|clk|vss \$213665 \$213666 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12795 VSS|anode|cathode|clk|vss \$213665 \$215496 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12796 \$215496 d|z$39 \$213667 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12797 \$213667 \$213666 \$215494 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12798 \$215494 \$213669 \$215493 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12799 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215493
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12800 \$213669 \$213667 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12801 \$213669 \$213666 \$213670 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12802 \$213670 \$213665 \$215229 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12803 \$213687 cp|i|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12804 VSS|anode|cathode|clk|vss \$213687 \$213688 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12805 VSS|anode|cathode|clk|vss \$213687 \$215489 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12806 \$215489 d|z$40 \$213689 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12807 \$213689 \$213688 \$215490 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12808 \$215490 \$213691 \$215491 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12809 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215491
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12810 \$213691 \$213689 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12811 \$213691 \$213688 \$213692 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12812 \$213692 \$213687 \$215230 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12813 \$213701 cp|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12814 VSS|anode|cathode|clk|vss \$213701 \$213702 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12815 VSS|anode|cathode|clk|vss \$213701 \$215475 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12816 \$215475 d|z$37 \$213703 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12817 \$213703 \$213702 \$215476 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12818 \$215476 \$213705 \$215477 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12819 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215477
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12820 \$213705 \$213703 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12821 \$213705 \$213702 \$213706 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12822 \$213706 \$213701 \$215231 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12823 \$213714 cp|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12824 VSS|anode|cathode|clk|vss \$213714 \$213715 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12825 VSS|anode|cathode|clk|vss \$213714 \$215464 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12826 \$215464 d|z$43 \$213716 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12827 \$213716 \$213715 \$215467 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12828 \$215467 \$213718 \$215468 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12829 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215468
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12830 \$213718 \$213716 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12831 \$213718 \$213715 \$213719 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12832 \$213719 \$213714 \$215232 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12833 VSS|anode|cathode|clk|vss cp|i|z$2 \$215799 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12834 VSS|anode|cathode|clk|vss \$215799 \$215504 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12835 \$215800 \$215504 \$215881 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12836 \$215881 \$215801 \$215879 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12837 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215879
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12838 \$215505 \$215799 \$215802 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12839 VSS|anode|cathode|clk|vss \$215799 \$215882 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12840 \$215882 d|z$50 \$215800 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12841 VSS|anode|cathode|clk|vss \$215800 \$215801 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12842 \$215801 \$215504 \$215505 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12843 VSS|anode|cathode|clk|vss \$215803 \$215802 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12844 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215933
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12845 \$215933 \$215505 \$215803 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12846 VSS|anode|cathode|clk|vss \$215803 a1|a2|q$6 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12847 VSS|anode|cathode|clk|vss a2|q$4 \$215932 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12848 \$215932 a1|b|d|z \$215804 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12849 VSS|anode|cathode|clk|vss \$215804 d|z$29 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12850 VSS|anode|cathode|clk|vss a1|a2|q$6 a3|zn$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12851 a3|zn$1 a2|q$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12852 VSS|anode|cathode|clk|vss a1|a2|q a4|zn$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12853 a4|zn$1 a2|q$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12854 z$31 cp|i|z$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12855 VSS|anode|cathode|clk|vss cp|i|z$2 \$215806 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12856 VSS|anode|cathode|clk|vss \$215806 \$215506 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12857 \$215807 \$215506 \$215891 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12858 \$215891 \$215808 \$215898 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12859 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215898
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12860 \$215507 \$215806 \$215809 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12861 VSS|anode|cathode|clk|vss \$215806 \$215892 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12862 \$215892 a1|b|d|z \$215807 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12863 VSS|anode|cathode|clk|vss \$215807 \$215808 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12864 \$215808 \$215506 \$215507 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12865 VSS|anode|cathode|clk|vss \$215810 \$215809 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12866 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215934
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12867 \$215934 \$215507 \$215810 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12868 VSS|anode|cathode|clk|vss \$215810 a1|a2|q$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12869 VSS|anode|cathode|clk|vss a2|i|q$2 \$215936 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12870 \$215936 a1|b|d|z \$215812 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12871 VSS|anode|cathode|clk|vss \$215812 d|s|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12872 \$215814 d|s|zn \$215815 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12873 \$215816 \$215509 \$215814 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12874 VSS|anode|cathode|clk|vss a1|i0|q$1 \$215816 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12875 VSS|anode|cathode|clk|vss DATA|core|i0|i1|p2c \$215815
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p
+ AD=0.244125p PS=2.27u PD=1.53u
M$12876 VSS|anode|cathode|clk|vss d|s|zn \$215509 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12877 VSS|anode|cathode|clk|vss \$215814 d|z$44 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12878 VSS|anode|cathode|clk|vss a2|zn$9 \$215943 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12879 \$215943 a1|i0|q a2|i|s|zn VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12880 \$215819 s|zn$1 \$215820 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12881 \$215821 \$215510 \$215819 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12882 VSS|anode|cathode|clk|vss i0|i1|q$4 \$215821 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12883 VSS|anode|cathode|clk|vss a1|i|i0|i1|q \$215820
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p
+ AD=0.244125p PS=2.27u PD=1.53u
M$12884 VSS|anode|cathode|clk|vss s|zn$1 \$215510 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12885 VSS|anode|cathode|clk|vss \$215819 d|z$42 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12886 VSS|anode|cathode|clk|vss cp|i|z$3 \$215822 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12887 VSS|anode|cathode|clk|vss \$215822 \$215511 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12888 \$215823 \$215511 \$215899 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12889 \$215899 \$215824 \$215900 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12890 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215900
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12891 \$215512 \$215822 \$215825 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12892 VSS|anode|cathode|clk|vss \$215822 \$215897 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12893 \$215897 d|z$46 \$215823 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12894 VSS|anode|cathode|clk|vss \$215823 \$215824 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12895 \$215824 \$215511 \$215512 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12896 VSS|anode|cathode|clk|vss \$215826 \$215825 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12897 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215944
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12898 \$215944 \$215512 \$215826 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12899 VSS|anode|cathode|clk|vss \$215826 a2|i|i0|i1|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$12900 VSS|anode|cathode|clk|vss a1|a2|q$2 a1|zn VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12901 a1|zn a2|q$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12902 VSS|anode|cathode|clk|vss cp|i|z$3 \$215828 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12903 VSS|anode|cathode|clk|vss \$215828 \$215513 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12904 \$215829 \$215513 \$215895 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12905 \$215895 \$215830 \$215896 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12906 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215896
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12907 \$215514 \$215828 \$215831 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12908 VSS|anode|cathode|clk|vss \$215828 \$215894 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12909 \$215894 d|z$47 \$215829 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12910 VSS|anode|cathode|clk|vss \$215829 \$215830 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12911 \$215830 \$215513 \$215514 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12912 VSS|anode|cathode|clk|vss \$215832 \$215831 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12913 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215947
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12914 \$215947 \$215514 \$215832 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12915 VSS|anode|cathode|clk|vss \$215832 R[18]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12916 VSS|anode|cathode|clk|vss cp|i|z$4 \$215834 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12917 VSS|anode|cathode|clk|vss \$215834 \$215515 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12918 \$215835 \$215515 \$215889 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12919 \$215889 \$215836 \$215890 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12920 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215890
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12921 \$215516 \$215834 \$215837 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12922 VSS|anode|cathode|clk|vss \$215834 \$215893 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12923 \$215893 d|z$36 \$215835 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12924 VSS|anode|cathode|clk|vss \$215835 \$215836 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12925 \$215836 \$215515 \$215516 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12926 VSS|anode|cathode|clk|vss \$215838 \$215837 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12927 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215949
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12928 \$215949 \$215516 \$215838 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12929 VSS|anode|cathode|clk|vss \$215838 R[39]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12930 VSS|anode|cathode|clk|vss cp|i|z$4 \$215839 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12931 VSS|anode|cathode|clk|vss \$215839 \$215517 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12932 \$215840 \$215517 \$215887 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12933 \$215887 \$215841 \$215888 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12934 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215888
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12935 \$215518 \$215839 \$215842 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12936 VSS|anode|cathode|clk|vss \$215839 \$215886 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12937 \$215886 d|z$48 \$215840 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12938 VSS|anode|cathode|clk|vss \$215840 \$215841 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12939 \$215841 \$215517 \$215518 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12940 VSS|anode|cathode|clk|vss \$215843 \$215842 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12941 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215951
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12942 \$215951 \$215518 \$215843 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12943 VSS|anode|cathode|clk|vss \$215843 R[23]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12944 \$215845 s|zn$2 \$215846 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12945 \$215847 \$215519 \$215845 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12946 VSS|anode|cathode|clk|vss R[22]|i0|q \$215847 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12947 VSS|anode|cathode|clk|vss i0|i1|q$3 \$215846 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12948 VSS|anode|cathode|clk|vss s|zn$2 \$215519 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12949 VSS|anode|cathode|clk|vss \$215845 d|z$45 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12950 VSS|anode|cathode|clk|vss cp|i|z$1 \$215849 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12951 VSS|anode|cathode|clk|vss \$215849 \$215520 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12952 \$215850 \$215520 \$215884 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12953 \$215884 \$215851 \$215885 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12954 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215885
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12955 \$215521 \$215849 \$215852 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12956 VSS|anode|cathode|clk|vss \$215849 \$215883 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12957 \$215883 d|z$45 \$215850 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12958 VSS|anode|cathode|clk|vss \$215850 \$215851 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12959 \$215851 \$215520 \$215521 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12960 VSS|anode|cathode|clk|vss \$215853 \$215852 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12961 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215950
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12962 \$215950 \$215521 \$215853 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12963 VSS|anode|cathode|clk|vss \$215853 R[22]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12964 \$215854 s|zn \$215855 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12965 \$215856 \$215522 \$215854 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12966 VSS|anode|cathode|clk|vss i0|i1|q$1 \$215856 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12967 VSS|anode|cathode|clk|vss R[35]|i1|q \$215855 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12968 VSS|anode|cathode|clk|vss s|zn \$215522 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12969 VSS|anode|cathode|clk|vss \$215854 d|z$49 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12970 VSS|anode|cathode|clk|vss cp|z$4 \$215857 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12971 VSS|anode|cathode|clk|vss \$215857 \$215523 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12972 \$215858 \$215523 \$215878 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12973 \$215878 \$215859 \$215880 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12974 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215880
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12975 \$215524 \$215857 \$215860 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12976 VSS|anode|cathode|clk|vss \$215857 \$215877 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12977 \$215877 d|z$49 \$215858 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12978 VSS|anode|cathode|clk|vss \$215858 \$215859 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12979 \$215859 \$215523 \$215524 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12980 VSS|anode|cathode|clk|vss \$215861 \$215860 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12981 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215946
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$12982 \$215946 \$215524 \$215861 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12983 VSS|anode|cathode|clk|vss \$215861 R[35]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12984 \$215862 s|zn$1 \$215863 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12985 \$215864 \$215525 \$215862 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12986 VSS|anode|cathode|clk|vss i0|i1|q$7 \$215864 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12987 VSS|anode|cathode|clk|vss i0|i1|q$3 \$215863 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12988 VSS|anode|cathode|clk|vss s|zn$1 \$215525 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12989 VSS|anode|cathode|clk|vss \$215862 d|z$35 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12990 \$215865 s|zn$1 \$215866 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12991 \$215867 \$215526 \$215865 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12992 VSS|anode|cathode|clk|vss i0|i1|q$3 \$215867 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12993 VSS|anode|cathode|clk|vss i0|i1|q$4 \$215866 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12994 VSS|anode|cathode|clk|vss s|zn$1 \$215526 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12995 VSS|anode|cathode|clk|vss \$215865 d|z$43 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12996 VSS|anode|cathode|clk|vss cp|z$4 \$215868 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12997 VSS|anode|cathode|clk|vss \$215868 \$215527 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12998 \$215869 \$215527 \$215875 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12999 \$215875 \$215870 \$215876 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13000 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215876
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13001 \$215528 \$215868 \$215871 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13002 VSS|anode|cathode|clk|vss \$215868 \$215874 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13003 \$215874 d|z$51 \$215869 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13004 VSS|anode|cathode|clk|vss \$215869 \$215870 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13005 \$215870 \$215527 \$215528 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13006 VSS|anode|cathode|clk|vss \$215872 \$215871 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13007 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$215941
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13008 \$215941 \$215528 \$215872 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13009 VSS|anode|cathode|clk|vss \$215872 R[53]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13010 d|z$50 \$217719 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13011 VSS|anode|cathode|clk|vss \$218627 \$218784 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13012 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219548
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13013 \$219548 \$217723 \$218627 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13014 VSS|anode|cathode|clk|vss \$218627 a1|a2|q$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13015 d|z$52 \$217725 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13016 a2|z$8 a2|i|q$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$13017 \$218785 a3|zn$2 \$219551 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13018 \$219551 a2|z$8 \$219550 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$13019 \$219550 a1|a2|q$7 a1|zn$1 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13020 \$218785 a4|zn$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13021 VSS|anode|cathode|clk|vss \$218628 \$218786 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13022 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219561
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13023 \$219561 \$217732 \$218628 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13024 VSS|anode|cathode|clk|vss \$218628 a2|i|q$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13025 VSS|anode|cathode|clk|vss \$218629 \$218787 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13026 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219567
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13027 \$219567 \$217736 \$218629 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13028 VSS|anode|cathode|clk|vss \$218629 a1|i0|q$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13029 VSS|anode|cathode|clk|vss \$218630 \$218788 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13030 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219568
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13031 \$219568 \$217740 \$218630 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13032 VSS|anode|cathode|clk|vss \$218630 a1|a3|i|i1|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13033 VSS|anode|cathode|clk|vss \$218631 \$218789 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13034 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219578
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13035 \$219578 \$217746 \$218631 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13036 VSS|anode|cathode|clk|vss \$218631 R[50]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13037 \$217748 s|zn$2 \$217747 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13038 \$217748 i0|i1|q$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13039 VSS|anode|cathode|clk|vss R[18]|i0|q \$217749 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13040 \$217749 \$217666 \$217747 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13041 VSS|anode|cathode|clk|vss s|zn$2 \$217666 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13042 VSS|anode|cathode|clk|vss \$217747 d|z$47 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13043 \$217751 s|zn$2 \$217750 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13044 \$217751 i0|i1|q$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13045 VSS|anode|cathode|clk|vss R[21]|i0|q \$217752 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13046 \$217752 \$217668 \$217750 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13047 VSS|anode|cathode|clk|vss s|zn$2 \$217668 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13048 VSS|anode|cathode|clk|vss \$217750 d|z$39 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13049 VSS|anode|cathode|clk|vss \$218632 \$218790 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13050 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219598
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13051 \$219598 \$217756 \$218632 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13052 VSS|anode|cathode|clk|vss \$218632 R[31]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13053 VSS|anode|cathode|clk|vss \$218633 \$218791 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13054 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219607
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13055 \$219607 \$217761 \$218633 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13056 VSS|anode|cathode|clk|vss \$218633 R[17]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13057 VSS|anode|cathode|clk|vss \$218634 \$218792 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13058 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219613
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13059 \$219613 \$217766 \$218634 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13060 VSS|anode|cathode|clk|vss \$218634 R[19]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13061 \$217769 s|zn$2 \$217768 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13062 \$217769 i0|i1|q$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13063 VSS|anode|cathode|clk|vss R[20]|i0|q \$217770 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13064 \$217770 \$217672 \$217768 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13065 VSS|anode|cathode|clk|vss s|zn$2 \$217672 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13066 VSS|anode|cathode|clk|vss \$217768 d|z$40 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13067 VSS|anode|cathode|clk|vss \$218635 \$218793 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13068 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219606
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13069 \$219606 \$217774 \$218635 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13070 VSS|anode|cathode|clk|vss \$218635 R[38]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13071 \$217777 s|zn$3 \$217776 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13072 \$217777 R[51]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13073 VSS|anode|cathode|clk|vss i0|i1|q$1 \$217778 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13074 \$217778 \$217674 \$217776 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13075 VSS|anode|cathode|clk|vss s|zn$3 \$217674 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13076 VSS|anode|cathode|clk|vss \$217776 d|z$53 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13077 \$217781 s|zn$3 \$217780 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13078 \$217781 R[49]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13079 VSS|anode|cathode|clk|vss i0|i1|q$6 \$217782 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13080 \$217782 \$217676 \$217780 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13081 VSS|anode|cathode|clk|vss s|zn$3 \$217676 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13082 VSS|anode|cathode|clk|vss \$217780 d|z$54 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13083 VSS|anode|cathode|clk|vss \$218636 \$218794 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13084 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219590
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13085 \$219590 \$217787 \$218636 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13086 VSS|anode|cathode|clk|vss \$218636 R[49]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13087 VSS|anode|cathode|clk|vss a1|a2|b|q|s \$219540
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p
+ AD=0.263525p PS=3.88u PD=1.465u
M$13088 \$219540 a1|b|d|z \$217719 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13089 \$217661 cp|i|z$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13090 VSS|anode|cathode|clk|vss \$217661 \$217720 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13091 VSS|anode|cathode|clk|vss \$217661 \$219545 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13092 \$219545 d|s|z \$217721 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13093 \$217721 \$217720 \$219544 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13094 \$219544 \$218407 \$219543 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13095 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219543
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13096 \$218407 \$217721 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13097 \$218407 \$217720 \$217723 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13098 \$217723 \$217661 \$218784 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13099 VSS|anode|cathode|clk|vss a2|q$7 \$219547 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13100 \$219547 a1|b|d|z \$217725 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13101 \$217662 cp|i|z$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13102 VSS|anode|cathode|clk|vss \$217662 \$217729 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13103 VSS|anode|cathode|clk|vss \$217662 \$219559 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13104 \$219559 d|s|zn \$217730 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13105 \$217730 \$217729 \$219555 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13106 \$219555 \$218408 \$219554 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13107 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219554
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13108 \$218408 \$217730 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13109 \$218408 \$217729 \$217732 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13110 \$217732 \$217662 \$218786 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13111 \$217663 cp|i|z$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13112 VSS|anode|cathode|clk|vss \$217663 \$217733 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13113 VSS|anode|cathode|clk|vss \$217663 \$219565 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13114 \$219565 d|z$44 \$217734 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13115 \$217734 \$217733 \$219564 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13116 \$219564 \$218409 \$219563 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13117 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219563
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13118 \$218409 \$217734 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13119 \$218409 \$217733 \$217736 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13120 \$217736 \$217663 \$218787 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13121 \$217664 cp|i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13122 VSS|anode|cathode|clk|vss \$217664 \$217737 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13123 VSS|anode|cathode|clk|vss \$217664 \$219566 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13124 \$219566 d|z$55 \$217738 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13125 \$217738 \$217737 \$219570 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13126 \$219570 \$218410 \$219569 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13127 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219569
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13128 \$218410 \$217738 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13129 \$218410 \$217737 \$217740 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13130 \$217740 \$217664 \$218788 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13131 \$217665 cp|i|z$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13132 VSS|anode|cathode|clk|vss \$217665 \$217742 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13133 VSS|anode|cathode|clk|vss \$217665 \$219572 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13134 \$219572 d|z$56 \$217743 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13135 \$217743 \$217742 \$219571 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13136 \$219571 \$218411 \$219581 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13137 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219581
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13138 \$218411 \$217743 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13139 \$218411 \$217742 \$217746 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13140 \$217746 \$217665 \$218789 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13141 \$217669 cp|i|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13142 VSS|anode|cathode|clk|vss \$217669 \$217753 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13143 VSS|anode|cathode|clk|vss \$217669 \$219594 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13144 \$219594 d|z$57 \$217754 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13145 \$217754 \$217753 \$219592 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13146 \$219592 \$218412 \$219591 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13147 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219591
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13148 \$218412 \$217754 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13149 \$218412 \$217753 \$217756 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13150 \$217756 \$217669 \$218790 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13151 \$217670 cp|i|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13152 VSS|anode|cathode|clk|vss \$217670 \$217758 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13153 VSS|anode|cathode|clk|vss \$217670 \$219602 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13154 \$219602 d|z$58 \$217759 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13155 \$217759 \$217758 \$219601 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13156 \$219601 \$218413 \$219600 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13157 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219600
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13158 \$218413 \$217759 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13159 \$218413 \$217758 \$217761 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13160 \$217761 \$217670 \$218791 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13161 \$217671 cp|i|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13162 VSS|anode|cathode|clk|vss \$217671 \$217763 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13163 VSS|anode|cathode|clk|vss \$217671 \$219611 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13164 \$219611 d|z$59 \$217764 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13165 \$217764 \$217763 \$219610 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13166 \$219610 \$218414 \$219609 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13167 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219609
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13168 \$218414 \$217764 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13169 \$218414 \$217763 \$217766 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13170 \$217766 \$217671 \$218792 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13171 \$217673 cp|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13172 VSS|anode|cathode|clk|vss \$217673 \$217771 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13173 VSS|anode|cathode|clk|vss \$217673 \$219612 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13174 \$219612 d|z$60 \$217772 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13175 \$217772 \$217771 \$219604 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13176 \$219604 \$218415 \$219603 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13177 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219603
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13178 \$218415 \$217772 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13179 \$218415 \$217771 \$217774 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13180 \$217774 \$217673 \$218793 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13181 \$217677 cp|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13182 VSS|anode|cathode|clk|vss \$217677 \$217784 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13183 VSS|anode|cathode|clk|vss \$217677 \$219595 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13184 \$219595 d|z$54 \$217785 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13185 \$217785 \$217784 \$219596 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13186 \$219596 \$218416 \$219597 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13187 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$219597
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13188 \$218416 \$217785 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13189 \$218416 \$217784 \$217787 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13190 \$217787 \$217677 \$218794 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13191 VSS|anode|cathode|clk|vss cp|i|z$5 \$219901 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13192 VSS|anode|cathode|clk|vss \$219901 \$219614 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13193 \$219902 \$219614 \$220008 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13194 \$220008 \$219903 \$220007 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13195 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220007
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13196 \$219615 \$219901 \$219904 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13197 VSS|anode|cathode|clk|vss \$219901 \$220009 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13198 \$220009 d|z$63 \$219902 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13199 VSS|anode|cathode|clk|vss \$219902 \$219903 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13200 \$219903 \$219614 \$219615 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13201 VSS|anode|cathode|clk|vss \$219905 \$219904 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13202 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220338
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13203 \$220338 \$219615 \$219905 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13204 VSS|anode|cathode|clk|vss \$219905 a2|q$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13205 VSS|anode|cathode|clk|vss cp|i|z$5 \$219906 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13206 VSS|anode|cathode|clk|vss \$219906 \$219616 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13207 \$219907 \$219616 \$220015 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13208 \$220015 \$219908 \$220019 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13209 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220019
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13210 \$219617 \$219906 \$219909 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13211 VSS|anode|cathode|clk|vss \$219906 \$220016 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13212 \$220016 d|z$52 \$219907 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13213 VSS|anode|cathode|clk|vss \$219907 \$219908 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13214 \$219908 \$219616 \$219617 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13215 VSS|anode|cathode|clk|vss \$219910 \$219909 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13216 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220339
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13217 \$220339 \$219617 \$219910 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13218 VSS|anode|cathode|clk|vss \$219910 a1|a2|q$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13219 VSS|anode|cathode|clk|vss cp|i|z$5 \$219912 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13220 VSS|anode|cathode|clk|vss \$219912 \$219618 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13221 \$219913 \$219618 \$220020 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13222 \$220020 \$219914 \$220025 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13223 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220025
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13224 \$219619 \$219912 \$219915 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13225 VSS|anode|cathode|clk|vss \$219912 \$220021 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13226 \$220021 d|z$64 \$219913 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13227 VSS|anode|cathode|clk|vss \$219913 \$219914 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13228 \$219914 \$219618 \$219619 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13229 VSS|anode|cathode|clk|vss \$219916 \$219915 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13230 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220342
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13231 \$220342 \$219619 \$219916 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13232 VSS|anode|cathode|clk|vss \$219916 a1|a2|b|q|s
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13233 \$219918 d|s|z \$219919 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13234 \$219920 \$219620 \$219918 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13235 VSS|anode|cathode|clk|vss a1|i0|q \$219920 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13236 VSS|anode|cathode|clk|vss DATA|core|i0|i1|p2c \$219919
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p
+ AD=0.244125p PS=2.27u PD=1.53u
M$13237 VSS|anode|cathode|clk|vss d|s|z \$219620 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13238 VSS|anode|cathode|clk|vss \$219918 d|z$41 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13239 VSS|anode|cathode|clk|vss a1|a2|q$5 \$220027 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13240 \$220027 a1|i0|q$1 \$219921 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13241 VSS|anode|cathode|clk|vss \$219921 a1|a2|a4|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13242 \$219922 s|zn$1 \$219923 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13243 \$219924 \$219621 \$219922 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13244 VSS|anode|cathode|clk|vss a1|i|i0|i1|q \$219924
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13245 VSS|anode|cathode|clk|vss a2|i|i0|i1|q \$219923
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p
+ AD=0.244125p PS=2.27u PD=1.53u
M$13246 VSS|anode|cathode|clk|vss s|zn$1 \$219621 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13247 VSS|anode|cathode|clk|vss \$219922 d|z$46 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13248 \$219925 s|zn$1 \$219926 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13249 \$219927 \$219622 \$219925 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13250 VSS|anode|cathode|clk|vss a2|i|i0|i1|q \$219927
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13251 VSS|anode|cathode|clk|vss a1|a3|i|i1|q \$219926
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p
+ AD=0.244125p PS=2.27u PD=1.53u
M$13252 VSS|anode|cathode|clk|vss s|zn$1 \$219622 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13253 VSS|anode|cathode|clk|vss \$219925 d|z$55 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13254 VSS|anode|cathode|clk|vss a1|zn$2 s|zn$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13255 s|zn$4 a2|zn$11 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13256 VSS|anode|cathode|clk|vss a1|i|i0|i1|q a2|a3|zn$1
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p
+ PS=2.53u PD=1.53u
M$13257 a2|a3|zn$1 a2|i|i0|i1|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p
+ PS=1.53u PD=2.53u
M$13258 \$219928 s|zn$3 \$219929 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13259 \$219930 \$219623 \$219928 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13260 VSS|anode|cathode|clk|vss i0|i1|q$2 \$219930 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13261 VSS|anode|cathode|clk|vss R[50]|i1|q \$219929 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13262 VSS|anode|cathode|clk|vss s|zn$3 \$219623 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13263 VSS|anode|cathode|clk|vss \$219928 d|z$56 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13264 VSS|anode|cathode|clk|vss cp|i|z$6 \$219931 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13265 VSS|anode|cathode|clk|vss \$219931 \$219624 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13266 \$219932 \$219624 \$220132 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13267 \$220132 \$219933 \$220129 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13268 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220129
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13269 \$219625 \$219931 \$219934 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13270 VSS|anode|cathode|clk|vss \$219931 \$220137 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13271 \$220137 d|z$65 \$219932 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13272 VSS|anode|cathode|clk|vss \$219932 \$219933 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13273 \$219933 \$219624 \$219625 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13274 VSS|anode|cathode|clk|vss \$219935 \$219934 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13275 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220373
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13276 \$220373 \$219625 \$219935 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13277 VSS|anode|cathode|clk|vss \$219935 R[54]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13278 \$219626 a1|a2|a4|z \$220355 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13279 \$220355 a1|a3|i|i1|q s|zn VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13280 VSS|anode|cathode|clk|vss a2|a3|zn$1 \$219626 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13281 VSS|anode|cathode|clk|vss a2|z$9 \$220158 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13282 \$220158 a1|a2|a4|z \$219937 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13283 VSS|anode|cathode|clk|vss \$219937 s|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13284 \$219938 s|z \$219939 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13285 \$219940 \$219627 \$219938 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13286 VSS|anode|cathode|clk|vss R[31]|i0|q \$219940 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13287 VSS|anode|cathode|clk|vss i0|i1|q$4 \$219939 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13288 VSS|anode|cathode|clk|vss s|z \$219627 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13289 VSS|anode|cathode|clk|vss \$219938 d|z$57 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13290 \$219941 s|zn$3 \$219942 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13291 \$219943 \$219628 \$219941 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13292 VSS|anode|cathode|clk|vss i0|i1|q$5 \$219943 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13293 VSS|anode|cathode|clk|vss R[52]|i1|q \$219942 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13294 VSS|anode|cathode|clk|vss s|zn$3 \$219628 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13295 VSS|anode|cathode|clk|vss \$219941 d|z$61 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13296 \$219945 s|zn$2 \$219946 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13297 \$219947 \$219629 \$219945 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13298 VSS|anode|cathode|clk|vss R[23]|i0|q \$219947 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13299 VSS|anode|cathode|clk|vss i0|i1|q$4 \$219946 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13300 VSS|anode|cathode|clk|vss s|zn$2 \$219629 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13301 VSS|anode|cathode|clk|vss \$219945 d|z$48 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13302 \$219948 s|zn$2 \$219949 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13303 \$219950 \$219630 \$219948 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13304 VSS|anode|cathode|clk|vss R[17]|i0|q \$219950 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13305 VSS|anode|cathode|clk|vss i0|i1|q$6 \$219949 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13306 VSS|anode|cathode|clk|vss s|zn$2 \$219630 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13307 VSS|anode|cathode|clk|vss \$219948 d|z$58 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13308 \$219951 s|zn$2 \$219952 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13309 \$219953 \$219631 \$219951 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13310 VSS|anode|cathode|clk|vss R[16]|i0|q \$219953 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13311 VSS|anode|cathode|clk|vss i0|i1|q \$219952 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13312 VSS|anode|cathode|clk|vss s|zn$2 \$219631 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13313 VSS|anode|cathode|clk|vss \$219951 d|z$62 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13314 VSS|anode|cathode|clk|vss cp|i|z$7 \$219955 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13315 VSS|anode|cathode|clk|vss \$219955 \$219632 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13316 \$219956 \$219632 \$220189 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13317 \$220189 \$219957 \$220191 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13318 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220191
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13319 \$219633 \$219955 \$219958 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13320 VSS|anode|cathode|clk|vss \$219955 \$220188 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13321 \$220188 d|z$62 \$219956 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13322 VSS|anode|cathode|clk|vss \$219956 \$219957 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13323 \$219957 \$219632 \$219633 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13324 VSS|anode|cathode|clk|vss \$219959 \$219958 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13325 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220388
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13326 \$220388 \$219633 \$219959 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13327 VSS|anode|cathode|clk|vss \$219959 R[16]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13328 \$219960 s|zn \$219961 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13329 \$219962 \$219634 \$219960 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13330 VSS|anode|cathode|clk|vss i0|i1|q$3 \$219962 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13331 VSS|anode|cathode|clk|vss R[38]|i1|q \$219961 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13332 VSS|anode|cathode|clk|vss s|zn \$219634 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13333 VSS|anode|cathode|clk|vss \$219960 d|z$60 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13334 VSS|anode|cathode|clk|vss cp|z$4 \$219963 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13335 VSS|anode|cathode|clk|vss \$219963 \$219635 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13336 \$219964 \$219635 \$220179 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13337 \$220179 \$219965 \$220180 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13338 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220180
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13339 \$219636 \$219963 \$219966 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13340 VSS|anode|cathode|clk|vss \$219963 \$220178 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13341 \$220178 d|z$66 \$219964 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13342 VSS|anode|cathode|clk|vss \$219964 \$219965 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13343 \$219965 \$219635 \$219636 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13344 VSS|anode|cathode|clk|vss \$219967 \$219966 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13345 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220386
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13346 \$220386 \$219636 \$219967 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13347 VSS|anode|cathode|clk|vss \$219967 R[48]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13348 VSS|anode|cathode|clk|vss cp|z$4 \$219969 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13349 VSS|anode|cathode|clk|vss \$219969 \$219637 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13350 \$219970 \$219637 \$220172 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13351 \$220172 \$219971 \$220173 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13352 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220173
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13353 \$219638 \$219969 \$219972 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13354 VSS|anode|cathode|clk|vss \$219969 \$220171 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13355 \$220171 d|z$53 \$219970 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13356 VSS|anode|cathode|clk|vss \$219970 \$219971 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13357 \$219971 \$219637 \$219638 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13358 VSS|anode|cathode|clk|vss \$219973 \$219972 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13359 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220385
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13360 \$220385 \$219638 \$219973 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13361 VSS|anode|cathode|clk|vss \$219973 R[51]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13362 VSS|anode|cathode|clk|vss cp|z$4 \$219974 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13363 VSS|anode|cathode|clk|vss \$219974 \$219639 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13364 \$219975 \$219639 \$220165 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13365 \$220165 \$219976 \$220166 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13366 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220166
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13367 \$219640 \$219974 \$219977 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13368 VSS|anode|cathode|clk|vss \$219974 \$220163 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13369 \$220163 d|z$67 \$219975 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13370 VSS|anode|cathode|clk|vss \$219975 \$219976 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13371 \$219976 \$219639 \$219640 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13372 VSS|anode|cathode|clk|vss \$219978 \$219977 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13373 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$220382
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13374 \$220382 \$219640 \$219978 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13375 VSS|anode|cathode|clk|vss \$219978 R[55]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13376 \$219980 s|zn$3 \$219981 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13377 \$219982 \$219641 \$219980 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13378 VSS|anode|cathode|clk|vss i0|i1|q$7 \$219982 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13379 VSS|anode|cathode|clk|vss R[53]|i1|q \$219981 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13380 VSS|anode|cathode|clk|vss s|zn$3 \$219641 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13381 VSS|anode|cathode|clk|vss \$219980 d|z$51 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13382 VSS|anode|cathode|clk|vss a1|a2|q$8 \$223800 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13383 \$223800 a1|b|d|z \$222044 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13384 d|z$63 \$222044 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13385 VSS|anode|cathode|clk|vss a1|a2|q$8 a3|zn$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13386 a3|zn$2 a2|q$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13387 VSS|anode|cathode|clk|vss a1|a2|q$9 \$223801 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13388 \$223801 a1|b|d|z \$222046 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13389 d|z$64 \$222046 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13390 \$222047 a1|a2|b|q|s \$222022 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13391 \$222047 i1|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13392 VSS|anode|cathode|clk|vss i0|z \$222048 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13393 \$222048 \$221966 \$222022 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13394 VSS|anode|cathode|clk|vss a1|a2|b|q|s \$221966
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$13395 VSS|anode|cathode|clk|vss \$222022 d|z$68 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13396 VSS|anode|cathode|clk|vss a1|a2|q$9 a4|zn$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13397 a4|zn$2 a1|a2|b|q|s VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13398 VSS|anode|cathode|clk|vss CEB|a1|core|i|p2c d|s|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p
+ PS=2.53u PD=1.53u
M$13399 d|s|zn a1|a2|q$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13400 a1|b|d|z CEB|a1|core|i|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$13401 VSS|anode|cathode|clk|vss a1|a2|q$5 \$223799 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13402 \$223799 a1|i0|q$1 a1|zn$2 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13403 \$222051 s|z$1 \$222023 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13404 \$222051 i0|i1|q$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13405 VSS|anode|cathode|clk|vss R[7]|i|i0|q \$222052
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13406 \$222052 \$221967 \$222023 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13407 VSS|anode|cathode|clk|vss s|z$1 \$221967 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13408 VSS|anode|cathode|clk|vss \$222023 d|z$69 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13409 cp|i|z$6 \$222024 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$13410 VSS|anode|cathode|clk|vss i|z$115 \$222024 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13411 \$222054 s|zn$4 \$222025 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13412 \$222054 i0|i1|q$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13413 VSS|anode|cathode|clk|vss R[47]|i0|q \$222055 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13414 \$222055 \$221969 \$222025 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13415 VSS|anode|cathode|clk|vss s|zn$4 \$221969 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13416 VSS|anode|cathode|clk|vss \$222025 d|z$70 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13417 z$32 cp|i|z$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$13418 VSS|anode|cathode|clk|vss a1|zn$14 \$222058 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13419 \$222058 a2|zn$32 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.263525p AD=0.374525p PS=1.465u PD=2.205u
M$13420 VSS|anode|cathode|clk|vss \$222058 i1|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.374525p AD=0.358775p PS=2.205u PD=2.4u
M$13421 \$223078 a2|i|i0|i1|q \$223798 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13422 \$223798 a1|z$15 a2|zn$12 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13423 \$223078 a1|a3|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13424 VSS|anode|cathode|clk|vss a1|zn$2 s|zn$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13425 s|zn$2 a2|zn$12 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13426 \$222061 s|zn$3 \$222026 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13427 \$222061 R[54]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13428 VSS|anode|cathode|clk|vss i0|i1|q$3 \$222062 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13429 \$222062 \$221971 \$222026 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13430 VSS|anode|cathode|clk|vss s|zn$3 \$221971 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13431 VSS|anode|cathode|clk|vss \$222026 d|z$65 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13432 \$223079 a1|a3|i|i1|q \$223796 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13433 \$223796 a2|i|i0|i1|q \$223795 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$13434 \$223795 a1|z$15 s|zn$3 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13435 \$223079 a1|a2|a4|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13436 VSS|anode|cathode|clk|vss a2|a3|z$1 \$223797 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13437 \$223797 a1|a3|z \$222063 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13438 a2|z$9 \$222063 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13439 i|z$115 \$222027 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$13440 VSS|anode|cathode|clk|vss CLK|core|i|p2c$1 \$222027
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$13441 VSS|anode|cathode|clk|vss \$222738 \$223080 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13442 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$223794
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13443 \$223794 \$222031 \$222738 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13444 VSS|anode|cathode|clk|vss \$222738 R[52]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13445 \$222065 s|zn$5 \$222032 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13446 \$222065 i0|i1|q$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13447 VSS|anode|cathode|clk|vss R[15]|i|i0|q \$222066
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13448 \$222066 \$221972 \$222032 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13449 VSS|anode|cathode|clk|vss s|zn$5 \$221972 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13450 VSS|anode|cathode|clk|vss \$222032 d|z$71 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13451 \$222068 s|zn$2 \$222033 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13452 \$222068 i0|i1|q$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13453 VSS|anode|cathode|clk|vss R[19]|i0|q \$222069 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13454 \$222069 \$221974 \$222033 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13455 VSS|anode|cathode|clk|vss s|zn$2 \$221974 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13456 VSS|anode|cathode|clk|vss \$222033 d|z$59 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13457 \$222070 s|zn$5 \$222034 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13458 \$222070 i0|i1|q$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13459 VSS|anode|cathode|clk|vss R[12]|i|i0|q \$222071
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13460 \$222071 \$221975 \$222034 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13461 VSS|anode|cathode|clk|vss s|zn$5 \$221975 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13462 VSS|anode|cathode|clk|vss \$222034 d|z$72 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13463 \$222073 s|z$1 \$222035 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13464 \$222073 i0|i1|q$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13465 VSS|anode|cathode|clk|vss R[4]|i|i0|q \$222074
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13466 \$222074 \$221976 \$222035 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13467 VSS|anode|cathode|clk|vss s|z$1 \$221976 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13468 VSS|anode|cathode|clk|vss \$222035 d|z$73 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13469 \$222076 s|zn$3 \$222036 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13470 \$222076 R[48]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13471 VSS|anode|cathode|clk|vss i0|i1|q \$222077 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13472 \$222077 \$221977 \$222036 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13473 VSS|anode|cathode|clk|vss s|zn$3 \$221977 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13474 VSS|anode|cathode|clk|vss \$222036 d|z$66 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13475 \$222078 s|zn$4 \$222037 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13476 \$222078 i0|i1|q$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13477 VSS|anode|cathode|clk|vss R[44]|i0|q \$222079 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13478 \$222079 \$221978 \$222037 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13479 VSS|anode|cathode|clk|vss s|zn$4 \$221978 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13480 VSS|anode|cathode|clk|vss \$222037 d|z$74 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13481 \$222081 s|zn$3 \$222038 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13482 \$222081 R[55]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13483 VSS|anode|cathode|clk|vss i0|i1|q$4 \$222082 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13484 \$222082 \$221979 \$222038 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13485 VSS|anode|cathode|clk|vss s|zn$3 \$221979 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13486 VSS|anode|cathode|clk|vss \$222038 d|z$67 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13487 \$222083 s|zn$6 \$222039 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13488 \$222083 R[63]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13489 VSS|anode|cathode|clk|vss i0|i1|q$4 \$222084 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13490 \$222084 \$221980 \$222039 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13491 VSS|anode|cathode|clk|vss s|zn$6 \$221980 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13492 VSS|anode|cathode|clk|vss \$222039 d|z$75 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13493 VSS|anode|cathode|clk|vss \$222739 \$223081 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13494 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$223790
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13495 \$223790 \$222043 \$222739 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13496 VSS|anode|cathode|clk|vss \$222739 R[63]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13497 \$222028 cp|i|z$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13498 VSS|anode|cathode|clk|vss \$222028 \$222029 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13499 VSS|anode|cathode|clk|vss \$222028 \$223791 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13500 \$223791 d|z$61 \$222064 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13501 \$222064 \$222029 \$223792 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13502 \$223792 \$222726 \$223793 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13503 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$223793
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13504 \$222726 \$222064 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13505 \$222726 \$222029 \$222031 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13506 \$222031 \$222028 \$223080 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13507 \$222040 cp|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13508 VSS|anode|cathode|clk|vss \$222040 \$222041 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13509 VSS|anode|cathode|clk|vss \$222040 \$223787 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13510 \$223787 d|z$75 \$222086 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13511 \$222086 \$222041 \$223788 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13512 \$223788 \$222729 \$223789 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13513 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$223789
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13514 \$222729 \$222086 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13515 \$222729 \$222041 \$222043 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13516 \$222043 \$222040 \$223081 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13517 \$223948 a2|i|s|zn \$223949 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13518 \$223951 \$223834 \$223948 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13519 VSS|anode|cathode|clk|vss i0|i1|q$8 \$223951 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13520 VSS|anode|cathode|clk|vss i0|i1|q$9 \$223949 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13521 VSS|anode|cathode|clk|vss a2|i|s|zn \$223834 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13522 VSS|anode|cathode|clk|vss \$223948 i0|z$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13523 \$223953 a1|a2|b|q|s \$223954 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13524 \$223956 \$223835 \$223953 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13525 VSS|anode|cathode|clk|vss i0|z$1 \$223956 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13526 VSS|anode|cathode|clk|vss i1|z$1 \$223954 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13527 VSS|anode|cathode|clk|vss a1|a2|b|q|s \$223835
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$13528 VSS|anode|cathode|clk|vss \$223953 d|z$76 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13529 z$33 cp|i|z$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$13530 VSS|anode|cathode|clk|vss i|z$115 \$223959 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13531 VSS|anode|cathode|clk|vss \$223959 cp|i|z$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13532 VSS|anode|cathode|clk|vss cp|i|z$5 \$223960 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13533 VSS|anode|cathode|clk|vss \$223960 \$223836 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13534 \$223961 \$223836 \$224024 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13535 \$224024 \$223962 \$224023 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13536 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224023
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13537 \$223837 \$223960 \$223963 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13538 VSS|anode|cathode|clk|vss \$223960 \$224025 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13539 \$224025 a2|d|z \$223961 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13540 VSS|anode|cathode|clk|vss \$223961 \$223962 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13541 \$223962 \$223836 \$223837 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13542 VSS|anode|cathode|clk|vss \$223964 \$223963 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13543 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224233
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13544 \$224233 \$223837 \$223964 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13545 VSS|anode|cathode|clk|vss \$223964 a2|q$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13546 VSS|anode|cathode|clk|vss a2|q$8 \$224237 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13547 \$224237 a1|b|d|z \$223966 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13548 VSS|anode|cathode|clk|vss \$223966 DOUT_EN|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13549 VSS|anode|cathode|clk|vss cp|i|z$6 \$223968 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13550 VSS|anode|cathode|clk|vss \$223968 \$223838 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13551 \$223969 \$223838 \$224027 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13552 \$224027 \$223970 \$224026 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13553 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224026
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13554 \$223839 \$223968 \$223971 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13555 VSS|anode|cathode|clk|vss \$223968 \$224028 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13556 \$224028 d|z$69 \$223969 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13557 VSS|anode|cathode|clk|vss \$223969 \$223970 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13558 \$223970 \$223838 \$223839 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13559 VSS|anode|cathode|clk|vss \$223972 \$223971 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13560 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224241
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13561 \$224241 \$223839 \$223972 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13562 VSS|anode|cathode|clk|vss \$223972 R[7]|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13563 VSS|anode|cathode|clk|vss cp|i|z$6 \$223973 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13564 VSS|anode|cathode|clk|vss \$223973 \$223840 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13565 \$223974 \$223840 \$224036 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13566 \$224036 \$223975 \$224034 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13567 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224034
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13568 \$223841 \$223973 \$223976 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13569 VSS|anode|cathode|clk|vss \$223973 \$224037 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13570 \$224037 d|z$70 \$223974 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13571 VSS|anode|cathode|clk|vss \$223974 \$223975 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13572 \$223975 \$223840 \$223841 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13573 VSS|anode|cathode|clk|vss \$223977 \$223976 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13574 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224244
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13575 \$224244 \$223841 \$223977 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13576 VSS|anode|cathode|clk|vss \$223977 R[47]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13577 a2|z$12 a2|i|i0|i1|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$13578 VSS|anode|cathode|clk|vss a2|z$10 \$224248 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13579 \$224248 a1|a2|a4|z \$223978 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13580 VSS|anode|cathode|clk|vss \$223978 s|z$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13581 VSS|anode|cathode|clk|vss a2|a3|zn$1 \$224246 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13582 \$224246 a1|a3|z \$223979 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13583 VSS|anode|cathode|clk|vss \$223979 a2|z$10 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13584 VSS|anode|cathode|clk|vss a1|zn$2 s|zn$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13585 s|zn$5 a2|zn$13 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13586 a1|a3|z a1|a3|i|i1|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$13587 VSS|anode|cathode|clk|vss cp|i|z$6 \$223980 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13588 VSS|anode|cathode|clk|vss \$223980 \$223842 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13589 \$223982 \$223842 \$224048 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13590 \$224048 \$223983 \$224046 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13591 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224046
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13592 \$223843 \$223980 \$223984 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13593 VSS|anode|cathode|clk|vss \$223980 \$224049 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13594 \$224049 d|z$78 \$223982 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13595 VSS|anode|cathode|clk|vss \$223982 \$223983 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13596 \$223983 \$223842 \$223843 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13597 VSS|anode|cathode|clk|vss \$223985 \$223984 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13598 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224256
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13599 \$224256 \$223843 \$223985 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13600 VSS|anode|cathode|clk|vss \$223985 R[43]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13601 \$223844 a1|a2|a4|z \$224252 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13602 \$224252 a1|a3|i|i1|q s|zn$6 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13603 VSS|anode|cathode|clk|vss a2|a3|z$1 \$223844 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13604 VSS|anode|cathode|clk|vss a2|i|i0|i1|q \$224257
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p
+ AD=0.263525p PS=3.88u PD=1.465u
M$13605 \$224257 a1|i|i0|i1|q \$223986 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13606 VSS|anode|cathode|clk|vss \$223986 a2|a3|z$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13607 VSS|anode|cathode|clk|vss cp|i|z$7 \$223987 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13608 VSS|anode|cathode|clk|vss \$223987 \$223845 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13609 \$223988 \$223845 \$224054 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13610 \$224054 \$223989 \$224055 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13611 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224055
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13612 \$223846 \$223987 \$223990 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13613 VSS|anode|cathode|clk|vss \$223987 \$224053 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13614 \$224053 d|z$79 \$223988 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13615 VSS|anode|cathode|clk|vss \$223988 \$223989 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13616 \$223989 \$223845 \$223846 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13617 VSS|anode|cathode|clk|vss \$223991 \$223990 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13618 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224260
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13619 \$224260 \$223846 \$223991 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13620 VSS|anode|cathode|clk|vss \$223991 R[46]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13621 VSS|anode|cathode|clk|vss cp|i|z$7 \$223993 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13622 VSS|anode|cathode|clk|vss \$223993 \$223847 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13623 \$223994 \$223847 \$224051 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13624 \$224051 \$223995 \$224052 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13625 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224052
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13626 \$223848 \$223993 \$223996 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13627 VSS|anode|cathode|clk|vss \$223993 \$224050 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13628 \$224050 d|z$71 \$223994 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13629 VSS|anode|cathode|clk|vss \$223994 \$223995 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13630 \$223995 \$223847 \$223848 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13631 VSS|anode|cathode|clk|vss \$223997 \$223996 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13632 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224269
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13633 \$224269 \$223848 \$223997 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13634 VSS|anode|cathode|clk|vss \$223997 R[15]|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13635 VSS|anode|cathode|clk|vss cp|i|z$7 \$223998 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13636 VSS|anode|cathode|clk|vss \$223998 \$223849 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13637 \$223999 \$223849 \$224044 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13638 \$224044 \$224000 \$224045 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13639 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224045
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13640 \$223850 \$223998 \$224001 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13641 VSS|anode|cathode|clk|vss \$223998 \$224047 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13642 \$224047 d|z$72 \$223999 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13643 VSS|anode|cathode|clk|vss \$223999 \$224000 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13644 \$224000 \$223849 \$223850 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13645 VSS|anode|cathode|clk|vss \$224002 \$224001 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13646 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224272
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13647 \$224272 \$223850 \$224002 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13648 VSS|anode|cathode|clk|vss \$224002 R[12]|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13649 VSS|anode|cathode|clk|vss cp|i|z$7 \$224003 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13650 VSS|anode|cathode|clk|vss \$224003 \$223851 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13651 \$224004 \$223851 \$224042 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13652 \$224042 \$224005 \$224043 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13653 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224043
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13654 \$223852 \$224003 \$224006 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13655 VSS|anode|cathode|clk|vss \$224003 \$224041 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13656 \$224041 d|z$73 \$224004 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13657 VSS|anode|cathode|clk|vss \$224004 \$224005 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13658 \$224005 \$223851 \$223852 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13659 VSS|anode|cathode|clk|vss \$224007 \$224006 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13660 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224297
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13661 \$224297 \$223852 \$224007 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13662 VSS|anode|cathode|clk|vss \$224007 R[4]|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13663 VSS|anode|cathode|clk|vss cp|z$4 \$224008 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13664 VSS|anode|cathode|clk|vss \$224008 \$223853 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13665 \$224009 \$223853 \$224039 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13666 \$224039 \$224010 \$224040 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13667 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224040
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13668 \$223854 \$224008 \$224011 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13669 VSS|anode|cathode|clk|vss \$224008 \$224038 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13670 \$224038 d|z$74 \$224009 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13671 VSS|anode|cathode|clk|vss \$224009 \$224010 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13672 \$224010 \$223853 \$223854 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13673 VSS|anode|cathode|clk|vss \$224012 \$224011 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13674 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224336
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13675 \$224336 \$223854 \$224012 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13676 VSS|anode|cathode|clk|vss \$224012 R[44]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13677 VSS|anode|cathode|clk|vss i|z$115 \$224013 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13678 VSS|anode|cathode|clk|vss \$224013 cp|z$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13679 \$224014 s|zn$6 \$224015 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13680 \$224016 \$223855 \$224014 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13681 VSS|anode|cathode|clk|vss i0|i1|q$5 \$224016 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13682 VSS|anode|cathode|clk|vss R[60]|i1|q \$224015 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13683 VSS|anode|cathode|clk|vss s|zn$6 \$223855 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13684 VSS|anode|cathode|clk|vss \$224014 d|z$77 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13685 VSS|anode|cathode|clk|vss cp|z$4 \$224018 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13686 VSS|anode|cathode|clk|vss \$224018 \$223856 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13687 \$224019 \$223856 \$224030 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13688 \$224030 \$224020 \$224031 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13689 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224031
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13690 \$223857 \$224018 \$224021 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13691 VSS|anode|cathode|clk|vss \$224018 \$224035 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13692 \$224035 d|z$77 \$224019 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13693 VSS|anode|cathode|clk|vss \$224019 \$224020 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13694 \$224020 \$223856 \$223857 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13695 VSS|anode|cathode|clk|vss \$224022 \$224021 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13696 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$224429
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13697 \$224429 \$223857 \$224022 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13698 VSS|anode|cathode|clk|vss \$224022 R[60]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13699 VSS|anode|cathode|clk|vss \$226404 RESET_B|RSTB|core|p2c
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$13700 VSS|anode|cathode|clk|vss \$226406 \$227138 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13701 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227837
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13702 \$227837 \$226131 \$226406 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13703 VSS|anode|cathode|clk|vss \$226406 i0|i1|q$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13704 VSS|anode|cathode|clk|vss \$226408 \$227139 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13705 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227841
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13706 \$227841 \$226135 \$226408 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13707 VSS|anode|cathode|clk|vss \$226408 i0|i1|q$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13708 VSS|anode|cathode|clk|vss \$226410 \$227140 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13709 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227846
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13710 \$227846 \$226139 \$226410 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13711 VSS|anode|cathode|clk|vss \$226410 i0|i1|q$10 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13712 VSS|anode|cathode|clk|vss \$226412 \$227141 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13713 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227845
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13714 \$227845 \$226143 \$226412 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13715 VSS|anode|cathode|clk|vss \$226412 DUT_Footer|R[10]|Vdn|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13716 \$226208 s|zn$5 \$226144 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13717 \$226208 i0|i1|q$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13718 VSS|anode|cathode|clk|vss DUT_Footer|R[10]|Vdn|i|i0|q \$226209
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13719 \$226209 \$226113 \$226144 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13720 VSS|anode|cathode|clk|vss s|zn$5 \$226113 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13721 VSS|anode|cathode|clk|vss \$226144 d|z$80 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13722 \$227142 a2|z$12 \$227840 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13723 \$227840 a1|i|i0|i1|q a2|zn$13 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13724 \$227142 a1|a3|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13725 \$226212 s|z$1 \$226145 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13726 \$226212 i0|i1|q$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13727 VSS|anode|cathode|clk|vss DUT_Header|R[3]|Vup|i|i0|q \$226213
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13728 \$226213 \$226114 \$226145 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13729 VSS|anode|cathode|clk|vss s|z$1 \$226114 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13730 VSS|anode|cathode|clk|vss \$226145 d|z$81 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13731 \$226215 s|zn$5 \$226146 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13732 \$226215 i0|i1|q$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13733 VSS|anode|cathode|clk|vss R[14]|i|i0|q \$226216
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13734 \$226216 \$226115 \$226146 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13735 VSS|anode|cathode|clk|vss s|zn$5 \$226115 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13736 VSS|anode|cathode|clk|vss \$226146 d|z$82 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13737 VSS|anode|cathode|clk|vss \$226416 \$227143 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13738 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227827
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13739 \$227827 \$226150 \$226416 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13740 VSS|anode|cathode|clk|vss \$226416 R[14]|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13741 a1|z$15 a1|i|i0|i1|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$13742 VSS|anode|cathode|clk|vss a1|zn$20 \$226219 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13743 \$226219 a2|zn$14 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.263525p AD=0.374525p PS=1.465u PD=2.205u
M$13744 VSS|anode|cathode|clk|vss \$226219 i1|z$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.374525p AD=0.358775p PS=2.205u PD=2.4u
M$13745 \$226221 s|zn$4 \$226151 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13746 \$226221 i0|i1|q$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13747 VSS|anode|cathode|clk|vss R[46]|i0|q \$226222 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13748 \$226222 \$226116 \$226151 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13749 VSS|anode|cathode|clk|vss s|zn$4 \$226116 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13750 VSS|anode|cathode|clk|vss \$226151 d|z$79 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13751 VSS|anode|cathode|clk|vss \$226418 \$227144 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13752 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227812
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13753 \$227812 \$226155 \$226418 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13754 VSS|anode|cathode|clk|vss \$226418 RO_control|R[1]|i|i0|nclk|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13755 VSS|anode|cathode|clk|vss \$226420 \$227145 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13756 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227810
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13757 \$227810 \$226159 \$226420 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13758 VSS|anode|cathode|clk|vss \$226420 DUT_Header|R[11]|Vup|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13759 \$226226 s|z$1 \$226160 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13760 \$226226 i0|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13761 VSS|anode|cathode|clk|vss R[0]|clk|i|i0|n_RO_control|q \$226227
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13762 \$226227 \$226117 \$226160 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13763 VSS|anode|cathode|clk|vss s|z$1 \$226117 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13764 VSS|anode|cathode|clk|vss \$226160 d|z$83 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13765 VSS|anode|cathode|clk|vss \$226423 \$227146 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13766 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227790
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13767 \$227790 \$226164 \$226423 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13768 VSS|anode|cathode|clk|vss \$226423 R[8]|clk|i|i0|n_RO_control|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13769 VSS|anode|cathode|clk|vss \$226425 \$227147 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13770 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227788
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13771 \$227788 \$226168 \$226425 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13772 VSS|anode|cathode|clk|vss \$226425 R[40]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13773 VSS|anode|cathode|clk|vss \$226427 \$227148 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13774 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227780
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13775 \$227780 \$226172 \$226427 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13776 VSS|anode|cathode|clk|vss \$226427 R[59]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13777 DATA|core|i0|i1|p2c \$227998 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$13778 \$226128 cp|i|z$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13779 VSS|anode|cathode|clk|vss \$226128 \$226129 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13780 VSS|anode|cathode|clk|vss \$226128 \$227831 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13781 \$227831 d|z$76 \$226203 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13782 \$226203 \$226129 \$227830 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13783 \$227830 \$226405 \$227829 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13784 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227829
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13785 \$226405 \$226203 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13786 \$226405 \$226129 \$226131 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13787 \$226131 \$226128 \$227138 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13788 \$226132 cp|i|z$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13789 VSS|anode|cathode|clk|vss \$226132 \$226133 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13790 VSS|anode|cathode|clk|vss \$226132 \$227836 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13791 \$227836 d|z$68 \$226204 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13792 \$226204 \$226133 \$227835 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13793 \$227835 \$226407 \$227834 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13794 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227834
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13795 \$226407 \$226204 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13796 \$226407 \$226133 \$226135 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13797 \$226135 \$226132 \$227139 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13798 \$226136 cp|i|z$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13799 VSS|anode|cathode|clk|vss \$226136 \$226137 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13800 VSS|anode|cathode|clk|vss \$226136 \$227839 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13801 \$227839 d|z$84 \$226205 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13802 \$226205 \$226137 \$227838 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13803 \$227838 \$226409 \$227847 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13804 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227847
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13805 \$226409 \$226205 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13806 \$226409 \$226137 \$226139 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13807 \$226139 \$226136 \$227140 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13808 \$226140 cp|i|z$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13809 VSS|anode|cathode|clk|vss \$226140 \$226141 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13810 VSS|anode|cathode|clk|vss \$226140 \$227842 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13811 \$227842 d|z$80 \$226207 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13812 \$226207 \$226141 \$227843 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13813 \$227843 \$226411 \$227844 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13814 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227844
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13815 \$226411 \$226207 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13816 \$226411 \$226141 \$226143 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13817 \$226143 \$226140 \$227141 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13818 \$226147 cp|i|z$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13819 VSS|anode|cathode|clk|vss \$226147 \$226148 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13820 VSS|anode|cathode|clk|vss \$226147 \$227832 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13821 \$227832 d|z$82 \$226218 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13822 \$226218 \$226148 \$227826 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13823 \$227826 \$226415 \$227825 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13824 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227825
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13825 \$226415 \$226218 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13826 \$226415 \$226148 \$226150 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13827 \$226150 \$226147 \$227143 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13828 \$226152 cp|i|z$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13829 VSS|anode|cathode|clk|vss \$226152 \$226153 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13830 VSS|anode|cathode|clk|vss \$226152 \$227818 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13831 \$227818 d|z$85 \$226223 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13832 \$226223 \$226153 \$227820 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13833 \$227820 \$226417 \$227821 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13834 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227821
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13835 \$226417 \$226223 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13836 \$226417 \$226153 \$226155 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13837 \$226155 \$226152 \$227144 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13838 \$226156 cp|i|z$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13839 VSS|anode|cathode|clk|vss \$226156 \$226157 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13840 VSS|anode|cathode|clk|vss \$226156 \$227817 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13841 \$227817 d|z$86 \$226225 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13842 \$226225 \$226157 \$227805 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13843 \$227805 \$226419 \$227808 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13844 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227808
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13845 \$226419 \$226225 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13846 \$226419 \$226157 \$226159 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13847 \$226159 \$226156 \$227145 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13848 \$226161 cp|i|z$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13849 VSS|anode|cathode|clk|vss \$226161 \$226162 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13850 VSS|anode|cathode|clk|vss \$226161 \$227799 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13851 \$227799 d|z$87 \$226229 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13852 \$226229 \$226162 \$227801 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13853 \$227801 \$226422 \$227802 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13854 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227802
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13855 \$226422 \$226229 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13856 \$226422 \$226162 \$226164 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13857 \$226164 \$226161 \$227146 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13858 \$226165 cp|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13859 VSS|anode|cathode|clk|vss \$226165 \$226166 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13860 VSS|anode|cathode|clk|vss \$226165 \$227794 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13861 \$227794 d|z$88 \$226230 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13862 \$226230 \$226166 \$227795 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13863 \$227795 \$226424 \$227796 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13864 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227796
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13865 \$226424 \$226230 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13866 \$226424 \$226166 \$226168 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13867 \$226168 \$226165 \$227147 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13868 \$226169 cp|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13869 VSS|anode|cathode|clk|vss \$226169 \$226170 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13870 VSS|anode|cathode|clk|vss \$226169 \$227789 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13871 \$227789 d|z$89 \$226231 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13872 \$226231 \$226170 \$227777 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13873 \$227777 \$226426 \$227776 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13874 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$227776
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13875 \$226426 \$226231 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13876 \$226426 \$226170 \$226172 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13877 \$226172 \$226169 \$227148 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13878 VSS|anode|cathode|clk|vss cp|i|z$5 \$227910 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13879 VSS|anode|cathode|clk|vss \$227910 \$227880 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13880 \$227911 \$227880 \$228215 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13881 \$228215 \$227913 \$228214 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13882 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$228214
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13883 \$227881 \$227910 \$227914 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13884 VSS|anode|cathode|clk|vss \$227910 \$228396 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13885 \$228396 d|z$90 \$227911 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13886 VSS|anode|cathode|clk|vss \$227911 \$227913 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13887 \$227913 \$227880 \$227881 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13888 VSS|anode|cathode|clk|vss \$227915 \$227914 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13889 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$228397
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13890 \$228397 \$227881 \$227915 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13891 VSS|anode|cathode|clk|vss \$227915 i0|i1|q$11 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13892 \$227917 a2|i|s|zn \$227918 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13893 \$227919 \$227882 \$227917 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13894 VSS|anode|cathode|clk|vss i0|i1|q$9 \$227919 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13895 VSS|anode|cathode|clk|vss i0|i1|q$11 \$227918 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13896 VSS|anode|cathode|clk|vss a2|i|s|zn \$227882 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13897 VSS|anode|cathode|clk|vss \$227917 i0|z$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13898 \$227921 a1|a2|b|q|s \$227922 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13899 \$227923 \$227883 \$227921 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13900 VSS|anode|cathode|clk|vss i0|z$2 \$227923 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13901 VSS|anode|cathode|clk|vss i1|z$3 \$227922 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13902 VSS|anode|cathode|clk|vss a1|a2|b|q|s \$227883
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$13903 VSS|anode|cathode|clk|vss \$227921 d|z$90 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13904 \$227924 a2|i|s|zn \$227925 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13905 \$227926 \$227884 \$227924 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13906 VSS|anode|cathode|clk|vss i0|i1|q$10 \$227926 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13907 VSS|anode|cathode|clk|vss i0|i1|q$8 \$227925 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13908 VSS|anode|cathode|clk|vss a2|i|s|zn \$227884 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13909 VSS|anode|cathode|clk|vss \$227924 i0|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13910 \$227927 a2|i|s|zn \$227928 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13911 \$227929 \$227885 \$227927 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13912 VSS|anode|cathode|clk|vss a1|i0|q$2 \$227929 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13913 VSS|anode|cathode|clk|vss i0|i1|q$10 \$227928 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13914 VSS|anode|cathode|clk|vss a2|i|s|zn \$227885 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13915 VSS|anode|cathode|clk|vss \$227927 i0|z$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13916 \$227931 a1|a2|b|q|s \$227932 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13917 \$227933 \$227886 \$227931 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13918 VSS|anode|cathode|clk|vss i0|z$3 \$227933 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13919 VSS|anode|cathode|clk|vss i1|zn \$227932 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13920 VSS|anode|cathode|clk|vss a1|a2|b|q|s \$227886
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$13921 VSS|anode|cathode|clk|vss \$227931 d|z$84 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13922 VSS|anode|cathode|clk|vss cp|i|z$6 \$227934 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13923 VSS|anode|cathode|clk|vss \$227934 \$227887 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13924 \$227935 \$227887 \$228226 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13925 \$228226 \$227936 \$228223 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13926 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$228223
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13927 \$227888 \$227934 \$227937 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13928 VSS|anode|cathode|clk|vss \$227934 \$228403 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13929 \$228403 d|z$91 \$227935 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13930 VSS|anode|cathode|clk|vss \$227935 \$227936 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13931 \$227936 \$227887 \$227888 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13932 VSS|anode|cathode|clk|vss \$227939 \$227937 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13933 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$228404
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13934 \$228404 \$227888 \$227939 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13935 VSS|anode|cathode|clk|vss \$227939 R[58]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13936 VSS|anode|cathode|clk|vss a2|zn$18 \$228407 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13937 \$228407 a1|zn$7 a1|zn$3 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13938 \$227889 a2|z$12 \$228406 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13939 \$228406 a1|i|i0|i1|q a2|zn$11 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13940 VSS|anode|cathode|clk|vss a1|a3|i|i1|q \$227889
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13941 \$227890 RD[39]|a2|z \$228409 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13942 \$228409 a1|a3|i|i1|q a1|zn$4 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13943 VSS|anode|cathode|clk|vss a2|a3|zn$1 \$227890 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13944 \$227891 RD[28]|a2|z \$228410 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13945 \$228410 a1|a3|z a2|zn$15 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13946 VSS|anode|cathode|clk|vss a2|a3|z$1 \$227891 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13947 VSS|anode|cathode|clk|vss cp|i|z$6 \$227944 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13948 VSS|anode|cathode|clk|vss \$227944 \$227892 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13949 \$227945 \$227892 \$228265 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13950 \$228265 \$227946 \$228264 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13951 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$228264
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13952 \$227893 \$227944 \$227947 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13953 VSS|anode|cathode|clk|vss \$227944 \$228411 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13954 \$228411 d|z$81 \$227945 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13955 VSS|anode|cathode|clk|vss \$227945 \$227946 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13956 \$227946 \$227892 \$227893 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13957 VSS|anode|cathode|clk|vss \$227948 \$227947 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13958 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$228412
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$13959 \$228412 \$227893 \$227948 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13960 VSS|anode|cathode|clk|vss \$227948 DUT_Header|R[3]|Vup|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$13961 VSS|anode|cathode|clk|vss a1|zn$18 \$227949 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13962 VSS|anode|cathode|clk|vss a2|zn$19 \$227949 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.374525p AD=0.263525p PS=2.205u PD=1.465u
M$13963 VSS|anode|cathode|clk|vss \$227949 i1|z$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.374525p AD=0.358775p PS=2.205u PD=2.4u
M$13964 \$227894 RD[33]|a2|z \$228413 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13965 \$228413 a1|a3|i|i1|q a1|zn$5 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13966 VSS|anode|cathode|clk|vss a2|a3|zn$1 \$227894 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13967 VSS|anode|cathode|clk|vss a2|zn$22 \$228415 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13968 \$228415 a1|zn$5 \$227951 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13969 VSS|anode|cathode|clk|vss \$227951 a2|z$11 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13970 VSS|anode|cathode|clk|vss a2|zn$16 \$228414 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13971 \$228414 a1|zn$8 \$227953 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13972 VSS|anode|cathode|clk|vss \$227953 a1|z$16 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13973 \$227895 RD[1]|a2|z \$228417 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13974 \$228417 a1|a3|z a2|zn$16 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13975 VSS|anode|cathode|clk|vss a2|a3|zn$1 \$227895 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13976 \$227896 RD[29]|a2|zn \$228416 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13977 \$228416 a1|a3|z a2|zn$17 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13978 VSS|anode|cathode|clk|vss a2|a3|z$1 \$227896 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13979 \$227897 RD[36]|a2|z \$228420 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13980 \$228420 a1|a3|i|i1|q a3|zn$4 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13981 VSS|anode|cathode|clk|vss a2|a3|zn$1 \$227897 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13982 \$227898 RD[35]|a2|z \$228422 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13983 \$228422 a1|a3|i|i1|q a3|zn$3 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13984 VSS|anode|cathode|clk|vss a2|a3|zn$1 \$227898 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13985 \$227958 s|z$1 \$227959 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13986 \$227960 \$227899 \$227958 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13987 VSS|anode|cathode|clk|vss RO_control|R[1]|i|i0|nclk|q \$227960
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$13988 VSS|anode|cathode|clk|vss i0|i1|q$6 \$227959 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13989 VSS|anode|cathode|clk|vss s|z$1 \$227899 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13990 VSS|anode|cathode|clk|vss \$227958 d|z$85 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13991 VSS|anode|cathode|clk|vss a2|zn$27 \$228424 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13992 \$228424 a1|zn$23 \$227961 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13993 VSS|anode|cathode|clk|vss \$227961 a1|z$17 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13994 VSS|anode|cathode|clk|vss a2|zn$35 \$228423 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13995 \$228423 a1|zn$10 \$227963 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13996 VSS|anode|cathode|clk|vss \$227963 a4|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13997 \$227965 s|zn$5 \$227966 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13998 \$227967 \$227900 \$227965 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13999 VSS|anode|cathode|clk|vss DUT_Header|R[11]|Vup|i|i0|q \$227967
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$14000 VSS|anode|cathode|clk|vss i0|i1|q$1 \$227966 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14001 VSS|anode|cathode|clk|vss s|zn$5 \$227900 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14002 VSS|anode|cathode|clk|vss \$227965 d|z$86 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14003 VSS|anode|cathode|clk|vss cp|i|z$7 \$227968 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14004 VSS|anode|cathode|clk|vss \$227968 \$227901 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14005 \$227969 \$227901 \$228266 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14006 \$228266 \$227970 \$228267 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14007 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$228267
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14008 \$227902 \$227968 \$227971 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14009 VSS|anode|cathode|clk|vss \$227968 \$228425 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14010 \$228425 d|z$83 \$227969 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14011 VSS|anode|cathode|clk|vss \$227969 \$227970 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14012 \$227970 \$227901 \$227902 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14013 VSS|anode|cathode|clk|vss \$227972 \$227971 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14014 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$228427
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14015 \$228427 \$227902 \$227972 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14016 VSS|anode|cathode|clk|vss \$227972 R[0]|clk|i|i0|n_RO_control|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14017 \$227973 s|z$1 \$227974 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14018 \$227975 \$227903 \$227973 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14019 VSS|anode|cathode|clk|vss R[6]|i|i0|q \$227975
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$14020 VSS|anode|cathode|clk|vss i0|i1|q$3 \$227974 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14021 VSS|anode|cathode|clk|vss s|z$1 \$227903 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14022 VSS|anode|cathode|clk|vss \$227973 d|z$92 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14023 \$227977 s|zn$5 \$227978 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14024 \$227979 \$227904 \$227977 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14025 VSS|anode|cathode|clk|vss R[8]|clk|i|i0|n_RO_control|q \$227979
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$14026 VSS|anode|cathode|clk|vss i0|i1|q \$227978 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14027 VSS|anode|cathode|clk|vss s|zn$5 \$227904 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14028 VSS|anode|cathode|clk|vss \$227977 d|z$87 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14029 \$227980 s|zn$5 \$227981 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14030 \$227982 \$227905 \$227980 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14031 VSS|anode|cathode|clk|vss RO_control|R[9]|i|i0|nclk|q \$227982
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$14032 VSS|anode|cathode|clk|vss i0|i1|q$6 \$227981 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14033 VSS|anode|cathode|clk|vss s|zn$5 \$227905 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14034 VSS|anode|cathode|clk|vss \$227980 d|z$93 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14035 \$227984 s|zn$4 \$227985 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14036 \$227986 \$227906 \$227984 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14037 VSS|anode|cathode|clk|vss R[40]|i0|q \$227986 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14038 VSS|anode|cathode|clk|vss i0|i1|q \$227985 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14039 VSS|anode|cathode|clk|vss s|zn$4 \$227906 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14040 VSS|anode|cathode|clk|vss \$227984 d|z$88 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14041 \$227987 s|zn$6 \$227988 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14042 \$227989 \$227907 \$227987 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14043 VSS|anode|cathode|clk|vss i0|i1|q$1 \$227989 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14044 VSS|anode|cathode|clk|vss R[59]|i1|q \$227988 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14045 VSS|anode|cathode|clk|vss s|zn$6 \$227907 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14046 VSS|anode|cathode|clk|vss \$227987 d|z$89 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14047 \$227990 s|zn$4 \$227991 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14048 \$227992 \$227908 \$227990 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14049 VSS|anode|cathode|clk|vss R[45]|i0|q \$227992 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14050 VSS|anode|cathode|clk|vss i0|i1|q$7 \$227991 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14051 VSS|anode|cathode|clk|vss s|zn$4 \$227908 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14052 VSS|anode|cathode|clk|vss \$227990 d|z$94 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14053 \$227994 s|zn$6 \$227995 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14054 \$227996 \$227909 \$227994 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14055 VSS|anode|cathode|clk|vss i0|i1|q$6 \$227996 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14056 VSS|anode|cathode|clk|vss R[57]|i1|q \$227995 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14057 VSS|anode|cathode|clk|vss s|zn$6 \$227909 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14058 VSS|anode|cathode|clk|vss \$227994 d|z$95 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14059 VSS|anode|cathode|clk|vss \$230542 \$230995 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14060 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231503
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14061 \$231503 \$230250 \$230542 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14062 VSS|anode|cathode|clk|vss \$230542 i0|i1|q$12 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14063 \$230253 a1|a2|b|q|s \$230252 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14064 \$230253 i1|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14065 VSS|anode|cathode|clk|vss i0|z$5 \$230254 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14066 \$230254 \$230228 \$230252 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14067 VSS|anode|cathode|clk|vss a1|a2|b|q|s \$230228
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14068 VSS|anode|cathode|clk|vss \$230252 d|z$96 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14069 \$230257 a2|i|s|zn \$230256 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14070 \$230257 i0|i1|q$12 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14071 VSS|anode|cathode|clk|vss i0|i1|q$13 \$230258 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14072 \$230258 \$230229 \$230256 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14073 VSS|anode|cathode|clk|vss a2|i|s|zn \$230229 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14074 VSS|anode|cathode|clk|vss \$230256 i0|z$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14075 a2|d|z a2|i|s|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14076 VSS|anode|cathode|clk|vss \$230546 \$230996 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14077 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231513
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14078 \$231513 \$230263 \$230546 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14079 VSS|anode|cathode|clk|vss \$230546 a1|i0|q$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14080 VSS|anode|cathode|clk|vss \$230548 \$230997 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14081 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231527
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14082 \$231527 \$230267 \$230548 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14083 VSS|anode|cathode|clk|vss \$230548 R[61]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14084 \$230271 s|zn$6 \$230270 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14085 \$230271 R[58]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14086 VSS|anode|cathode|clk|vss i0|i1|q$2 \$230272 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14087 \$230272 \$230232 \$230270 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14088 VSS|anode|cathode|clk|vss s|zn$6 \$230232 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14089 VSS|anode|cathode|clk|vss \$230270 d|z$91 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14090 \$230998 RD[4]|a2|z \$231532 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14091 \$231532 a1|a3|z a1|zn$6 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14092 \$230998 a2|a3|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14093 \$230999 a1|a3|i|i1|q \$231540 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14094 \$231540 a2|z$12 \$231538 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14095 \$231538 a1|i|i0|i1|q a4|zn$3 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14096 \$230999 RD[43]|a4|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14097 \$231000 a1|a3|z \$231536 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14098 \$231536 a2|z$12 \$231535 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14099 \$231535 a1|i|i0|i1|q a1|zn$7 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14100 \$231000 RD[12]|a4|zn VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14101 \$231001 a3|zn$4 \$231543 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14102 \$231543 a2|zn$15 \$231542 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14103 \$231542 a1|zn$6 a2|zn$20 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14104 \$231001 a4|zn$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14105 \$230278 s|zn$4 \$230277 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14106 \$230278 i0|i1|q$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14107 VSS|anode|cathode|clk|vss R[43]|i0|q \$230279 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14108 \$230279 \$230233 \$230277 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14109 VSS|anode|cathode|clk|vss s|zn$4 \$230233 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14110 VSS|anode|cathode|clk|vss \$230277 d|z$78 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14111 \$231002 RD[25]|a2|zn \$231549 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14112 \$231549 a1|a3|z a4|zn$4 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14113 \$231002 a2|a3|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14114 \$231003 a1|a3|z \$231548 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14115 \$231548 a2|i|i0|i1|q \$231553 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14116 \$231553 a1|z$15 a2|zn$21 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14117 \$231003 RD[19]|a4|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14118 \$231004 a3|zn$5 \$231552 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14119 \$231552 a2|z$11 \$231551 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14120 \$231551 a1|z$16 i1|zn VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14121 \$231004 a4|zn$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14122 \$231005 a1|a3|z \$231555 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14123 \$231555 a2|i|i0|i1|q \$231554 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14124 \$231554 a1|z$15 a1|zn$8 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14125 \$231005 RD[17]|a4|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14126 \$231006 a1|a3|z \$231560 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14127 \$231560 a2|i|i0|i1|q \$231559 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14128 \$231559 a1|z$15 a1|zn$9 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14129 \$231006 RD[23]|a4|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14130 a4|z$1 \$230285 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14131 \$231007 a1|a3|i|i1|q \$231562 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14132 \$231562 a2|z$12 \$231561 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14133 \$231561 a1|i|i0|i1|q a3|zn$5 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14134 \$231007 RD[41]|a4|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14135 \$231008 a1|a3|z \$231568 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14136 \$231568 a2|z$12 \$231567 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14137 \$231567 a1|i|i0|i1|q a2|zn$22 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14138 \$231008 RD[9]|a4|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14139 \$231009 a1|a3|i|i1|q \$231564 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14140 \$231564 a2|z$12 \$231573 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14141 \$231573 a1|i|i0|i1|q a2|zn$23 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14142 \$231009 RD[46]|a4|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14143 \$231010 RD[38]|a2|z \$231571 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14144 \$231571 a1|a3|i|i1|q a1|zn$10 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14145 \$231010 a2|a3|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14146 \$231011 RD[7]|a2|zn \$231576 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14147 \$231576 a1|a3|z a2|zn$24 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14148 \$231011 a2|a3|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14149 z$34 cp|i|z$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14150 cp|i|z$7 \$230293 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$14151 VSS|anode|cathode|clk|vss i|z$115 \$230293 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14152 VSS|anode|cathode|clk|vss \$230552 \$231012 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14153 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231590
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14154 \$231590 \$230297 \$230552 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14155 VSS|anode|cathode|clk|vss \$230552 DUT_Footer|R[2]|Vdn|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14156 VSS|anode|cathode|clk|vss \$230554 \$231013 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14157 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231592
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14158 \$231592 \$230302 \$230554 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14159 VSS|anode|cathode|clk|vss \$230554 R[41]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14160 \$230305 s|zn$6 \$230304 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14161 \$230305 R[56]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14162 VSS|anode|cathode|clk|vss i0|i1|q \$230306 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14163 \$230306 \$230236 \$230304 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14164 VSS|anode|cathode|clk|vss s|zn$6 \$230236 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14165 VSS|anode|cathode|clk|vss \$230304 d|z$97 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14166 VSS|anode|cathode|clk|vss \$230556 \$231014 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14167 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231612
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14168 \$231612 \$230311 \$230556 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14169 VSS|anode|cathode|clk|vss \$230556 R[56]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14170 \$230313 s|zn$6 \$230312 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14171 \$230313 R[62]|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14172 VSS|anode|cathode|clk|vss i0|i1|q$3 \$230314 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14173 \$230314 \$230238 \$230312 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14174 VSS|anode|cathode|clk|vss s|zn$6 \$230238 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14175 VSS|anode|cathode|clk|vss \$230312 d|z$98 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14176 \$230227 cp|i|z$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14177 VSS|anode|cathode|clk|vss \$230227 \$230247 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14178 VSS|anode|cathode|clk|vss \$230227 \$231499 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14179 \$231499 d|z$99 \$230248 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14180 \$230248 \$230247 \$231497 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14181 \$231497 \$230541 \$231496 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14182 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231496
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14183 \$230541 \$230248 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14184 \$230541 \$230247 \$230250 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14185 \$230250 \$230227 \$230995 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14186 \$230230 cp|i|z$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14187 VSS|anode|cathode|clk|vss \$230230 \$230260 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14188 VSS|anode|cathode|clk|vss \$230230 \$231510 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14189 \$231510 d|z$100 \$230261 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14190 \$230261 \$230260 \$231517 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14191 \$231517 \$230545 \$231518 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14192 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231518
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14193 \$230545 \$230261 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14194 \$230545 \$230260 \$230263 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14195 \$230263 \$230230 \$230996 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14196 \$230231 cp|i|z$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14197 VSS|anode|cathode|clk|vss \$230231 \$230264 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14198 VSS|anode|cathode|clk|vss \$230231 \$231522 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14199 \$231522 d|z$101 \$230265 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14200 \$230265 \$230264 \$231520 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14201 \$231520 \$230547 \$231519 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14202 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231519
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14203 \$230547 \$230265 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14204 \$230547 \$230264 \$230267 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14205 \$230267 \$230231 \$230997 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14206 VSS|anode|cathode|clk|vss a1|zn$3 \$230269 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14207 \$230269 a2|zn$20 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.263525p AD=0.374525p PS=1.465u PD=2.205u
M$14208 VSS|anode|cathode|clk|vss \$230269 i1|z$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.374525p AD=0.358775p PS=2.205u PD=2.4u
M$14209 VSS|anode|cathode|clk|vss a2|zn$25 \$231556 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14210 \$231556 a1|zn$13 \$230285 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14211 \$230234 cp|i|z$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14212 VSS|anode|cathode|clk|vss \$230234 \$230294 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14213 VSS|anode|cathode|clk|vss \$230234 \$231578 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14214 \$231578 d|z$102 \$230295 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14215 \$230295 \$230294 \$231585 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14216 \$231585 \$230551 \$231583 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14217 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231583
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14218 \$230551 \$230295 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14219 \$230551 \$230294 \$230297 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14220 \$230297 \$230234 \$231012 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14221 \$230235 cp|i|z$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14222 VSS|anode|cathode|clk|vss \$230235 \$230299 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14223 VSS|anode|cathode|clk|vss \$230235 \$231586 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14224 \$231586 d|z$103 \$230300 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14225 \$230300 \$230299 \$231596 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14226 \$231596 \$230553 \$231595 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14227 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231595
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14228 \$230553 \$230300 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14229 \$230553 \$230299 \$230302 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14230 \$230302 \$230235 \$231013 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14231 \$230237 cp|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14232 VSS|anode|cathode|clk|vss \$230237 \$230308 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14233 VSS|anode|cathode|clk|vss \$230237 \$231602 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14234 \$231602 d|z$97 \$230309 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14235 \$230309 \$230308 \$231608 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14236 \$231608 \$230555 \$231607 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14237 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$231607
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14238 \$230555 \$230309 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14239 \$230555 \$230308 \$230311 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14240 \$230311 \$230237 \$231014 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14241 VSS|anode|cathode|clk|vss cp|i|z$5 \$232162 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14242 VSS|anode|cathode|clk|vss \$232162 \$232070 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14243 \$232163 \$232070 \$232469 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14244 \$232469 \$232164 \$232467 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14245 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232467
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14246 \$232071 \$232162 \$232165 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14247 VSS|anode|cathode|clk|vss \$232162 \$232470 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14248 \$232470 d|z$104 \$232163 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14249 VSS|anode|cathode|clk|vss \$232163 \$232164 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14250 \$232164 \$232070 \$232071 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14251 VSS|anode|cathode|clk|vss \$232166 \$232165 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14252 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232472
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14253 \$232472 \$232071 \$232166 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14254 VSS|anode|cathode|clk|vss \$232166 i0|i1|q$13 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14255 VSS|anode|cathode|clk|vss cp|i|z$5 \$232167 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14256 VSS|anode|cathode|clk|vss \$232167 \$232072 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14257 \$232168 \$232072 \$232475 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14258 \$232475 \$232169 \$232474 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14259 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232474
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14260 \$232073 \$232167 \$232170 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14261 VSS|anode|cathode|clk|vss \$232167 \$232473 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14262 \$232473 d|z$96 \$232168 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14263 VSS|anode|cathode|clk|vss \$232168 \$232169 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14264 \$232169 \$232072 \$232073 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14265 VSS|anode|cathode|clk|vss \$232171 \$232170 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14266 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232476
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14267 \$232476 \$232073 \$232171 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14268 VSS|anode|cathode|clk|vss \$232171 a1|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14269 VSS|anode|cathode|clk|vss cp|i|z$5 \$232173 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14270 VSS|anode|cathode|clk|vss \$232173 \$232075 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14271 \$232174 \$232075 \$232479 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14272 \$232479 \$232175 \$232478 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14273 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232478
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14274 \$232076 \$232173 \$232176 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14275 VSS|anode|cathode|clk|vss \$232173 \$232480 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14276 \$232480 d|z$105 \$232174 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14277 VSS|anode|cathode|clk|vss \$232174 \$232175 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14278 \$232175 \$232075 \$232076 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14279 VSS|anode|cathode|clk|vss \$232177 \$232176 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14280 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232481
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14281 \$232481 \$232076 \$232177 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14282 VSS|anode|cathode|clk|vss \$232177 DOUT_DAT|c2p|core|i|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14283 \$232178 a1|zn$12 \$232077 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14284 VSS|anode|cathode|clk|vss b|z \$232077 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.4015p AD=0.2905p PS=2.27u PD=1.53u
M$14285 VSS|anode|cathode|clk|vss \$232178 d|z$100 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.4015p AD=0.3955p PS=2.27u PD=2.53u
M$14286 \$232178 a2|zn$29 \$232077 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14287 VSS|anode|cathode|clk|vss cp|i|z$5 \$232179 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14288 VSS|anode|cathode|clk|vss \$232179 \$232078 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14289 \$232180 \$232078 \$232487 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14290 \$232487 \$232181 \$232486 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14291 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232486
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14292 \$232079 \$232179 \$232182 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14293 VSS|anode|cathode|clk|vss \$232179 \$232488 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14294 \$232488 d|z$106 \$232180 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14295 VSS|anode|cathode|clk|vss \$232180 \$232181 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14296 \$232181 \$232078 \$232079 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14297 VSS|anode|cathode|clk|vss \$232183 \$232182 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14298 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232489
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14299 \$232489 \$232079 \$232183 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14300 VSS|anode|cathode|clk|vss \$232183 R[5]|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14301 \$232185 s|zn$6 \$232186 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14302 \$232187 \$232080 \$232185 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14303 VSS|anode|cathode|clk|vss i0|i1|q$7 \$232187 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14304 VSS|anode|cathode|clk|vss R[61]|i1|q \$232186 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14305 VSS|anode|cathode|clk|vss s|zn$6 \$232080 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14306 VSS|anode|cathode|clk|vss \$232185 d|z$101 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14307 \$232081 a1|a3|i|i1|q \$232493 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14308 \$232493 a2|z$12 \$232492 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14309 \$232492 a1|i|i0|i1|q a3|zn$6 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14310 VSS|anode|cathode|clk|vss RD[40]|a4|z \$232081
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14311 \$232082 a1|a3|z \$232495 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14312 \$232495 a2|i|i0|i1|q \$232494 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14313 \$232494 a1|z$15 a2|zn$18 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14314 VSS|anode|cathode|clk|vss RD[20]|a4|zn \$232082
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14315 \$232083 a1|a3|z \$232497 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14316 \$232497 a2|i|i0|i1|q \$232496 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14317 \$232496 a1|z$15 a3|zn$7 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14318 VSS|anode|cathode|clk|vss RD[16]|a4|zn \$232083
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14319 \$232084 a1|a3|i|i1|q \$232500 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14320 \$232500 a2|z$12 \$232499 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14321 \$232499 a1|i|i0|i1|q a4|zn$5 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14322 VSS|anode|cathode|clk|vss RD[44]|a4|z \$232084
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14323 \$232085 a1|a3|z \$232498 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14324 \$232498 a2|i|i0|i1|q \$232501 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14325 \$232501 a1|z$15 a2|zn$26 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14326 VSS|anode|cathode|clk|vss RD[18]|a4|zn \$232085
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14327 \$232086 a3|zn$7 \$232503 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14328 \$232503 a2|zn$28 \$232502 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14329 \$232502 a1|zn$17 a1|zn$12 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14330 VSS|anode|cathode|clk|vss a4|zn$7 \$232086 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14331 \$232087 RD[0]|a2|z \$232504 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14332 \$232504 a1|a3|z a2|zn$28 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14333 VSS|anode|cathode|clk|vss a2|a3|zn$1 \$232087 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14334 \$232088 a3|zn$3 \$232506 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14335 \$232506 a2|zn$21 \$232507 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14336 \$232507 a1|zn$21 a2|zn$19 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14337 VSS|anode|cathode|clk|vss a4|zn$3 \$232088 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14338 \$232089 a1|a3|z \$232505 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14339 \$232505 a2|i|i0|i1|q \$232508 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14340 \$232508 a1|z$15 a2|zn$27 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14341 VSS|anode|cathode|clk|vss RD[22]|a4|zn \$232089
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14342 \$232090 a1|a3|z \$232510 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14343 \$232510 a2|z$12 \$232509 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14344 \$232509 a1|i|i0|i1|q a1|zn$11 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14345 VSS|anode|cathode|clk|vss RD[13]|a4|zn \$232090
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14346 \$232092 a1|a3|z \$232512 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14347 \$232512 a2|z$12 \$232511 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14348 \$232511 a1|i|i0|i1|q a1|zn$13 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14349 VSS|anode|cathode|clk|vss RD[15]|a4|zn \$232092
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14350 \$232093 a3|zn$10 \$232514 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14351 \$232514 a2|zn$34 \$232513 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14352 \$232513 a1|zn$22 a2|zn$14 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14353 VSS|anode|cathode|clk|vss a4|zn$8 \$232093 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14354 \$232094 a3|zn$11 \$232519 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14355 \$232519 a2|z$13 \$232518 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14356 \$232518 a1|zn$4 i1|zn$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14357 VSS|anode|cathode|clk|vss a4|z$1 \$232094 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14358 \$232095 a1|a3|i|i1|q \$232521 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14359 \$232521 a2|z$12 \$232520 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14360 \$232520 a1|i|i0|i1|q a4|zn$6 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14361 VSS|anode|cathode|clk|vss RD[42]|a4|z \$232095
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14362 \$232096 a1|a3|i|i1|q \$232523 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14363 \$232523 a2|z$12 \$232522 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14364 \$232522 a1|i|i0|i1|q a4|zn$8 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14365 VSS|anode|cathode|clk|vss RD[45]|a4|z \$232096
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14366 \$232097 a3|zn$8 \$232525 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14367 \$232525 a2|zn$23 \$232524 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14368 \$232524 a1|z$17 i1|zn$2 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14369 VSS|anode|cathode|clk|vss a4|z \$232097 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14370 \$232098 RD[30]|a2|z \$232529 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14371 \$232529 a1|a3|z a3|zn$8 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14372 VSS|anode|cathode|clk|vss a2|a3|z$1 \$232098 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14373 \$232196 s|z$1 \$232197 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14374 \$232198 \$232099 \$232196 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14375 VSS|anode|cathode|clk|vss DUT_Footer|R[2]|Vdn|i|i0|q \$232198
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$14376 VSS|anode|cathode|clk|vss i0|i1|q$2 \$232197 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14377 VSS|anode|cathode|clk|vss s|z$1 \$232099 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14378 VSS|anode|cathode|clk|vss \$232196 d|z$102 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14379 VSS|anode|cathode|clk|vss cp|i|z$7 \$232199 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14380 VSS|anode|cathode|clk|vss \$232199 \$232100 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14381 \$232200 \$232100 \$232569 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14382 \$232569 \$232201 \$232565 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14383 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232565
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14384 \$232101 \$232199 \$232202 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14385 VSS|anode|cathode|clk|vss \$232199 \$232579 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14386 \$232579 d|z$107 \$232200 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14387 VSS|anode|cathode|clk|vss \$232200 \$232201 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14388 \$232201 \$232100 \$232101 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14389 VSS|anode|cathode|clk|vss \$232203 \$232202 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14390 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232586
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14391 \$232586 \$232101 \$232203 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14392 VSS|anode|cathode|clk|vss \$232203 R[13]|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14393 VSS|anode|cathode|clk|vss cp|z$4 \$232205 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14394 VSS|anode|cathode|clk|vss \$232205 \$232102 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14395 \$232206 \$232102 \$232652 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14396 \$232652 \$232207 \$232641 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14397 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232641
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14398 \$232103 \$232205 \$232208 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14399 VSS|anode|cathode|clk|vss \$232205 \$232607 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14400 \$232607 d|z$93 \$232206 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14401 VSS|anode|cathode|clk|vss \$232206 \$232207 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14402 \$232207 \$232102 \$232103 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14403 VSS|anode|cathode|clk|vss \$232209 \$232208 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14404 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232655
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14405 \$232655 \$232103 \$232209 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14406 VSS|anode|cathode|clk|vss \$232209 RO_control|R[9]|i|i0|nclk|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14407 VSS|anode|cathode|clk|vss cp|z$4 \$232210 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14408 VSS|anode|cathode|clk|vss \$232210 \$232104 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14409 \$232211 \$232104 \$232659 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14410 \$232659 \$232212 \$232658 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14411 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232658
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14412 \$232105 \$232210 \$232213 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14413 VSS|anode|cathode|clk|vss \$232210 \$232661 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14414 \$232661 d|z$108 \$232211 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14415 VSS|anode|cathode|clk|vss \$232211 \$232212 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14416 \$232212 \$232104 \$232105 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14417 VSS|anode|cathode|clk|vss \$232214 \$232213 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14418 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232663
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14419 \$232663 \$232105 \$232214 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14420 VSS|anode|cathode|clk|vss \$232214 R[42]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14421 VSS|anode|cathode|clk|vss cp|z$4 \$232216 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14422 VSS|anode|cathode|clk|vss \$232216 \$232106 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14423 \$232217 \$232106 \$232660 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14424 \$232660 \$232218 \$232662 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14425 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232662
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14426 \$232107 \$232216 \$232219 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14427 VSS|anode|cathode|clk|vss \$232216 \$232656 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14428 \$232656 d|z$95 \$232217 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14429 VSS|anode|cathode|clk|vss \$232217 \$232218 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14430 \$232218 \$232106 \$232107 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14431 VSS|anode|cathode|clk|vss \$232220 \$232219 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14432 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$232654
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14433 \$232654 \$232107 \$232220 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14434 VSS|anode|cathode|clk|vss \$232220 R[57]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14435 \$234141 a1|a2|b|q|s \$234140 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14436 \$234141 i1|z$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14437 VSS|anode|cathode|clk|vss i0|z$6 \$234142 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14438 \$234142 \$233988 \$234140 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14439 VSS|anode|cathode|clk|vss a1|a2|b|q|s \$233988
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14440 VSS|anode|cathode|clk|vss \$234140 d|z$104 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14441 \$234144 a2|i|s|zn \$234143 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14442 \$234144 i0|i1|q$13 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14443 VSS|anode|cathode|clk|vss i0|i1|q$11 \$234145 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14444 \$234145 \$233989 \$234143 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14445 VSS|anode|cathode|clk|vss a2|i|s|zn \$233989 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14446 VSS|anode|cathode|clk|vss \$234143 i0|z$6 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14447 \$234147 a2|i|s|zn \$234146 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14448 \$234147 a1|i1|q VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14449 VSS|anode|cathode|clk|vss i0|i1|q$12 \$234148 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14450 \$234148 \$233990 \$234146 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14451 VSS|anode|cathode|clk|vss a2|i|s|zn \$233990 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14452 VSS|anode|cathode|clk|vss \$234146 i0|z$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14453 \$234150 a1|a2|b|q|s \$234149 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14454 \$234150 i1|zn$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14455 VSS|anode|cathode|clk|vss i0|z$4 \$234151 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14456 \$234151 \$233991 \$234149 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14457 VSS|anode|cathode|clk|vss a1|a2|b|q|s \$233991
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14458 VSS|anode|cathode|clk|vss \$234149 d|z$99 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14459 d|z$105 \$234152 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14460 \$234415 a1|i0|q$2 \$235358 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14461 \$235358 a2|i|s|zn VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.4015p PS=1.53u PD=2.27u
M$14462 VSS|anode|cathode|clk|vss a1|a2|b|q|s \$234415
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.4015p AD=0.3955p
+ PS=2.27u PD=2.53u
M$14463 b|z \$234415 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14464 \$235181 a2|zn$30 \$235372 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14465 \$235372 a1|a2|b|q|s a2|zn$29 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14466 \$235181 a3|zn$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14467 \$234157 s|z$1 \$234156 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14468 \$234157 i0|i1|q$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14469 VSS|anode|cathode|clk|vss R[5]|i|i0|q \$234158
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$14470 \$234158 \$233992 \$234156 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14471 VSS|anode|cathode|clk|vss s|z$1 \$233992 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14472 VSS|anode|cathode|clk|vss \$234156 d|z$106 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14473 VSS|anode|cathode|clk|vss a2|zn$31 \$235376 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14474 \$235376 a1|zn$15 a1|zn$14 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14475 \$235182 RD[32]|a2|z \$235383 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14476 \$235383 a1|a3|i|i1|q a2|zn$30 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14477 \$235182 a2|a3|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14478 \$235183 RD[34]|a2|z \$235380 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14479 \$235380 a1|a3|i|i1|q a1|zn$15 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14480 \$235183 a2|a3|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14481 \$235184 RD[2]|a2|z \$235389 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14482 \$235389 a1|a3|z a3|zn$9 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14483 \$235184 a2|a3|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14484 \$235185 a1|a3|z \$235387 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14485 \$235387 a2|z$12 \$235385 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14486 \$235385 a1|i|i0|i1|q a2|zn$31 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14487 \$235185 RD[10]|a4|zn VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14488 \$235186 a1|a3|z \$235394 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14489 \$235394 a2|z$12 \$235393 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14490 \$235393 a1|i|i0|i1|q a1|zn$16 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14491 \$235186 RD[11]|a4|zn VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14492 \$235187 a3|zn$9 \$235400 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14493 \$235400 a2|zn$26 \$235399 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14494 \$235399 a1|zn$19 a2|zn$32 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14495 \$235187 a4|zn$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14496 \$235188 a1|a3|z \$235397 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14497 \$235397 a2|z$12 \$235396 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14498 \$235396 a1|i|i0|i1|q a1|zn$17 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14499 \$235188 RD[8]|a4|z VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14500 VSS|anode|cathode|clk|vss a2|zn$33 \$235403 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14501 \$235403 a1|zn$16 a1|zn$18 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14502 \$235189 RD[24]|a2|z \$235402 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14503 \$235402 a1|a3|z a4|zn$7 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14504 \$235189 a2|a3|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14505 \$235190 RD[26]|a2|z \$235406 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14506 \$235406 a1|a3|z a1|zn$19 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14507 \$235190 a2|a3|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14508 \$235191 RD[37]|a2|z \$235405 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14509 \$235405 a1|a3|i|i1|q a3|zn$10 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14510 \$235191 a2|a3|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14511 \$235192 RD[27]|a2|zn \$235408 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14512 \$235408 a1|a3|z a2|zn$33 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14513 \$235192 a2|a3|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14514 \$235193 a1|a3|z \$235407 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14515 \$235407 a2|i|i0|i1|q \$235413 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14516 \$235413 a1|z$15 a2|zn$34 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14517 \$235193 RD[21]|a4|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14518 \$235194 RD[31]|a2|zn \$235411 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14519 \$235411 a1|a3|z a3|zn$11 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14520 \$235194 a2|a3|z$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14521 a2|z$13 \$234173 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14522 VSS|anode|cathode|clk|vss a2|zn$17 \$235414 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14523 \$235414 a1|zn$11 a1|zn$20 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14524 \$235195 a1|a3|i|i1|q \$235429 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14525 \$235429 a2|z$12 \$235428 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14526 \$235428 a1|i|i0|i1|q a2|zn$25 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14527 \$235195 RD[47]|a4|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14528 \$235196 a1|a3|z \$235424 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14529 \$235424 a2|z$12 \$235423 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14530 \$235423 a1|i|i0|i1|q a2|zn$35 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14531 \$235196 RD[14]|a4|zn VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p
+ PS=2.53u PD=4.01u
M$14532 \$235197 RD[3]|a2|z \$235442 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14533 \$235442 a1|a3|z a1|zn$21 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14534 \$235197 a2|a3|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14535 \$235198 RD[5]|a2|zn \$235470 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14536 \$235470 a1|a3|z a1|zn$22 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14537 \$235198 a2|a3|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14538 \$235199 RD[6]|a2|zn \$235457 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14539 \$235457 a1|a3|z a1|zn$23 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14540 \$235199 a2|a3|zn$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14541 \$234180 s|zn$5 \$234179 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14542 \$234180 i0|i1|q$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14543 VSS|anode|cathode|clk|vss R[13]|i|i0|q \$234181
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$14544 \$234181 \$233993 \$234179 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14545 VSS|anode|cathode|clk|vss s|zn$5 \$233993 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14546 VSS|anode|cathode|clk|vss \$234179 d|z$107 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14547 VSS|anode|cathode|clk|vss \$234417 \$235200 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14548 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$235516
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14549 \$235516 \$234186 \$234417 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14550 VSS|anode|cathode|clk|vss \$234417 R[6]|i|i0|q
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14551 \$234188 s|zn$4 \$234187 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14552 \$234188 i0|i1|q$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14553 VSS|anode|cathode|clk|vss R[41]|i0|q \$234189 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14554 \$234189 \$233994 \$234187 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14555 VSS|anode|cathode|clk|vss s|zn$4 \$233994 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14556 VSS|anode|cathode|clk|vss \$234187 d|z$103 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14557 \$234191 s|zn$4 \$234190 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14558 \$234191 i0|i1|q$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14559 VSS|anode|cathode|clk|vss R[42]|i0|q \$234192 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14560 \$234192 \$233995 \$234190 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14561 VSS|anode|cathode|clk|vss s|zn$4 \$233995 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14562 VSS|anode|cathode|clk|vss \$234190 d|z$108 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14563 VSS|anode|cathode|clk|vss \$234419 \$235201 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14564 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$235568
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14565 \$235568 \$234197 \$234419 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14566 VSS|anode|cathode|clk|vss \$234419 R[45]|i0|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14567 VSS|anode|cathode|clk|vss \$234421 \$235202 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14568 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$235576
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p
+ AD=0.2905p PS=2.27u PD=1.53u
M$14569 \$235576 \$234202 \$234421 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14570 VSS|anode|cathode|clk|vss \$234421 R[62]|i1|q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14571 VSS|anode|cathode|clk|vss a2|d|z \$235354 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14572 \$235354 a1|i1|q \$234152 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14573 VSS|anode|cathode|clk|vss a2|zn$24 \$235420 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14574 \$235420 a1|zn$9 \$234173 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14575 \$234182 cp|i|z$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14576 VSS|anode|cathode|clk|vss \$234182 \$234183 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14577 VSS|anode|cathode|clk|vss \$234182 \$235496 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14578 \$235496 d|z$92 \$234184 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14579 \$234184 \$234183 \$235525 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14580 \$235525 \$234416 \$235523 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14581 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$235523
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14582 \$234416 \$234184 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14583 \$234416 \$234183 \$234186 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14584 \$234186 \$234182 \$235200 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14585 \$234193 cp|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14586 VSS|anode|cathode|clk|vss \$234193 \$234194 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14587 VSS|anode|cathode|clk|vss \$234193 \$235553 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14588 \$235553 d|z$94 \$234195 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14589 \$234195 \$234194 \$235550 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14590 \$235550 \$234418 \$235549 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14591 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$235549
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14592 \$234418 \$234195 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14593 \$234418 \$234194 \$234197 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14594 \$234197 \$234193 \$235201 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14595 \$234198 cp|z$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14596 VSS|anode|cathode|clk|vss \$234198 \$234199 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14597 VSS|anode|cathode|clk|vss \$234198 \$235587 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14598 \$235587 d|z$98 \$234200 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14599 \$234200 \$234199 \$235584 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14600 \$235584 \$234420 \$235582 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14601 VSS|anode|cathode|clk|vss RST|a1|b|cdn|core|i|p2c \$235582
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14602 \$234420 \$234200 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14603 \$234420 \$234199 \$234202 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14604 \$234202 \$234198 \$235202 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14605 \$235203 RO_control|R[9]|i|i0|nclk|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=15.6u AS=5.304p AD=5.304p
+ PS=39.36u PD=39.36u
M$14617 \$235203 Vin|Vout Vin VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u
+ W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14621 Vin R[8]|clk|i|i0|n_RO_control|q \$235205 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14622 Vin R[8]|clk|i|i0|n_RO_control|q DUT_gate|core|p2c$1
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p
+ PS=3.28u PD=3.28u
M$14623 \$235206 DUT_Footer|R[10]|Vdn|i|i0|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=15.6u AS=5.304p AD=5.304p
+ PS=39.36u PD=39.36u
M$14635 \$235206 Vin Vin|Vout|core|extra_load|padres VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14639 Vin|Vout|core|extra_load|padres R[8]|clk|i|i0|n_RO_control|q
+ Drain_Sense|Vout|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u
+ W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14640 Vin|Vout|core|extra_load|padres R[8]|clk|i|i0|n_RO_control|q
+ Drain_Force|Vout|core|padres VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u
+ W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14644 VSS|anode|cathode|clk|vss Vin|Vout|core|extra_load|padres Vout
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14648 \$235211 VSS|anode|cathode|clk|vss Vout VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14649 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss Vout
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p
+ PS=3.28u PD=3.28u
M$14650 VSS|anode|cathode|clk|vss Vout IN|Vout VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14654 Vin$1 VSS|anode|cathode|clk|vss IN|Vout VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14655 Vin$2 VSS|anode|cathode|clk|vss IN|Vout VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14656 \$235935 D|Q_N \$236439 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1428p AD=0.0609p PS=1.52u PD=0.71u
M$14657 \$236439 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0609p AD=0.1626p
+ PS=0.71u PD=1.415u
M$14658 VSS|anode|cathode|clk|vss \$236455 \$235757 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1626p AD=0.2516p PS=1.415u PD=2.16u
M$14659 \$235939 \$236456 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u PD=0.8u
M$14660 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$236442
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.0378p
+ PS=0.8u PD=0.6u
M$14661 \$236442 \$235940 \$236456 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0378p AD=0.1428p PS=0.6u PD=1.52u
M$14662 VSS|anode|cathode|clk|vss \$235940 D|Q_N VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.2849p PS=2.16u PD=2.25u
M$14663 \$235941 \$235940 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u PD=1.12u
M$14664 VSS|anode|cathode|clk|vss \$235941 Q VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$14665 \$235943 D|Q_N$1 \$236448 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0609p PS=1.52u PD=0.71u
M$14666 \$236448 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0609p AD=0.1626p
+ PS=0.71u PD=1.415u
M$14667 VSS|anode|cathode|clk|vss \$236457 \$235758 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1626p AD=0.2516p PS=1.415u PD=2.16u
M$14668 \$235947 \$236458 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u PD=0.8u
M$14669 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$236450
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.0378p
+ PS=0.8u PD=0.6u
M$14670 \$236450 \$235948 \$236458 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0378p AD=0.1428p PS=0.6u PD=1.52u
M$14671 VSS|anode|cathode|clk|vss \$235948 D|Q_N$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.2849p PS=2.16u PD=2.25u
M$14672 \$235949 \$235948 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u PD=1.12u
M$14673 VSS|anode|cathode|clk|vss \$235949 Q$1 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$14674 \$235951 D|Q_N$2 \$236453 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0609p PS=1.52u PD=0.71u
M$14675 \$236453 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0609p AD=0.1626p
+ PS=0.71u PD=1.415u
M$14676 VSS|anode|cathode|clk|vss \$236459 \$235759 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1626p AD=0.2516p PS=1.415u PD=2.16u
M$14677 \$235955 \$236460 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u PD=0.8u
M$14678 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$236454
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.0378p
+ PS=0.8u PD=0.6u
M$14679 \$236454 \$235956 \$236460 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0378p AD=0.1428p PS=0.6u PD=1.52u
M$14680 VSS|anode|cathode|clk|vss \$235956 D|Q_N$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.2849p PS=2.16u PD=2.25u
M$14681 \$235957 \$235956 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u PD=1.12u
M$14682 VSS|anode|cathode|clk|vss \$235957 Q$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$14683 \$235959 D|Q_N$3 \$236451 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0609p PS=1.52u PD=0.71u
M$14684 \$236451 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0609p AD=0.1626p
+ PS=0.71u PD=1.415u
M$14685 VSS|anode|cathode|clk|vss \$236461 \$235760 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1626p AD=0.2516p PS=1.415u PD=2.16u
M$14686 \$235963 \$236462 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u PD=0.8u
M$14687 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$236445
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.0378p
+ PS=0.8u PD=0.6u
M$14688 \$236445 \$235964 \$236462 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0378p AD=0.1428p PS=0.6u PD=1.52u
M$14689 VSS|anode|cathode|clk|vss \$235964 D|Q_N$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.2849p PS=2.16u PD=2.25u
M$14690 \$235965 \$235964 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u PD=1.12u
M$14691 VSS|anode|cathode|clk|vss \$235965 Q$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$14692 \$235967 D|Q_N$4 \$236441 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0609p PS=1.52u PD=0.71u
M$14693 \$236441 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0609p AD=0.1626p
+ PS=0.71u PD=1.415u
M$14694 VSS|anode|cathode|clk|vss \$236463 \$235761 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1626p AD=0.2516p PS=1.415u PD=2.16u
M$14695 \$235971 \$236464 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u PD=0.8u
M$14696 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$236440
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.0378p
+ PS=0.8u PD=0.6u
M$14697 \$236440 \$235972 \$236464 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0378p AD=0.1428p PS=0.6u PD=1.52u
M$14698 VSS|anode|cathode|clk|vss \$235972 D|Q_N$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.2849p PS=2.16u PD=2.25u
M$14699 \$235973 \$235972 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u PD=1.12u
M$14700 VSS|anode|cathode|clk|vss \$235973 OUT|Q|c2p|core|i
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p
+ PS=1.12u PD=2.16u
M$14701 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$236436
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.1701p AD=0.0378p
+ PS=1.65u PD=0.6u
M$14702 \$236436 \$235757 \$235937 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0378p AD=0.1428p PS=0.6u PD=1.52u
M$14703 \$235935 \$235938 \$236455 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1296p AD=0.0798p PS=1.52u PD=0.8u
M$14704 \$236455 \$236468 \$235937 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0798p AD=0.2373p PS=0.8u PD=1.97u
M$14705 VSS|anode|cathode|clk|vss \$235938 \$236468 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$14706 VSS|anode|cathode|clk|vss IN|Vout \$235938 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$14707 \$235940 \$235938 \$235939 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.12665p AD=0.1428p PS=1.145u PD=1.52u
M$14708 \$235757 \$236468 \$235940 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.74u AS=0.3473p AD=0.12665p PS=2.71u PD=1.145u
M$14709 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$236446
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.1701p AD=0.0378p
+ PS=1.65u PD=0.6u
M$14710 \$236446 \$235758 \$235945 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0378p AD=0.1428p PS=0.6u PD=1.52u
M$14711 \$235943 \$235946 \$236457 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1296p AD=0.0798p PS=1.52u PD=0.8u
M$14712 \$236457 \$236469 \$235945 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0798p AD=0.2373p PS=0.8u PD=1.97u
M$14713 VSS|anode|cathode|clk|vss \$235946 \$236469 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$14714 VSS|anode|cathode|clk|vss Q \$235946 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$14715 \$235948 \$235946 \$235947 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.12665p AD=0.1428p PS=1.145u PD=1.52u
M$14716 \$235758 \$236469 \$235948 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.74u AS=0.3473p AD=0.12665p PS=2.71u PD=1.145u
M$14717 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$236452
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.1701p AD=0.0378p
+ PS=1.65u PD=0.6u
M$14718 \$236452 \$235759 \$235953 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0378p AD=0.1428p PS=0.6u PD=1.52u
M$14719 \$235951 \$235954 \$236459 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1296p AD=0.0798p PS=1.52u PD=0.8u
M$14720 \$236459 \$236470 \$235953 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0798p AD=0.2373p PS=0.8u PD=1.97u
M$14721 VSS|anode|cathode|clk|vss \$235954 \$236470 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$14722 VSS|anode|cathode|clk|vss Q$1 \$235954 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$14723 \$235956 \$235954 \$235955 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.12665p AD=0.1428p PS=1.145u PD=1.52u
M$14724 \$235759 \$236470 \$235956 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.74u AS=0.3473p AD=0.12665p PS=2.71u PD=1.145u
M$14725 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$236447
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.1701p AD=0.0378p
+ PS=1.65u PD=0.6u
M$14726 \$236447 \$235760 \$235961 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0378p AD=0.1428p PS=0.6u PD=1.52u
M$14727 \$235959 \$235962 \$236461 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1296p AD=0.0798p PS=1.52u PD=0.8u
M$14728 \$236461 \$236471 \$235961 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0798p AD=0.2373p PS=0.8u PD=1.97u
M$14729 VSS|anode|cathode|clk|vss \$235962 \$236471 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$14730 VSS|anode|cathode|clk|vss Q$2 \$235962 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$14731 \$235964 \$235962 \$235963 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.12665p AD=0.1428p PS=1.145u PD=1.52u
M$14732 \$235760 \$236471 \$235964 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.74u AS=0.3473p AD=0.12665p PS=2.71u PD=1.145u
M$14733 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$236443
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.1701p AD=0.0378p
+ PS=1.65u PD=0.6u
M$14734 \$236443 \$235761 \$235969 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0378p AD=0.1428p PS=0.6u PD=1.52u
M$14735 \$235967 \$235970 \$236463 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1296p AD=0.0798p PS=1.52u PD=0.8u
M$14736 \$236463 \$236472 \$235969 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0798p AD=0.2373p PS=0.8u PD=1.97u
M$14737 VSS|anode|cathode|clk|vss \$235970 \$236472 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$14738 VSS|anode|cathode|clk|vss Q$3 \$235970 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$14739 \$235972 \$235970 \$235971 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.12665p AD=0.1428p PS=1.145u PD=1.52u
M$14740 \$235761 \$236472 \$235972 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.74u AS=0.3473p AD=0.12665p PS=2.71u PD=1.145u
M$14741 Vin|Vout VSS|anode|cathode|clk|vss Vin$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14742 Vin|Vout VSS|anode|cathode|clk|vss Vin$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14743 Vin|Vout Vout$1 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14747 Vout$1 VSS|anode|cathode|clk|vss Vin$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14748 Vout$1 VSS|anode|cathode|clk|vss Vin$6 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14749 Vout$1 Vout$2 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14753 Vout$2 VSS|anode|cathode|clk|vss Vin$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14754 Vout$2 VSS|anode|cathode|clk|vss Vin$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14755 Vout$2 Vout$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14759 Vout$3 VSS|anode|cathode|clk|vss Vin$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14760 Vout$3 VSS|anode|cathode|clk|vss Vin$10 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14761 Vout$3 Vout$4 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14765 Vout$4 VSS|anode|cathode|clk|vss Vin$11 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14766 Vout$4 VSS|anode|cathode|clk|vss Vin$12 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14767 Vout$4 Vout$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14771 Vout$5 VSS|anode|cathode|clk|vss Vin$13 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14772 Vout$5 VSS|anode|cathode|clk|vss Vin$14 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14773 Vout$5 Vout$6 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14777 Vout$6 VSS|anode|cathode|clk|vss Vin$15 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14778 Vout$6 VSS|anode|cathode|clk|vss Vin$16 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14779 Vout$6 Vout$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14783 Vout$7 VSS|anode|cathode|clk|vss Vin$17 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14784 Vout$7 VSS|anode|cathode|clk|vss Vin$18 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14785 Vout$7 Vout$8 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14789 Vout$8 VSS|anode|cathode|clk|vss Vin$19 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14790 Vout$8 VSS|anode|cathode|clk|vss Vin$20 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14791 Vout$8 IN|Vout VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$14795 VSS|anode|cathode|clk|vss i \$247856 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14796 VSS|anode|cathode|clk|vss \$247856 RD[4]|a2|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14797 VSS|anode|cathode|clk|vss \$248626 RD[25]|a2|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14798 VSS|anode|cathode|clk|vss i$1 \$247857 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14799 VSS|anode|cathode|clk|vss \$247857 RD[2]|a2|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14800 RD[39]|a2|z \$247858 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14801 VSS|anode|cathode|clk|vss R[7]|i|i0|q \$247858
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14802 RD[20]|a4|zn \$248627 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14803 RD[16]|a4|zn \$248628 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14804 RD[11]|a4|zn \$248629 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14805 VSS|anode|cathode|clk|vss \$248630 RD[27]|a2|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14806 VSS|anode|cathode|clk|vss \$248631 RD[18]|a4|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14807 VSS|anode|cathode|clk|vss \$249521 \$249521 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14808 VSS|anode|cathode|clk|vss R[5]|i|i0|q \$247859
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14809 VSS|anode|cathode|clk|vss \$247859 RD[37]|a2|z
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p
+ PS=2.27u PD=2.53u
M$14810 VSS|anode|cathode|clk|vss \$248632 RD[15]|a4|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14811 VSS|anode|cathode|clk|vss \$249522 \$249522 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14812 VSS|anode|cathode|clk|vss \$248633 RD[10]|a4|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14813 VSS|anode|cathode|clk|vss \$248634 RD[12]|a4|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14814 VSS|anode|cathode|clk|vss i$2 \$247860 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14815 VSS|anode|cathode|clk|vss \$247860 RD[0]|a2|z VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14816 VSS|anode|cathode|clk|vss \$248635 RD[14]|a4|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14817 VSS|anode|cathode|clk|vss \$249523 \$249523 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14818 VSS|anode|cathode|clk|vss \$249524 \$249524 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14819 VSS|anode|cathode|clk|vss R[14]|i|i0|q \$247861
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14820 VSS|anode|cathode|clk|vss \$247861 RD[46]|a4|z
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p
+ PS=2.27u PD=2.53u
M$14821 RD[1]|a2|z \$247862 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$14822 VSS|anode|cathode|clk|vss i$3 \$247862 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14823 \$249525 \$249525 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14824 RD[44]|a4|z \$247863 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14825 VSS|anode|cathode|clk|vss R[12]|i|i0|q \$247863
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14826 RD[29]|a2|zn \$248636 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14827 \$249526 \$249526 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14828 \$249527 \$249527 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14829 RD[31]|a2|zn \$248637 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14830 RD[3]|a2|z \$247864 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$14831 VSS|anode|cathode|clk|vss i$4 \$247864 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14832 VSS|anode|cathode|clk|vss R[15]|i|i0|q \$247865
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14833 VSS|anode|cathode|clk|vss \$247865 RD[47]|a4|z
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p
+ PS=2.27u PD=2.53u
M$14834 VSS|anode|cathode|clk|vss \$248638 RD[5]|a2|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14835 RD[6]|a2|zn \$248639 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14836 RD[7]|a2|zn \$248640 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14837 RD[45]|a4|z \$247866 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14838 VSS|anode|cathode|clk|vss R[13]|i|i0|q \$247866
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14839 RD[36]|a2|z \$247867 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14840 VSS|anode|cathode|clk|vss R[4]|i|i0|q \$247867
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14841 RD[38]|a2|z \$247868 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14842 VSS|anode|cathode|clk|vss R[6]|i|i0|q \$247868
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14843 RD[43]|a4|z \$247869 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14844 VSS|anode|cathode|clk|vss DUT_Header|R[11]|Vup|i|i0|q \$247869
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14845 RD[34]|a2|z \$247870 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14846 VSS|anode|cathode|clk|vss DUT_Footer|R[2]|Vdn|i|i0|q \$247870
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14847 RD[42]|a4|z \$247871 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14848 VSS|anode|cathode|clk|vss DUT_Footer|R[10]|Vdn|i|i0|q \$247871
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14849 RD[33]|a2|z \$247872 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14850 VSS|anode|cathode|clk|vss RO_control|R[1]|i|i0|nclk|q \$247872
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14851 RD[35]|a2|z \$247873 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14852 VSS|anode|cathode|clk|vss DUT_Header|R[3]|Vup|i|i0|q \$247873
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14853 RD[40]|a4|z \$247874 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14854 VSS|anode|cathode|clk|vss R[8]|clk|i|i0|n_RO_control|q \$247874
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14855 RD[32]|a2|z \$247875 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14856 VSS|anode|cathode|clk|vss R[0]|clk|i|i0|n_RO_control|q \$247875
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14857 RD[41]|a4|z \$247876 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p
+ PS=2.53u PD=2.27u
M$14858 VSS|anode|cathode|clk|vss RO_control|R[9]|i|i0|nclk|q \$247876
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p
+ AD=0.19775p PS=2.27u PD=1.83u
M$14859 VSS|anode|cathode|clk|vss \$250730 RD[22]|a4|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14860 VSS|anode|cathode|clk|vss \$250731 RD[13]|a4|zn
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p
+ PS=2.53u PD=2.53u
M$14861 \$249966 \$249966 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14862 VSS|anode|cathode|clk|vss \$252776 DUT_gate|core|p2c
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$14863 CLK|core|i|p2c$1 \$254718 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$14864 VSS|anode|cathode|clk|vss Vin|Vout$1 Vin|Vout$2
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14868 Vin$21 VSS|anode|cathode|clk|vss Vin|Vout$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14869 Vin$22 VSS|anode|cathode|clk|vss Vin|Vout$2 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14870 VSS|anode|cathode|clk|vss Vin|Vout$2 Vin|Vout$3
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14874 Vin$23 VSS|anode|cathode|clk|vss Vin|Vout$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14875 Vin$24 VSS|anode|cathode|clk|vss Vin|Vout$3 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14876 VSS|anode|cathode|clk|vss Vin|Vout$3 Vin|Vout$4
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14880 Vin$25 VSS|anode|cathode|clk|vss Vin|Vout$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14881 Vin$26 VSS|anode|cathode|clk|vss Vin|Vout$4 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14882 VSS|anode|cathode|clk|vss Vin|Vout$4 Vin|Vout$5
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14886 Vin$27 VSS|anode|cathode|clk|vss Vin|Vout$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14887 Vin$28 VSS|anode|cathode|clk|vss Vin|Vout$5 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14888 VSS|anode|cathode|clk|vss Vin|Vout$5 Vin|Vout$6
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14892 Vin$29 VSS|anode|cathode|clk|vss Vin|Vout$6 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14893 Vin$30 VSS|anode|cathode|clk|vss Vin|Vout$6 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14894 VSS|anode|cathode|clk|vss Vin|Vout$6 Vin|Vout$7
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14898 Vin$31 VSS|anode|cathode|clk|vss Vin|Vout$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14899 Vin$32 VSS|anode|cathode|clk|vss Vin|Vout$7 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14900 VSS|anode|cathode|clk|vss Vin|Vout$7 Vin|Vout$8
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14904 Vin$33 VSS|anode|cathode|clk|vss Vin|Vout$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14905 Vin$34 VSS|anode|cathode|clk|vss Vin|Vout$8 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14906 VSS|anode|cathode|clk|vss Vin|Vout$8 Vin|Vout$9
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14910 Vin$35 VSS|anode|cathode|clk|vss Vin|Vout$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14911 Vin$36 VSS|anode|cathode|clk|vss Vin|Vout$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14912 VSS|anode|cathode|clk|vss Vin|Vout$9 Vin|Vout$10
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14916 Vin$37 VSS|anode|cathode|clk|vss Vin|Vout$10 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14917 Vin$38 VSS|anode|cathode|clk|vss Vin|Vout$10 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14918 VSS|anode|cathode|clk|vss Vin|Vout$10 Vin|Vout$11
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14922 Vin$39 VSS|anode|cathode|clk|vss Vin|Vout$11 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14923 Vin$40 VSS|anode|cathode|clk|vss Vin|Vout$11 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14924 VSS|anode|cathode|clk|vss Vin|Vout$11 Vin|Vout$12
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14928 Vin$41 VSS|anode|cathode|clk|vss Vin|Vout$12 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14929 Vin$42 VSS|anode|cathode|clk|vss Vin|Vout$12 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14930 VSS|anode|cathode|clk|vss Vin|Vout$12 Vin|Vout$13
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14934 Vin$43 VSS|anode|cathode|clk|vss Vin|Vout$13 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14935 Vin$44 VSS|anode|cathode|clk|vss Vin|Vout$13 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14936 VSS|anode|cathode|clk|vss Vin|Vout$13 Vin|Vout$14
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14940 Vin$45 VSS|anode|cathode|clk|vss Vin|Vout$14 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14941 Vin$46 VSS|anode|cathode|clk|vss Vin|Vout$14 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14942 VSS|anode|cathode|clk|vss Vin|Vout$14 Vin|Vout$15
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14946 Vin$47 VSS|anode|cathode|clk|vss Vin|Vout$15 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14947 Vin$48 VSS|anode|cathode|clk|vss Vin|Vout$15 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14948 VSS|anode|cathode|clk|vss Vin|Vout$15 Vin|Vout$16
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14952 Vin$49 VSS|anode|cathode|clk|vss Vin|Vout$16 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14953 Vin$50 VSS|anode|cathode|clk|vss Vin|Vout$16 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14954 VSS|anode|cathode|clk|vss Vin|Vout$16 Vin|Vout$17
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14958 Vin$51 VSS|anode|cathode|clk|vss Vin|Vout$17 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14959 Vin$52 VSS|anode|cathode|clk|vss Vin|Vout$17 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14960 VSS|anode|cathode|clk|vss Vin|Vout$17 Vin|Vout$18
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14964 Vin$53 VSS|anode|cathode|clk|vss Vin|Vout$18 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14965 Vin$54 VSS|anode|cathode|clk|vss Vin|Vout$18 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14966 VSS|anode|cathode|clk|vss Vin|Vout$18 Vin|Vout$19
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14970 Vin$55 VSS|anode|cathode|clk|vss Vin|Vout$19 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14971 Vin$56 VSS|anode|cathode|clk|vss Vin|Vout$19 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14972 VSS|anode|cathode|clk|vss Vin|Vout$19 Vin|Vout$20
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14976 Vin$57 VSS|anode|cathode|clk|vss Vin|Vout$20 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14977 Vin$58 VSS|anode|cathode|clk|vss Vin|Vout$20 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14978 VSS|anode|cathode|clk|vss Vin|Vout$20 Vin|Vout$21
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14982 Vin$59 VSS|anode|cathode|clk|vss Vin|Vout$21 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14983 Vin$60 VSS|anode|cathode|clk|vss Vin|Vout$21 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14984 VSS|anode|cathode|clk|vss Vin|Vout$21 Vin|Vout$22
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14988 Vin$61 VSS|anode|cathode|clk|vss Vin|Vout$22 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14989 Vin$62 VSS|anode|cathode|clk|vss Vin|Vout$22 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14990 VSS|anode|cathode|clk|vss Vin|Vout$22 Vin|Vout$23
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$14994 Vin$63 VSS|anode|cathode|clk|vss Vin|Vout$23 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14995 Vin$64 VSS|anode|cathode|clk|vss Vin|Vout$23 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$14996 VSS|anode|cathode|clk|vss Vin|Vout$23 Vin|Vout$24
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15000 Vin$65 VSS|anode|cathode|clk|vss Vin|Vout$24 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15001 Vin$66 VSS|anode|cathode|clk|vss Vin|Vout$24 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15002 VSS|anode|cathode|clk|vss Vin|Vout$24 Vin|Vout$25
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15006 Vin$67 VSS|anode|cathode|clk|vss Vin|Vout$25 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15007 Vin$68 VSS|anode|cathode|clk|vss Vin|Vout$25 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15008 VSS|anode|cathode|clk|vss Vin|Vout$25 Vin|Vout$26
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15012 Vin$69 VSS|anode|cathode|clk|vss Vin|Vout$26 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15013 Vin$70 VSS|anode|cathode|clk|vss Vin|Vout$26 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15014 VSS|anode|cathode|clk|vss Vin|Vout$26 Vin|Vout$27
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15018 Vin$71 VSS|anode|cathode|clk|vss Vin|Vout$27 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15019 Vin$72 VSS|anode|cathode|clk|vss Vin|Vout$27 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15020 VSS|anode|cathode|clk|vss Vin|Vout$27 Vin|Vout$28
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15024 Vin$73 VSS|anode|cathode|clk|vss Vin|Vout$28 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15025 Vin$74 VSS|anode|cathode|clk|vss Vin|Vout$28 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15026 VSS|anode|cathode|clk|vss Vin|Vout$28 Vin|Vout$29
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15030 Vin$75 VSS|anode|cathode|clk|vss Vin|Vout$29 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15031 Vin$76 VSS|anode|cathode|clk|vss Vin|Vout$29 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15032 VSS|anode|cathode|clk|vss Vin|Vout$29 Vin|Vout$30
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15036 Vin$77 VSS|anode|cathode|clk|vss Vin|Vout$30 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15037 Vin$78 VSS|anode|cathode|clk|vss Vin|Vout$30 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15038 VSS|anode|cathode|clk|vss Vin|Vout$30 Vin|Vout$31
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15042 Vin$79 VSS|anode|cathode|clk|vss Vin|Vout$31 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15043 Vin$80 VSS|anode|cathode|clk|vss Vin|Vout$31 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15044 VSS|anode|cathode|clk|vss Vin|Vout$31 Vin|Vout$32
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15048 Vin$81 VSS|anode|cathode|clk|vss Vin|Vout$32 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15049 Vin$82 VSS|anode|cathode|clk|vss Vin|Vout$32 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15050 VSS|anode|cathode|clk|vss Vin|Vout$32 Vin|Vout$33
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15054 Vin$83 VSS|anode|cathode|clk|vss Vin|Vout$33 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15055 Vin$84 VSS|anode|cathode|clk|vss Vin|Vout$33 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15056 VSS|anode|cathode|clk|vss Vin|Vout$33 Vin|Vout$34
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15060 Vin$85 VSS|anode|cathode|clk|vss Vin|Vout$34 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15061 Vin$86 VSS|anode|cathode|clk|vss Vin|Vout$34 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15062 VSS|anode|cathode|clk|vss Vin|Vout$34 Vin|Vout$35
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15066 Vin$87 VSS|anode|cathode|clk|vss Vin|Vout$35 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15067 Vin$88 VSS|anode|cathode|clk|vss Vin|Vout$35 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15068 VSS|anode|cathode|clk|vss Vin|Vout$35 Vin|Vout$36
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15072 Vin$89 VSS|anode|cathode|clk|vss Vin|Vout$36 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15073 Vin$90 VSS|anode|cathode|clk|vss Vin|Vout$36 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15074 VSS|anode|cathode|clk|vss Vin|Vout$36 Vin|Vout$37
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15078 Vin$91 VSS|anode|cathode|clk|vss Vin|Vout$37 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15079 Vin$92 VSS|anode|cathode|clk|vss Vin|Vout$37 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15080 VSS|anode|cathode|clk|vss Vin|Vout$37 Vin|Vout$38
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15084 Vin$93 VSS|anode|cathode|clk|vss Vin|Vout$38 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15085 Vin$94 VSS|anode|cathode|clk|vss Vin|Vout$38 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15086 VSS|anode|cathode|clk|vss Vin|Vout$38 Vin|Vout$39
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15090 Vin$95 VSS|anode|cathode|clk|vss Vin|Vout$39 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15091 Vin$96 VSS|anode|cathode|clk|vss Vin|Vout$39 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15092 VSS|anode|cathode|clk|vss Vin|Vout$39 Vin|Vout$40
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15096 Vin$97 VSS|anode|cathode|clk|vss Vin|Vout$40 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15097 Vin$98 VSS|anode|cathode|clk|vss Vin|Vout$40 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15098 VSS|anode|cathode|clk|vss Vin|Vout$40 Vin|Vout$41
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15102 Vin$99 VSS|anode|cathode|clk|vss Vin|Vout$41 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15103 Vin$100 VSS|anode|cathode|clk|vss Vin|Vout$41 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15104 VSS|anode|cathode|clk|vss Vin|Vout$41 Vin|Vout$42
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15108 Vin$101 VSS|anode|cathode|clk|vss Vin|Vout$42 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15109 Vin$102 VSS|anode|cathode|clk|vss Vin|Vout$42 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15110 VSS|anode|cathode|clk|vss Vin|Vout$42 Vin|Vout$43
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15114 Vin$103 VSS|anode|cathode|clk|vss Vin|Vout$43 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15115 Vin$104 VSS|anode|cathode|clk|vss Vin|Vout$43 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15116 VSS|anode|cathode|clk|vss Vin|Vout$43 Vout$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$15120 Vin$105 VSS|anode|cathode|clk|vss Vout$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15121 Vin$106 VSS|anode|cathode|clk|vss Vout$9 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15122 \$270151 RO_control|R[1]|i|i0|nclk|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=15.6u AS=5.304p AD=5.304p
+ PS=39.36u PD=39.36u
M$15134 \$270151 Vout$9 Vin$107 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u
+ W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$15138 Vin$107 R[0]|clk|i|i0|n_RO_control|q \$270153 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15139 Vin$107 R[0]|clk|i|i0|n_RO_control|q DUT_gate|core|p2c
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p
+ PS=3.28u PD=3.28u
M$15140 \$270154 DUT_Footer|R[2]|Vdn|i|i0|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=15.6u AS=5.304p AD=5.304p
+ PS=39.36u PD=39.36u
M$15152 \$270154 Vin$107 Vin|Vout|core|extra_load|padres$1
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15156 Vin|Vout|core|extra_load|padres$1 R[0]|clk|i|i0|n_RO_control|q
+ Drain_Sense|Vout|core|padres$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u
+ W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15157 Vin|Vout|core|extra_load|padres$1 R[0]|clk|i|i0|n_RO_control|q
+ Drain_Force|Vout|core|padres$1 VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u
+ W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$15161 VSS|anode|cathode|clk|vss Vin|Vout|core|extra_load|padres$1 Vin$110
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15165 \$270157 VSS|anode|cathode|clk|vss Vin$110 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15166 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss Vin$110
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p
+ PS=3.28u PD=3.28u
M$15167 VSS|anode|cathode|clk|vss Vin$110 IN|Vin|Vout VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p PS=13.12u PD=13.12u
M$15171 Vin$108 VSS|anode|cathode|clk|vss IN|Vin|Vout VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15172 Vin$109 VSS|anode|cathode|clk|vss IN|Vin|Vout VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15173 Vin|Vout$1 VSS|anode|cathode|clk|vss Vin$111 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15174 Vin|Vout$1 VSS|anode|cathode|clk|vss Vin$112 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15175 Vin|Vout$1 Vin|Vout$44 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15179 Vin|Vout$44 VSS|anode|cathode|clk|vss Vin$113 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15180 Vin|Vout$44 VSS|anode|cathode|clk|vss Vin$114 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15181 Vin|Vout$44 Vin|Vout$45 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15185 Vin|Vout$45 VSS|anode|cathode|clk|vss Vin$115 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15186 Vin|Vout$45 VSS|anode|cathode|clk|vss Vin$116 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15187 Vin|Vout$45 Vin|Vout$46 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15191 Vin|Vout$46 VSS|anode|cathode|clk|vss Vin$117 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15192 Vin|Vout$46 VSS|anode|cathode|clk|vss Vin$118 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15193 Vin|Vout$46 Vin|Vout$47 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15197 Vin|Vout$47 VSS|anode|cathode|clk|vss Vin$119 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15198 Vin|Vout$47 VSS|anode|cathode|clk|vss Vin$120 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15199 Vin|Vout$47 Vin|Vout$48 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15203 Vin|Vout$48 VSS|anode|cathode|clk|vss Vin$121 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15204 Vin|Vout$48 VSS|anode|cathode|clk|vss Vin$122 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15205 Vin|Vout$48 Vin|Vout$49 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15209 Vin|Vout$49 VSS|anode|cathode|clk|vss Vin$123 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15210 Vin|Vout$49 VSS|anode|cathode|clk|vss Vin$124 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15211 Vin|Vout$49 Vin|Vout$50 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15215 Vin|Vout$50 VSS|anode|cathode|clk|vss Vin$125 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15216 Vin|Vout$50 VSS|anode|cathode|clk|vss Vin$126 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15217 Vin|Vout$50 Vin|Vout$51 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15221 Vin|Vout$51 VSS|anode|cathode|clk|vss Vin$127 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15222 Vin|Vout$51 VSS|anode|cathode|clk|vss Vin$128 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15223 Vin|Vout$51 Vin|Vout$52 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15227 Vin|Vout$52 VSS|anode|cathode|clk|vss Vin$129 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15228 Vin|Vout$52 VSS|anode|cathode|clk|vss Vin$130 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15229 Vin|Vout$52 Vin|Vout$53 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15233 Vin|Vout$53 VSS|anode|cathode|clk|vss Vin$131 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15234 Vin|Vout$53 VSS|anode|cathode|clk|vss Vin$132 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15235 Vin|Vout$53 Vin|Vout$54 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15239 Vin|Vout$54 VSS|anode|cathode|clk|vss Vin$133 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15240 Vin|Vout$54 VSS|anode|cathode|clk|vss Vin$134 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15241 Vin|Vout$54 Vin|Vout$55 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15245 Vin|Vout$55 VSS|anode|cathode|clk|vss Vin$135 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15246 Vin|Vout$55 VSS|anode|cathode|clk|vss Vin$136 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15247 Vin|Vout$55 Vin|Vout$56 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15251 Vin|Vout$56 VSS|anode|cathode|clk|vss Vin$137 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15252 Vin|Vout$56 VSS|anode|cathode|clk|vss Vin$138 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15253 Vin|Vout$56 Vin|Vout$57 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15257 Vin|Vout$57 VSS|anode|cathode|clk|vss Vin$139 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15258 Vin|Vout$57 VSS|anode|cathode|clk|vss Vin$140 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15259 Vin|Vout$57 Vin|Vout$58 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15263 Vin|Vout$58 VSS|anode|cathode|clk|vss Vin$141 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15264 Vin|Vout$58 VSS|anode|cathode|clk|vss Vin$142 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15265 Vin|Vout$58 Vin|Vout$59 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15269 Vin|Vout$59 VSS|anode|cathode|clk|vss Vin$143 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15270 Vin|Vout$59 VSS|anode|cathode|clk|vss Vin$144 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15271 Vin|Vout$59 Vin|Vout$60 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15275 Vin|Vout$60 VSS|anode|cathode|clk|vss Vin$145 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15276 Vin|Vout$60 VSS|anode|cathode|clk|vss Vin$146 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15277 Vin|Vout$60 Vin|Vout$61 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15281 Vin|Vout$61 VSS|anode|cathode|clk|vss Vin$147 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15282 Vin|Vout$61 VSS|anode|cathode|clk|vss Vin$148 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15283 Vin|Vout$61 Vin|Vout$62 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15287 Vin|Vout$62 VSS|anode|cathode|clk|vss Vin$149 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15288 Vin|Vout$62 VSS|anode|cathode|clk|vss Vin$150 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15289 Vin|Vout$62 Vin|Vout$63 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15293 Vin|Vout$63 VSS|anode|cathode|clk|vss Vin$151 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15294 Vin|Vout$63 VSS|anode|cathode|clk|vss Vin$152 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15295 Vin|Vout$63 Vin|Vout$64 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15299 Vin|Vout$64 VSS|anode|cathode|clk|vss Vin$153 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15300 Vin|Vout$64 VSS|anode|cathode|clk|vss Vin$154 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15301 Vin|Vout$64 Vin|Vout$65 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15305 Vin|Vout$65 VSS|anode|cathode|clk|vss Vin$155 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15306 Vin|Vout$65 VSS|anode|cathode|clk|vss Vin$156 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15307 Vin|Vout$65 Vin|Vout$66 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15311 Vin|Vout$66 VSS|anode|cathode|clk|vss Vin$157 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15312 Vin|Vout$66 VSS|anode|cathode|clk|vss Vin$158 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15313 Vin|Vout$66 Vin|Vout$67 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15317 Vin|Vout$67 VSS|anode|cathode|clk|vss Vin$159 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15318 Vin|Vout$67 VSS|anode|cathode|clk|vss Vin$160 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15319 Vin|Vout$67 Vin|Vout$68 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15323 Vin|Vout$68 VSS|anode|cathode|clk|vss Vin$161 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15324 Vin|Vout$68 VSS|anode|cathode|clk|vss Vin$162 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15325 Vin|Vout$68 Vin|Vout$69 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15329 Vin|Vout$69 VSS|anode|cathode|clk|vss Vin$163 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15330 Vin|Vout$69 VSS|anode|cathode|clk|vss Vin$164 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15331 Vin|Vout$69 Vin|Vout$70 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15335 Vin|Vout$70 VSS|anode|cathode|clk|vss Vin$165 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15336 Vin|Vout$70 VSS|anode|cathode|clk|vss Vin$166 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15337 Vin|Vout$70 Vin|Vout$71 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15341 Vin|Vout$71 VSS|anode|cathode|clk|vss Vin$167 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15342 Vin|Vout$71 VSS|anode|cathode|clk|vss Vin$168 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15343 Vin|Vout$71 Vin|Vout$72 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15347 Vin|Vout$72 VSS|anode|cathode|clk|vss Vin$169 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15348 Vin|Vout$72 VSS|anode|cathode|clk|vss Vin$170 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15349 Vin|Vout$72 Vin|Vout$73 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15353 Vin|Vout$73 VSS|anode|cathode|clk|vss Vin$171 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15354 Vin|Vout$73 VSS|anode|cathode|clk|vss Vin$172 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15355 Vin|Vout$73 Vin|Vout$74 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15359 Vin|Vout$74 VSS|anode|cathode|clk|vss Vin$173 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15360 Vin|Vout$74 VSS|anode|cathode|clk|vss Vin$174 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15361 Vin|Vout$74 Vin|Vout$75 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15365 Vin|Vout$75 VSS|anode|cathode|clk|vss Vin$175 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15366 Vin|Vout$75 VSS|anode|cathode|clk|vss Vin$176 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15367 Vin|Vout$75 Vin|Vout$76 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15371 Vin|Vout$76 VSS|anode|cathode|clk|vss Vin$177 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15372 Vin|Vout$76 VSS|anode|cathode|clk|vss Vin$178 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15373 Vin|Vout$76 Vin|Vout$77 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15377 Vin|Vout$77 VSS|anode|cathode|clk|vss Vin$179 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15378 Vin|Vout$77 VSS|anode|cathode|clk|vss Vin$180 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15379 Vin|Vout$77 Vin|Vout$78 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15383 Vin|Vout$78 VSS|anode|cathode|clk|vss Vin$181 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15384 Vin|Vout$78 VSS|anode|cathode|clk|vss Vin$182 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15385 Vin|Vout$78 Vin|Vout$79 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15389 Vin|Vout$79 VSS|anode|cathode|clk|vss Vin$183 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15390 Vin|Vout$79 VSS|anode|cathode|clk|vss Vin$184 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15391 Vin|Vout$79 Vin|Vout$80 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15395 Vin|Vout$80 VSS|anode|cathode|clk|vss Vin$185 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15396 Vin|Vout$80 VSS|anode|cathode|clk|vss Vin$186 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15397 Vin|Vout$80 Vin|Vout$81 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15401 Vin|Vout$81 VSS|anode|cathode|clk|vss Vin$187 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15402 Vin|Vout$81 VSS|anode|cathode|clk|vss Vin$188 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15403 Vin|Vout$81 Vin|Vout$82 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15407 Vin|Vout$82 VSS|anode|cathode|clk|vss Vin$189 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15408 Vin|Vout$82 VSS|anode|cathode|clk|vss Vin$190 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15409 Vin|Vout$82 Vin|Vout$83 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15413 Vin|Vout$83 VSS|anode|cathode|clk|vss Vin$191 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15414 Vin|Vout$83 VSS|anode|cathode|clk|vss Vin$192 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15415 Vin|Vout$83 Vin|Vout$84 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15419 Vin|Vout$84 VSS|anode|cathode|clk|vss Vin$193 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15420 Vin|Vout$84 VSS|anode|cathode|clk|vss Vin$194 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15421 Vin|Vout$84 Vin|Vout$85 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15425 Vin|Vout$85 VSS|anode|cathode|clk|vss Vin$195 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15426 Vin|Vout$85 VSS|anode|cathode|clk|vss Vin$196 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15427 Vin|Vout$85 Vin|Vout$86 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15431 Vin|Vout$86 VSS|anode|cathode|clk|vss Vin$197 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15432 Vin|Vout$86 VSS|anode|cathode|clk|vss Vin$198 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15433 Vin|Vout$86 Vin|Vout$87 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15437 Vin|Vout$87 VSS|anode|cathode|clk|vss Vin$199 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15438 Vin|Vout$87 VSS|anode|cathode|clk|vss Vin$200 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15439 Vin|Vout$87 Vin|Vout$88 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15443 Vin|Vout$88 VSS|anode|cathode|clk|vss Vin$201 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15444 Vin|Vout$88 VSS|anode|cathode|clk|vss Vin$202 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15445 Vin|Vout$88 Vin|Vout$89 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15449 Vin|Vout$89 VSS|anode|cathode|clk|vss Vin$203 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15450 Vin|Vout$89 VSS|anode|cathode|clk|vss Vin$204 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15451 Vin|Vout$89 Vin|Vout$90 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15455 Vin|Vout$90 VSS|anode|cathode|clk|vss Vin$205 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15456 Vin|Vout$90 VSS|anode|cathode|clk|vss Vin$206 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15457 Vin|Vout$90 Vin|Vout$91 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15461 Vin|Vout$91 VSS|anode|cathode|clk|vss Vin$207 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15462 Vin|Vout$91 VSS|anode|cathode|clk|vss Vin$208 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15463 Vin|Vout$91 Vin|Vout$92 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15467 Vin|Vout$92 VSS|anode|cathode|clk|vss Vin$209 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15468 Vin|Vout$92 VSS|anode|cathode|clk|vss Vin$210 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15469 Vin|Vout$92 Vin|Vout$93 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15473 Vin|Vout$93 VSS|anode|cathode|clk|vss Vin$211 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15474 Vin|Vout$93 VSS|anode|cathode|clk|vss Vin$212 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15475 Vin|Vout$93 Vin|Vout$94 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15479 Vin|Vout$94 VSS|anode|cathode|clk|vss Vin$213 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15480 Vin|Vout$94 VSS|anode|cathode|clk|vss Vin$214 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15481 Vin|Vout$94 Vin|Vout$95 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15485 Vin|Vout$95 VSS|anode|cathode|clk|vss Vin$215 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15486 Vin|Vout$95 VSS|anode|cathode|clk|vss Vin$216 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15487 Vin|Vout$95 Vin|Vout$96 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15491 Vin|Vout$96 VSS|anode|cathode|clk|vss Vin$217 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15492 Vin|Vout$96 VSS|anode|cathode|clk|vss Vin$218 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.45u W=1.3u AS=0.442p AD=0.442p PS=3.28u PD=3.28u
M$15493 Vin|Vout$96 IN|Vin|Vout VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.45u W=5.2u AS=1.768p AD=1.768p
+ PS=13.12u PD=13.12u
M$15497 VSS|anode|cathode|clk|vss \$278874 DUT_gate|core|p2c$1
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$15498 OUT|Q|c2p|core|i$1 \$279336 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p
+ PS=2.16u PD=1.12u
M$15499 VSS|anode|cathode|clk|vss \$279856 \$279336 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$15500 D|Q_N$5 \$279856 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2849p AD=0.2516p PS=2.25u PD=2.16u
M$15501 \$279338 \$279856 \$279780 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0378p PS=1.52u PD=0.6u
M$15502 \$279780 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0378p AD=0.0798p
+ PS=0.6u PD=0.8u
M$15503 VSS|anode|cathode|clk|vss \$279338 \$279339 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u PD=1.52u
M$15504 \$279340 \$279857 \$279856 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.74u AS=0.3473p AD=0.12665p PS=2.71u PD=1.145u
M$15505 \$279856 \$279562 \$279339 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.12665p AD=0.1428p PS=1.145u PD=1.52u
M$15506 VSS|anode|cathode|clk|vss Q$4 \$279562 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$15507 VSS|anode|cathode|clk|vss \$279562 \$279857 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$15508 \$279564 \$279857 \$279859 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.2373p AD=0.0798p PS=1.97u PD=0.8u
M$15509 \$279859 \$279562 \$279563 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0798p AD=0.1296p PS=0.8u PD=1.52u
M$15510 \$279564 \$279340 \$279775 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0378p PS=1.52u PD=0.6u
M$15511 \$279775 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0378p AD=0.1701p
+ PS=0.6u PD=1.65u
M$15512 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$279777
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.1626p AD=0.0609p
+ PS=1.415u PD=0.71u
M$15513 \$279777 D|Q_N$5 \$279563 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0609p AD=0.1428p PS=0.71u PD=1.52u
M$15514 VSS|anode|cathode|clk|vss \$279859 \$279340 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1626p AD=0.2516p PS=1.415u PD=2.16u
M$15515 Q$4 \$279341 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u PD=1.12u
M$15516 VSS|anode|cathode|clk|vss \$279860 \$279341 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$15517 D|Q_N$6 \$279860 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2849p AD=0.2516p PS=2.25u PD=2.16u
M$15518 \$279343 \$279860 \$279773 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0378p PS=1.52u PD=0.6u
M$15519 \$279773 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0378p AD=0.0798p
+ PS=0.6u PD=0.8u
M$15520 VSS|anode|cathode|clk|vss \$279343 \$279344 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u PD=1.52u
M$15521 \$279345 \$279861 \$279860 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.74u AS=0.3473p AD=0.12665p PS=2.71u PD=1.145u
M$15522 \$279860 \$279565 \$279344 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.12665p AD=0.1428p PS=1.145u PD=1.52u
M$15523 VSS|anode|cathode|clk|vss Q$5 \$279565 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$15524 VSS|anode|cathode|clk|vss \$279565 \$279861 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$15525 \$279567 \$279861 \$279863 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.2373p AD=0.0798p PS=1.97u PD=0.8u
M$15526 \$279863 \$279565 \$279566 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0798p AD=0.1296p PS=0.8u PD=1.52u
M$15527 \$279567 \$279345 \$279770 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0378p PS=1.52u PD=0.6u
M$15528 \$279770 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0378p AD=0.1701p
+ PS=0.6u PD=1.65u
M$15529 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$279771
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.1626p AD=0.0609p
+ PS=1.415u PD=0.71u
M$15530 \$279771 D|Q_N$6 \$279566 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0609p AD=0.1428p PS=0.71u PD=1.52u
M$15531 VSS|anode|cathode|clk|vss \$279863 \$279345 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1626p AD=0.2516p PS=1.415u PD=2.16u
M$15532 Q$5 \$279346 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u PD=1.12u
M$15533 VSS|anode|cathode|clk|vss \$279864 \$279346 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$15534 D|Q_N$7 \$279864 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2849p AD=0.2516p PS=2.25u PD=2.16u
M$15535 \$279348 \$279864 \$279767 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0378p PS=1.52u PD=0.6u
M$15536 \$279767 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0378p AD=0.0798p
+ PS=0.6u PD=0.8u
M$15537 VSS|anode|cathode|clk|vss \$279348 \$279349 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u PD=1.52u
M$15538 \$279350 \$279865 \$279864 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.74u AS=0.3473p AD=0.12665p PS=2.71u PD=1.145u
M$15539 \$279864 \$279568 \$279349 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.12665p AD=0.1428p PS=1.145u PD=1.52u
M$15540 VSS|anode|cathode|clk|vss Q$6 \$279568 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$15541 VSS|anode|cathode|clk|vss \$279568 \$279865 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$15542 \$279570 \$279865 \$279867 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.2373p AD=0.0798p PS=1.97u PD=0.8u
M$15543 \$279867 \$279568 \$279569 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0798p AD=0.1296p PS=0.8u PD=1.52u
M$15544 \$279570 \$279350 \$279764 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0378p PS=1.52u PD=0.6u
M$15545 \$279764 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0378p AD=0.1701p
+ PS=0.6u PD=1.65u
M$15546 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$279760
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.1626p AD=0.0609p
+ PS=1.415u PD=0.71u
M$15547 \$279760 D|Q_N$7 \$279569 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0609p AD=0.1428p PS=0.71u PD=1.52u
M$15548 VSS|anode|cathode|clk|vss \$279867 \$279350 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1626p AD=0.2516p PS=1.415u PD=2.16u
M$15549 Q$6 \$279351 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u PD=1.12u
M$15550 VSS|anode|cathode|clk|vss \$279868 \$279351 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$15551 D|Q_N$8 \$279868 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2849p AD=0.2516p PS=2.25u PD=2.16u
M$15552 \$279353 \$279868 \$279758 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0378p PS=1.52u PD=0.6u
M$15553 \$279758 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0378p AD=0.0798p
+ PS=0.6u PD=0.8u
M$15554 VSS|anode|cathode|clk|vss \$279353 \$279354 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u PD=1.52u
M$15555 \$279355 \$279869 \$279868 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.74u AS=0.3473p AD=0.12665p PS=2.71u PD=1.145u
M$15556 \$279868 \$279571 \$279354 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.12665p AD=0.1428p PS=1.145u PD=1.52u
M$15557 VSS|anode|cathode|clk|vss Q$7 \$279571 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$15558 VSS|anode|cathode|clk|vss \$279571 \$279869 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$15559 \$279573 \$279869 \$279871 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.2373p AD=0.0798p PS=1.97u PD=0.8u
M$15560 \$279871 \$279571 \$279572 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0798p AD=0.1296p PS=0.8u PD=1.52u
M$15561 \$279573 \$279355 \$279759 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0378p PS=1.52u PD=0.6u
M$15562 \$279759 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0378p AD=0.1701p
+ PS=0.6u PD=1.65u
M$15563 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$279755
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.1626p AD=0.0609p
+ PS=1.415u PD=0.71u
M$15564 \$279755 D|Q_N$8 \$279572 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0609p AD=0.1428p PS=0.71u PD=1.52u
M$15565 VSS|anode|cathode|clk|vss \$279871 \$279355 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1626p AD=0.2516p PS=1.415u PD=2.16u
M$15566 Q$7 \$279356 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u PD=1.12u
M$15567 VSS|anode|cathode|clk|vss \$279872 \$279356 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$15568 D|Q_N$9 \$279872 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.2849p AD=0.2516p PS=2.25u PD=2.16u
M$15569 \$279358 \$279872 \$279754 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0378p PS=1.52u PD=0.6u
M$15570 \$279754 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0378p AD=0.0798p
+ PS=0.6u PD=0.8u
M$15571 VSS|anode|cathode|clk|vss \$279358 \$279359 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u PD=1.52u
M$15572 \$279360 \$279873 \$279872 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.74u AS=0.3473p AD=0.12665p PS=2.71u PD=1.145u
M$15573 \$279872 \$279574 \$279359 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.12665p AD=0.1428p PS=1.145u PD=1.52u
M$15574 VSS|anode|cathode|clk|vss IN|Vin|Vout \$279574
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p
+ AD=0.2516p PS=1.805u PD=2.16u
M$15575 VSS|anode|cathode|clk|vss \$279574 \$279873 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.317325p AD=0.2516p PS=1.805u PD=2.16u
M$15576 \$279576 \$279873 \$279874 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.2373p AD=0.0798p PS=1.97u PD=0.8u
M$15577 \$279874 \$279574 \$279575 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0798p AD=0.1296p PS=0.8u PD=1.52u
M$15578 \$279576 \$279360 \$279750 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.1428p AD=0.0378p PS=1.52u PD=0.6u
M$15579 \$279750 RESET_B|RSTB|core|p2c VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.0378p AD=0.1701p
+ PS=0.6u PD=1.65u
M$15580 VSS|anode|cathode|clk|vss RESET_B|RSTB|core|p2c \$279751
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=0.42u AS=0.1626p AD=0.0609p
+ PS=1.415u PD=0.71u
M$15581 \$279751 D|Q_N$9 \$279575 VSS|anode|cathode|clk|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.0609p AD=0.1428p PS=0.71u PD=1.52u
M$15582 VSS|anode|cathode|clk|vss \$279874 \$279360 VSS|anode|cathode|clk|vss
+ sg13_lv_nmos L=0.13u W=0.74u AS=0.1626p AD=0.2516p PS=1.415u PD=2.16u
M$15583 CEB|a1|core|i|p2c \$280694 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$15584 VSS|anode|cathode|clk|vss OUT|Q|c2p|core|i$1 \$304122
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$15585 VSS|anode|cathode|clk|vss OUT|Q|c2p|core|i$1 \$304123
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$15586 VSS|anode|cathode|clk|vss OUT|Q|c2p|core|i \$304124
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$15587 VSS|anode|cathode|clk|vss OUT|Q|c2p|core|i \$304125
+ VSS|anode|cathode|clk|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$15588 VSSIO|anode|cathode|guard|iovss \$40710 AVDD|anode|cathode|pad|vdd
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p
+ PS=110.9u PD=110.9u
M$15608 VSSIO|anode|cathode|guard|iovss gate|ngate|o
+ anode|cathode|pad|pad_adc_result_0_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$15616 VSSIO|anode|cathode|guard|iovss gate|ngate|o$1
+ anode|cathode|pad|pad_adc_result_1_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$15624 VSSIO|anode|cathode|guard|iovss gate|ngate|o$2
+ anode|cathode|pad|pad_adc_result_2_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$15632 VSSIO|anode|cathode|guard|iovss gate|ngate|o$3
+ anode|cathode|pad|pad_adc_result_3_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$15640 VSSIO|anode|cathode|guard|iovss gate|ngate|o$4
+ anode|cathode|pad|pad_adc_result_4_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$15648 VSSIO|anode|cathode|guard|iovss gate|ngate|o$5
+ anode|cathode|pad|pad_adc_valid_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$15656 VSSIO|anode|cathode|guard|iovss gate|ngate|o$6
+ anode|cathode|pad|pad_adc_sample_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$15664 \$63424 RESULT[0]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15665 VSS|anode|cathode|clk|vss \$63550 \$63425 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15666 VSS|anode|cathode|clk|vss \$63425 gate|ngate|o
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15667 \$63426 RESULT[0]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15668 VSS|anode|cathode|clk|vss \$63551 \$63427 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15669 VSS|anode|cathode|clk|vss \$63427 gate|o|pgate
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15670 \$63428 RESULT[1]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15671 VSS|anode|cathode|clk|vss \$63553 \$63429 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15672 VSS|anode|cathode|clk|vss \$63429 gate|ngate|o$1
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15673 \$63430 RESULT[1]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15674 VSS|anode|cathode|clk|vss \$63554 \$63431 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15675 VSS|anode|cathode|clk|vss \$63431 gate|o|pgate$1
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15676 \$63432 RESULT[2]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15677 VSS|anode|cathode|clk|vss \$63556 \$63433 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15678 VSS|anode|cathode|clk|vss \$63433 gate|ngate|o$2
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15679 \$63434 RESULT[2]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15680 VSS|anode|cathode|clk|vss \$63557 \$63435 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15681 VSS|anode|cathode|clk|vss \$63435 gate|o|pgate$2
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15682 \$63436 RESULT[3]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15683 VSS|anode|cathode|clk|vss \$63559 \$63437 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15684 VSS|anode|cathode|clk|vss \$63437 gate|ngate|o$3
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15685 \$63438 RESULT[3]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15686 VSS|anode|cathode|clk|vss \$63560 \$63439 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15687 VSS|anode|cathode|clk|vss \$63439 gate|o|pgate$3
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15688 \$63440 RESULT[4]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15689 VSS|anode|cathode|clk|vss \$63562 \$63441 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15690 VSS|anode|cathode|clk|vss \$63441 gate|ngate|o$4
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15691 \$63442 RESULT[4]|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15692 VSS|anode|cathode|clk|vss \$63563 \$63443 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15693 VSS|anode|cathode|clk|vss \$63443 gate|o|pgate$4
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15694 \$63444 VALID|a3|c2p|core|i|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15695 VSS|anode|cathode|clk|vss \$63565 \$63445 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15696 VSS|anode|cathode|clk|vss \$63445 gate|ngate|o$5
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15697 \$63446 VALID|a3|c2p|core|i|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15698 VSS|anode|cathode|clk|vss \$63566 \$63447 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15699 VSS|anode|cathode|clk|vss \$63447 gate|o|pgate$5
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15700 \$63448 SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15701 VSS|anode|cathode|clk|vss \$63568 \$63449 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15702 VSS|anode|cathode|clk|vss \$63449 gate|ngate|o$6
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15703 \$63450 SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15704 VSS|anode|cathode|clk|vss \$63569 \$63451 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15705 VSS|anode|cathode|clk|vss \$63451 gate|o|pgate$6
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$15706 VSS|anode|cathode|clk|vss core \$64422 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$15707 VSS|anode|cathode|clk|vss core$1 \$64424 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$15708 VSS|anode|cathode|clk|vss core$2 \$90525 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$15709 VSSIO|anode|cathode|guard|iovss \$104012
+ anode|cathode|pad|pad_adc_vrefp_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$15729 VSSIO|anode|cathode|guard|iovss in|pin2 gate|out
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.5u W=108u AS=23.22p AD=20.52p
+ PS=131.16u PD=112.56u
M$15735 VSSIO|anode|cathode|guard|iovss in|pin2 VSSIO|anode|cathode|guard|iovss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=9.5u W=126u AS=23.94p AD=26.64p
+ PS=131.32u PD=149.92u
M$15755 VSSIO|anode|cathode|guard|iovss gate|out VDD|pad|pin1|supply|vdd
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.6u W=756.8u AS=344.608p AD=349.36p
+ PS=931.04u PD=933.2u
M$15927 VSSIO|anode|cathode|guard|iovss \$123933
+ anode|cathode|pad|pad_adc_vrefn_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$15947 VSSIO|anode|cathode|guard|iovss \$144244
+ anode|cathode|pad|pad_adc_vin_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$15967 VSSIO|anode|cathode|guard|iovss in|pin2$1 gate|out$1
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.5u W=108u AS=23.22p AD=20.52p
+ PS=131.16u PD=112.56u
M$15973 VSSIO|anode|cathode|guard|iovss in|pin2$1
+ VSSIO|anode|cathode|guard|iovss VSS|anode|cathode|clk|vss sg13_hv_nmos L=9.5u
+ W=126u AS=23.94p AD=26.64p PS=131.32u PD=149.92u
M$15993 VSSIO|anode|cathode|guard|iovss gate|out$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.6u W=756.8u AS=344.608p AD=349.36p PS=931.04u PD=933.2u
M$16165 VSSIO|anode|cathode|guard|iovss \$165240
+ anode|cathode|pad|pad_adc_vip_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$16185 VSSIO|anode|cathode|guard|iovss gate|ngate|o$7
+ anode|cathode|pad|pad_miso_pad VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.6u
+ W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$16193 \$198890 DOUT_DAT|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$16194 VSS|anode|cathode|clk|vss \$198889 \$199478 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$16195 VSS|anode|cathode|clk|vss \$199478 gate|ngate|o$7
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$16196 \$200225 DOUT_DAT|c2p|core|i|q VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$16197 VSS|anode|cathode|clk|vss \$200224 \$200540 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$16198 VSS|anode|cathode|clk|vss \$200540 gate|o|pgate$7
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$16199 \$226404 core$3 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$16200 VSS|anode|cathode|clk|vss core$4 \$227998 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$16201 \$252776 core$5 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$16202 VSS|anode|cathode|clk|vss core$6 \$254718 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$16203 \$278874 core$7 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$16204 VSS|anode|cathode|clk|vss core$8 \$280694 VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$16205 gate|o|pgate$8 \$306590 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$16206 \$306590 \$304122 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p PS=4.48u PD=2.28u
M$16207 VSS|anode|cathode|clk|vss OUT|Q|c2p|core|i$1 \$306591
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p
+ PS=2.28u PD=4.48u
M$16208 gate|ngate|o$8 \$306593 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$16209 \$306593 \$304123 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p PS=4.48u PD=2.28u
M$16210 VSS|anode|cathode|clk|vss OUT|Q|c2p|core|i$1 \$306594
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p
+ PS=2.28u PD=4.48u
M$16211 gate|o|pgate$9 \$306596 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$16212 \$306596 \$304124 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p PS=4.48u PD=2.28u
M$16213 VSS|anode|cathode|clk|vss OUT|Q|c2p|core|i \$306597
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p
+ PS=2.28u PD=4.48u
M$16214 gate|ngate|o$9 \$306599 VSS|anode|cathode|clk|vss
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p
+ PS=4.48u PD=4.48u
M$16215 \$306599 \$304125 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p PS=4.48u PD=2.28u
M$16216 VSS|anode|cathode|clk|vss OUT|Q|c2p|core|i \$306600
+ VSS|anode|cathode|clk|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p
+ PS=2.28u PD=4.48u
M$16217 VSSIO|anode|cathode|guard|iovss \$329246
+ anode|cathode|pad|pad_RO_101_Drain_Force_pad VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$16237 VSSIO|anode|cathode|guard|iovss \$329247
+ anode|cathode|pad|pad_RO_101_Drain_Sense_pad VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$16257 VSSIO|anode|cathode|guard|iovss \$329248
+ anode|cathode|pad|pad_RO_101_extra_load_pad VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$16277 VSSIO|anode|cathode|guard|iovss \$329249
+ anode|cathode|pad|pad_RO_13_Drain_Force_pad VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$16297 VSSIO|anode|cathode|guard|iovss \$329250
+ anode|cathode|pad|pad_RO_13_Drain_Sense_pad VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$16317 VSSIO|anode|cathode|guard|iovss \$329251
+ anode|cathode|pad|pad_RO_13_extra_load_pad VSS|anode|cathode|clk|vss
+ sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$16337 VSSIO|anode|cathode|guard|iovss \$329252
+ ROVDD|VDD|anode|cathode|nclk|pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$16357 VSSIO|anode|cathode|guard|iovss \$329253
+ RO2VDD|VDD|anode|cathode|nclk|pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$16377 VSSIO|anode|cathode|guard|iovss gate|ngate|o$8
+ anode|cathode|pad|pad_RO_101_Vout_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$16385 VSSIO|anode|cathode|guard|iovss gate|ngate|o$9
+ anode|cathode|pad|pad_RO_13_Vout_pad VSS|anode|cathode|clk|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$16393 RST|a1|b|cdn|core|i|p2c \$64422 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16394 CLK|core|i|p2c \$64424 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p PS=10.18u PD=10.18u
M$16395 \$63550 RESULT[0]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16396 \$63551 RESULT[0]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16397 \$63553 RESULT[1]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16398 \$63554 RESULT[1]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16399 \$63556 RESULT[2]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16400 \$63557 RESULT[2]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16401 \$63559 RESULT[3]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16402 \$63560 RESULT[3]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16403 \$63562 RESULT[4]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16404 \$63563 RESULT[4]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16405 \$63565 VALID|a3|c2p|core|i|z VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16406 \$63566 VALID|a3|c2p|core|i|z VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16407 \$63568 SAMPLE|a1|c2p|core|i|z VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16408 \$63569 SAMPLE|a1|c2p|core|i|z VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$16409 \$89657 \$89973 \$89657 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16445 \$89658 \$89974 \$89658 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16481 \$89659 \$89975 \$89659 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16517 \$89660 \$89976 \$89660 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16553 \$89661 \$89977 \$89661 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16589 \$89662 \$89978 \$89662 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16625 \$89663 \$89979 \$89663 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16661 \$89664 \$89980 \$89664 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16697 \$89665 \$89981 \$89665 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16733 \$89666 \$89982 \$89666 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16769 GO|a2|core|p2c \$90525 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p PS=10.18u PD=10.18u
M$17130 \$91501 a2|zn d|zn VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$17131 d|zn a1|z \$91501 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$17132 \$91501 b|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$17133 \$94761 \$95239 \$94761 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$17145 \$89973 z$6 \$92959 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17146 \$92959 zn$1 \$92959 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17148 \$89973 zn$1 \$89973 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17161 \$92960 z$6 \$89973 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17164 \$92960 zn$1 \$92960 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17177 \$92961 z$6 \$89973 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17180 \$92961 zn$1 \$92961 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17181 \$94762 \$95240 \$94762 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1382.4u AS=590.976p AD=590.976p PS=2482.56u PD=2482.56u
M$17193 \$89974 z$6 \$92962 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17194 \$92962 zn$1 \$92962 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17196 \$89974 zn$1 \$89974 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17209 \$92963 z$6 \$89974 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17212 \$92963 zn$1 \$92963 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17225 \$92964 z$6 \$89974 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17228 \$92964 zn$1 \$92964 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17241 \$89975 z$6 \$92965 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17242 \$92965 zn$1 \$92965 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17244 \$89975 zn$1 \$89975 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17257 \$92966 z$6 \$89975 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17260 \$92966 zn$1 \$92966 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17273 \$92967 z$6 \$89975 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17276 \$92967 zn$1 \$92967 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17289 \$89976 z$6 \$92968 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17290 \$92968 zn$1 \$92968 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17292 \$89976 zn$1 \$89976 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17305 \$92969 z$6 \$89976 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17308 \$92969 zn$1 \$92969 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17321 \$92970 z$6 \$89976 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17324 \$92970 zn$1 \$92970 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17337 \$89977 z$6 \$92971 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17338 \$92971 zn$1 \$92971 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17340 \$89977 zn$1 \$89977 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17353 \$92972 z$6 \$89977 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17356 \$92972 zn$1 \$92972 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17369 \$92973 z$6 \$89977 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17372 \$92973 zn$1 \$92973 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17385 \$89978 z$6 \$92974 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17386 \$92974 zn$1 \$92974 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17388 \$89978 zn$1 \$89978 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17401 \$92975 z$6 \$89978 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17404 \$92975 zn$1 \$92975 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17417 \$92976 z$6 \$89978 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17420 \$92976 zn$1 \$92976 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17433 \$89979 z$6 \$92977 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17434 \$92977 zn$1 \$92977 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17436 \$89979 zn$1 \$89979 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17449 \$92978 z$6 \$89979 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17452 \$92978 zn$1 \$92978 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17465 \$92979 z$6 \$89979 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17468 \$92979 zn$1 \$92979 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17481 \$89980 z$6 \$92980 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17482 \$92980 zn$1 \$92980 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17484 \$89980 zn$1 \$89980 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17497 \$92981 z$6 \$89980 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17500 \$92981 zn$1 \$92981 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17513 \$92982 z$6 \$89980 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17516 \$92982 zn$1 \$92982 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17529 \$89981 z$6 \$92983 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17530 \$92983 zn$1 \$92983 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17532 \$89981 zn$1 \$89981 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17545 \$92984 z$6 \$89981 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17548 \$92984 zn$1 \$92984 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17561 \$92985 z$6 \$89981 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17564 \$92985 zn$1 \$92985 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17565 \$94763 \$95241 \$94763 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$17577 \$89982 z$6 \$92986 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17578 \$92986 zn$1 \$92986 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17580 \$89982 zn$1 \$89982 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17593 \$92987 z$6 \$89982 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17596 \$92987 zn$1 \$92987 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17609 \$92988 z$6 \$89982 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17612 \$92988 zn$1 \$92988 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17613 VDD|pad|pin1|supply|vdd a1|z$3 \$94525 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$17614 \$94525 a2|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$17615 VDD|pad|pin1|supply|vdd \$94525 d|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$17616 b|zn$1 a1|a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$17617 VDD|pad|pin1|supply|vdd GO|a2|core|p2c b|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$17618 b|zn$1 a2|a3|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$17619 a1|z$1 a1|b|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$17620 a1|z$2 a1|b|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$17981 \$100188 \$100549 \$100188 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$17993 \$95239 z$6 \$98170 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17994 \$98170 zn$1 \$98170 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17996 \$95239 zn$1 \$95239 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$18009 \$98171 z$6 \$95239 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18012 \$98171 zn$1 \$98171 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18025 \$98172 z$6 \$95239 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18028 \$98172 zn$1 \$98172 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18041 \$95240 z$3 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=19.2u
+ AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$18042 a2 z$1 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u
+ AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$18044 \$95240 z$1 \$95240 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$18057 VIP|core|padres z$7 \$95240 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=19.2u AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$18058 \$95240 z$4 \$95240 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$18060 VIP|core|padres z$4 VIP|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$18073 VIN|core|padres z$2 \$95240 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=19.2u AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$18074 \$95240 zn \$95240 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$18076 VIN|core|padres zn VIN|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$18125 \$100189 \$100550 \$100189 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=691.2u AS=295.488p AD=295.488p PS=1241.28u PD=1241.28u
M$18413 \$100190 \$100551 \$100190 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$18425 \$95241 z$6 \$98175 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18426 \$98175 zn$1 \$98175 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18428 \$95241 zn$1 \$95241 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$18441 \$98176 z$6 \$95241 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18444 \$98176 zn$1 \$98176 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18457 \$98177 z$6 \$95241 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18460 \$98177 zn$1 \$98177 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18461 \$97466 \$97411 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$18462 VDD|pad|pin1|supply|vdd cp|z \$97411 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$18463 \$99070 \$98923 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$18464 VDD|pad|pin1|supply|vdd cp|z$1 \$98923 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$18465 \$97412 \$97411 \$97567 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$18466 \$97567 \$97467 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$18467 \$98590 \$97466 \$97562 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$18468 \$97562 \$98130 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$18469 \$97566 d|z$1 \$97412 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$18470 VDD|pad|pin1|supply|vdd \$97412 \$97467 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$18471 VDD|pad|pin1|supply|vdd \$97466 \$97566 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$18472 \$97467 \$97411 \$98590 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$18473 VDD|pad|pin1|supply|vdd \$98590 \$98130 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$18474 VDD|pad|pin1|supply|vdd \$99070 \$100074 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$18475 \$100074 d|zn$1 \$98924 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$18476 \$98924 \$98923 \$100082 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$18477 VDD|pad|pin1|supply|vdd \$98926 \$100082 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$18478 \$98926 \$98924 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$18479 \$98926 \$98923 \$98925 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$18480 \$98925 \$99070 \$100080 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$18481 VDD|pad|pin1|supply|vdd \$99071 \$100080 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$18482 VDD|pad|pin1|supply|vdd \$98925 \$99071 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$18483 \$96412 a2|zn$1 d|zn$1 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$18484 d|zn$1 a1|z$4 \$96412 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$18485 \$96412 b|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$18486 b|i|q$1 \$98130 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$18487 RESULT[3]|c2p|core|i|q \$99071 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$18848 \$105761 \$106210 \$105761 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$18860 \$100549 z$6 \$104013 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18861 \$104013 zn$1 \$104013 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18863 \$100549 zn$1 \$100549 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$18876 \$104014 z$6 \$100549 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18879 \$104014 zn$1 \$104014 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18892 \$104015 z$6 \$100549 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18895 \$104015 zn$1 \$104015 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18992 \$105762 \$106211 \$105762 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=345.6u AS=147.744p AD=147.744p PS=620.64u PD=620.64u
M$19004 \$100550 z$7 VREFH|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$19005 VREFH|core|padres z$4 VREFH|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$19007 \$100550 z$4 \$100550 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19020 a2 z$9 \$100550 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u
+ AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$19021 \$100550 z \$100550 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19023 a2 z a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19036 a2$1 z$8 \$100550 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$19037 \$100550 z$5 \$100550 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19039 a2$1 z$5 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19280 \$105763 \$106212 \$105763 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19292 \$100551 z$6 \$104018 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19293 \$104018 zn$1 \$104018 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19295 \$100551 zn$1 \$100551 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$19308 \$104019 z$6 \$100551 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19311 \$104019 zn$1 \$104019 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19324 \$104020 z$6 \$100551 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19327 \$104020 zn$1 \$104020 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19328 \$102321 \$102317 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$19329 VDD|pad|pin1|supply|vdd cp|z$1 \$102317 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$19330 \$106213 a2|z$2 b|zn VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$19331 b|zn a1|i|q \$106213 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$19332 \$106213 RST|a1|b|cdn|core|i|p2c VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p
+ PS=2.03u PD=3.53u
M$19333 VDD|pad|pin1|supply|vdd \$102321 \$103372 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$19334 \$103372 d|zn$2 \$102318 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$19335 \$102318 \$102317 \$103377 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$19336 VDD|pad|pin1|supply|vdd \$102322 \$103377 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$19337 \$102322 \$102318 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$19338 \$102322 \$102317 \$102319 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$19339 \$102319 \$102321 \$103376 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$19340 VDD|pad|pin1|supply|vdd \$102599 \$103376 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$19341 VDD|pad|pin1|supply|vdd \$102319 \$102599 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$19342 VDD|pad|pin1|supply|vdd a1|z$3 \$105439 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$19343 \$105439 a2|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$19344 VDD|pad|pin1|supply|vdd \$105439 d|z$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$19345 \$106214 a2|zn$2 d|zn$3 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$19346 d|zn$3 a1|z$5 \$106214 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$19347 \$106214 b|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$19348 RESULT[0]|c2p|core|i|q \$102599 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$19709 a1|z$5 RESULT[2]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$19710 b|zn$2 a1|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$19711 VDD|pad|pin1|supply|vdd a2|i|q b|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$19712 b|zn$2 a1|a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$19713 \$107103 \$106574 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$19714 VDD|pad|pin1|supply|vdd cp|z \$106574 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$19715 \$106575 \$106574 \$107099 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$19716 \$107099 \$107104 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$19717 \$107535 \$107103 \$107098 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$19718 \$107098 \$107450 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$19719 \$107146 d|z \$106575 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$19720 VDD|pad|pin1|supply|vdd \$106575 \$107104 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$19721 VDD|pad|pin1|supply|vdd \$107103 \$107146 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$19722 \$107104 \$106574 \$107535 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$19723 VDD|pad|pin1|supply|vdd \$107535 \$107450 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$19724 b|i|q \$107450 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$19725 a1|z$6 a1|b|i|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$19726 \$110666 \$111316 \$110666 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19738 \$106210 z$6 \$108873 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19739 \$108873 zn$1 \$108873 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19741 \$106210 zn$1 \$106210 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$19754 \$108874 z$6 \$106210 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19757 \$108874 zn$1 \$108874 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19770 \$108875 z$6 \$106210 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19773 \$108875 zn$1 \$108875 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19870 \$110667 \$111317 \$110667 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=172.8u AS=73.872p AD=73.872p PS=310.32u PD=310.32u
M$19882 \$106211 z$7 VREFH|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19885 \$106211 z$4 \$106211 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19898 a2 z$12 \$106211 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19899 \$106211 z$11 \$106211 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19901 a2 z$11 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19914 a2$1 z$10 \$106211 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19915 \$106211 z$13 \$106211 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19917 a2$1 z$13 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19918 \$110668 \$111318 \$110668 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19966 \$110669 \$111319 \$110669 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20158 \$110670 \$111320 \$110670 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20170 \$106212 z$6 \$108876 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20171 \$108876 zn$1 \$108876 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20173 \$106212 zn$1 \$106212 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20186 \$108877 z$6 \$106212 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20189 \$108877 zn$1 \$108877 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20202 \$108878 z$6 \$106212 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20205 \$108878 zn$1 \$108878 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20206 \$109960 \$109381 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20207 VDD|pad|pin1|supply|vdd cp|z \$109381 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20208 \$109382 \$109381 \$109826 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$20209 \$109826 \$109383 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$20210 \$110568 \$109960 \$109822 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$20211 \$109822 \$109961 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$20212 \$109997 d|z$2 \$109382 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$20213 VDD|pad|pin1|supply|vdd \$109382 \$109383 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$20214 VDD|pad|pin1|supply|vdd \$109960 \$109997 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$20215 \$109383 \$109381 \$110568 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$20216 VDD|pad|pin1|supply|vdd \$110568 \$109961 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$20217 a1|z$8 RESULT[1]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$20218 VDD|pad|pin1|supply|vdd a2|d|zn \$109359 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20219 \$109359 a1|z$9 d|zn$4 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$20220 d|zn$4 b|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20221 VDD|pad|pin1|supply|vdd a2|zn$3 \$109354 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20222 \$109354 a1|z$6 d|zn$5 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$20223 d|zn$5 b|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20224 b|q \$109961 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$20225 VDD|pad|pin1|supply|vdd i|z$3 \$108456 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$20226 VDD|pad|pin1|supply|vdd \$108456 cp|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$20587 a1|a2|a3|z RST|a1|b|cdn|core|i|p2c VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$20588 VDD|pad|pin1|supply|vdd i|z$3 \$111321 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$20589 VDD|pad|pin1|supply|vdd \$111321 cp|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$20590 \$111624 \$111123 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20591 VDD|pad|pin1|supply|vdd cp|z$1 \$111123 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20592 VDD|pad|pin1|supply|vdd \$111624 \$112415 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$20593 \$112415 d|zn \$111124 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$20594 \$111124 \$111123 \$112416 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$20595 VDD|pad|pin1|supply|vdd \$111322 \$112416 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$20596 \$111322 \$111124 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$20597 \$111322 \$111123 \$111125 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$20598 \$111125 \$111624 \$112417 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$20599 VDD|pad|pin1|supply|vdd \$111626 \$112417 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$20600 VDD|pad|pin1|supply|vdd \$111125 \$111626 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$20601 RESULT[4]|c2p|core|i|q \$111626 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$20602 \$115923 \$116062 \$115923 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20614 \$111316 z$6 \$114146 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20615 \$114146 zn$1 \$114146 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20617 \$111316 zn$1 \$111316 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20630 \$114147 z$6 \$111316 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20633 \$114147 zn$1 \$114147 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20646 \$114148 z$6 \$111316 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20649 \$114148 zn$1 \$114148 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20650 \$115924 \$116063 \$115924 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20698 \$115925 \$116064 \$115925 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20746 \$115926 \$116065 \$115926 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20758 \$111317 z$7 VREFH|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$20761 \$111317 z$4 \$111317 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20774 a2 z$14 \$111317 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$20775 \$111317 z$15 \$111317 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20777 a2 z$15 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20790 a2$1 z$18 \$111317 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$20791 \$111317 z$19 \$111317 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20793 a2$1 z$19 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20794 \$115927 \$116066 \$115927 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20806 \$111318 z$7 VREFH|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20809 \$111318 z$4 \$111318 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20822 a2 z$16 \$111318 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20823 \$111318 z$25 \$111318 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20825 a2 z$25 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20838 a2$1 z$21 \$111318 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20839 \$111318 z$23 \$111318 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20841 a2$1 z$23 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20842 \$115928 \$116067 \$115928 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20854 \$111319 z$7 VREFH|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20857 \$111319 z$4 \$111319 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20870 a2 z$17 \$111319 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20871 \$111319 zn$2 \$111319 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20873 a2 zn$2 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20886 a2$1 z$17 \$111319 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20889 a2$1 zn$2 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20890 \$115929 \$116068 \$115929 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20938 \$115930 \$116069 \$115930 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20986 \$115931 \$116070 \$115931 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$21034 \$115932 \$116071 \$115932 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$21046 \$111320 z$6 \$114150 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21047 \$114150 zn$1 \$114150 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21049 \$111320 zn$1 \$111320 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21062 \$114151 z$6 \$111320 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21065 \$114151 zn$1 \$114151 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21078 \$114152 z$6 \$111320 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21081 \$114152 zn$1 \$114152 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21082 \$114426 \$114135 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21083 VDD|pad|pin1|supply|vdd cp|z \$114135 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21084 VDD|pad|pin1|supply|vdd \$114426 \$115337 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$21085 \$115337 d|z$3 \$114136 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$21086 \$114136 \$114135 \$115332 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$21087 VDD|pad|pin1|supply|vdd \$114153 \$115332 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$21088 \$114153 \$114136 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$21089 \$114153 \$114135 \$114137 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$21090 \$114137 \$114426 \$115333 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$21091 VDD|pad|pin1|supply|vdd \$114513 \$115333 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$21092 VDD|pad|pin1|supply|vdd \$114137 \$114513 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$21093 VDD|pad|pin1|supply|vdd a1|z$7 \$112921 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21094 \$112921 a2|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$21095 VDD|pad|pin1|supply|vdd \$112921 SAMPLE|a1|c2p|core|i|z
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p
+ PS=2.03u PD=3.53u
M$21096 b|i|q$3 \$114513 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$21457 AVDD|anode|cathode|pad|vdd i|z$2 \$125722 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21459 AVDD|anode|cathode|pad|vdd \$125722 i|z$10 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$21463 AVDD|anode|cathode|pad|vdd i|zn \$123934 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21465 AVDD|anode|cathode|pad|vdd \$123934 i|z$5 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$21469 \$116062 z$6 \$119299 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21470 \$119299 zn$1 \$119299 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21471 AVDD|anode|cathode|pad|vdd \$125725 \$125726 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21472 \$125724 i|z$10 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21473 \$123935 i|z|zn$3 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21474 AVDD|anode|cathode|pad|vdd \$123605 \$123936 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21476 \$125725 \$125724 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21477 AVDD|anode|cathode|pad|vdd \$125726 i|z$11 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21478 \$123605 \$123935 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21479 AVDD|anode|cathode|pad|vdd \$123936 i|z$1 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21480 \$116062 zn$1 \$116062 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21481 AVDD|anode|cathode|pad|vdd \$126465 i|z$109 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21483 AVDD|anode|cathode|pad|vdd i|z$14 \$126465 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21484 \$123938 i|z$6 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21490 AVDD|anode|cathode|pad|vdd \$123938 i|z|zn AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21506 \$119300 z$6 \$116062 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21507 AVDD|anode|cathode|pad|vdd i|zn$5 \$125728 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21513 AVDD|anode|cathode|pad|vdd \$125728 z$7 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21531 \$119300 zn$1 \$119300 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21532 \$119301 z$6 \$116062 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21535 \$119301 zn$1 \$119301 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21536 \$116063 z$6 \$119302 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21537 \$119302 zn$1 \$119302 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21539 \$116063 zn$1 \$116063 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21540 \$119303 z$6 \$116063 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21543 \$119303 zn$1 \$119303 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21544 \$119304 z$6 \$116063 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21547 \$119304 zn$1 \$119304 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21548 \$116064 z$6 \$119305 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21549 \$119305 zn$1 \$119305 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21551 \$116064 zn$1 \$116064 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21552 \$119306 z$6 \$116064 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21555 \$119306 zn$1 \$119306 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21556 \$119307 z$6 \$116064 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21559 \$119307 zn$1 \$119307 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21560 \$123941 i|z$7 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21566 AVDD|anode|cathode|pad|vdd \$123941 z$21 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21582 \$116065 z$6 \$119308 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21583 AVDD|anode|cathode|pad|vdd i|zn$2 \$125729 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21589 AVDD|anode|cathode|pad|vdd \$125729 i|z|zn$1 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21605 \$119308 zn$1 \$119308 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21607 \$116065 zn$1 \$116065 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21608 \$119309 z$6 \$116065 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21611 \$119309 zn$1 \$119309 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21612 \$119310 z$6 \$116065 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21615 \$119310 zn$1 \$119310 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21616 \$116066 z$6 \$119311 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21617 \$119311 zn$1 \$119311 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21619 \$116066 zn$1 \$116066 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21620 \$119312 z$6 \$116066 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21621 AVDD|anode|cathode|pad|vdd i|z$16 \$125731 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21627 AVDD|anode|cathode|pad|vdd \$125731 z$15 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21645 \$119312 zn$1 \$119312 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21646 \$119313 z$6 \$116066 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21649 \$119313 zn$1 \$119313 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21650 \$116067 z$6 \$119314 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21651 \$119314 zn$1 \$119314 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21653 \$116067 zn$1 \$116067 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21654 \$119315 z$6 \$116067 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21657 \$119315 zn$1 \$119315 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21658 \$119316 z$6 \$116067 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21661 \$119316 zn$1 \$119316 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21662 \$116068 z$6 \$119317 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21663 \$119317 zn$1 \$119317 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21665 \$116068 zn$1 \$116068 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21666 \$119318 z$6 \$116068 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21669 \$119318 zn$1 \$119318 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21670 \$119319 z$6 \$116068 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21673 AVDD|anode|cathode|pad|vdd \$125733 \$125734 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21674 \$125732 i|zn$8 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21675 \$119319 zn$1 \$119319 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21676 \$125733 \$125732 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21677 AVDD|anode|cathode|pad|vdd \$125734 i|z$12 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21678 i|zn$1 i|z|zn$1 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21686 \$116069 z$6 \$119320 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21687 \$119320 zn$1 \$119320 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21689 \$116069 zn$1 \$116069 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21690 \$119321 z$6 \$116069 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21693 \$119321 zn$1 \$119321 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21694 \$119322 z$6 \$116069 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21697 \$119322 zn$1 \$119322 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21698 \$116070 z$6 \$119323 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21699 \$119323 zn$1 \$119323 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21700 AVDD|anode|cathode|pad|vdd \$125738 \$125739 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21701 \$125737 i|z$15 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21703 \$125738 \$125737 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21704 AVDD|anode|cathode|pad|vdd \$125739 i|z$13 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21705 \$116070 zn$1 \$116070 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21706 AVDD|anode|cathode|pad|vdd RESULT[1]|c2p|core|i|q \$125741
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p
+ AD=2.8813375p PS=12.07u PD=12.18u
M$21712 AVDD|anode|cathode|pad|vdd \$125741 i|z|zn$2 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21728 \$119324 z$6 \$116070 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21731 \$119324 zn$1 \$119324 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21732 \$119325 z$6 \$116070 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21735 \$119325 zn$1 \$119325 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21736 AVDD|anode|cathode|pad|vdd \$125744 \$125745 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21737 \$125743 i|z|zn$5 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21738 \$116071 z$6 \$119326 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21739 AVDD|anode|cathode|pad|vdd \$124161 i|z$9 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21741 AVDD|anode|cathode|pad|vdd i|z$8 \$124161 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21742 \$125744 \$125743 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21743 AVDD|anode|cathode|pad|vdd \$125745 i|z$81 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21744 \$119326 zn$1 \$119326 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21746 \$116071 zn$1 \$116071 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21747 \$119327 z$6 \$116071 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21750 \$119327 zn$1 \$119327 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21751 \$119328 z$6 \$116071 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$21754 \$119328 zn$1 \$119328 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$21755 VDD|pad|pin1|supply|vdd a1|i|q \$120240 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$21756 VDD|pad|pin1|supply|vdd a2|i|q \$120241 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.4185p PS=2.03u PD=2.03u
M$21757 \$120241 \$120240 \$120242 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.4185p AD=0.249p PS=2.03u PD=1.43u
M$21758 \$120242 a1|i|q \$120243 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.249p AD=0.249p PS=1.43u PD=1.43u
M$21759 VDD|pad|pin1|supply|vdd \$120241 \$120243 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.249p PS=2.03u PD=1.43u
M$21760 VDD|pad|pin1|supply|vdd \$120242 a2|a3|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$21761 \$118852 i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.339p AD=0.4185p PS=2.33u PD=2.03u
M$21762 VDD|pad|pin1|supply|vdd \$118852 i|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$21763 a2|zn$4 a1|b|i|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21764 VDD|pad|pin1|supply|vdd a1|a2|a3|z a2|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$21765 a2|zn$4 a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21766 \$125747 \$125626 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21767 VDD|pad|pin1|supply|vdd cp|z$2 \$125626 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21768 \$123943 \$123606 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21769 VDD|pad|pin1|supply|vdd cp|z$2 \$123606 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21770 a2|z$2 a2|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$21771 \$125627 \$125626 \$126068 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$21772 \$126068 \$125748 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$21773 \$126892 \$125747 \$126083 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$21774 \$126083 \$126468 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$21775 \$126100 d|zn$8 \$125627 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$21776 VDD|pad|pin1|supply|vdd \$125627 \$125748 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$21777 VDD|pad|pin1|supply|vdd \$125747 \$126100 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$21778 \$125748 \$125626 \$126892 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$21779 VDD|pad|pin1|supply|vdd \$126892 \$126468 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$21780 a2|z$3 \$120244 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21781 VDD|pad|pin1|supply|vdd b|i|q$2 \$121694 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$21782 \$121694 a1|b|i|q$1 \$120244 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$21783 \$120244 a2|zn$5 \$121694 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21784 VDD|pad|pin1|supply|vdd \$123943 \$125498 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$21785 \$125498 d|zn$7 \$123607 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$21786 \$123607 \$123606 \$125473 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$21787 VDD|pad|pin1|supply|vdd \$123944 \$125473 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$21788 \$123944 \$123607 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$21789 \$123944 \$123606 \$123608 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$21790 \$123608 \$123943 \$125476 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$21791 VDD|pad|pin1|supply|vdd \$124164 \$125476 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$21792 VDD|pad|pin1|supply|vdd \$123608 \$124164 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$21793 VDD|pad|pin1|supply|vdd a2|zn$3 \$119232 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21794 \$119232 a1|z$10 d|zn$6 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$21795 d|zn$6 b|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21796 z$20 i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$21797 VDD|pad|pin1|supply|vdd a1|i|q \$120245 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21798 \$120245 a2|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$21799 VDD|pad|pin1|supply|vdd \$120245 VALID|a3|c2p|core|i|z
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p
+ PS=2.03u PD=3.53u
M$21800 a1|b|i|q$3 \$126468 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$21801 RESULT[1]|c2p|core|i|q \$124164 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$21802 AVDD|anode|cathode|pad|vdd \$127549 i|z$75 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21804 AVDD|anode|cathode|pad|vdd i|z \$127549 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21805 i|z|zn$1 i|zn$1 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21813 \$127371 i|z$67 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21819 AVDD|anode|cathode|pad|vdd \$127371 z$4 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21835 \$127372 i|z$17 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21836 AVDD|anode|cathode|pad|vdd \$127110 \$127373 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21837 \$127110 \$127372 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21838 AVDD|anode|cathode|pad|vdd \$127373 i|z$19 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21839 AVDD|anode|cathode|pad|vdd \$127550 i|z$20 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21841 AVDD|anode|cathode|pad|vdd i|z$26 \$127550 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21842 AVDD|anode|cathode|pad|vdd \$127552 i|z$21 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21844 AVDD|anode|cathode|pad|vdd i|z$27 \$127552 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21845 \$127378 i|z$22 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21851 AVDD|anode|cathode|pad|vdd \$127378 z$12 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21867 \$127379 RESULT[4]|c2p|core|i|q AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p
+ AD=2.713175p PS=12.18u PD=12.07u
M$21873 AVDD|anode|cathode|pad|vdd \$127379 i|z|zn$4 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21889 \$127382 i|z$23 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21895 AVDD|anode|cathode|pad|vdd \$127382 a1|i|z|zn
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p
+ PS=32.48u PD=33.98u
M$21911 \$127384 i|z$18 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21912 AVDD|anode|cathode|pad|vdd \$127112 \$127385 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21913 \$127112 \$127384 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21914 AVDD|anode|cathode|pad|vdd \$127385 i|z$31 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21915 i|zn$3 i|z|zn$5 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21923 \$127387 RESULT[2]|c2p|core|i|q AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p
+ AD=2.713175p PS=12.18u PD=12.07u
M$21929 AVDD|anode|cathode|pad|vdd \$127387 i|z|zn$5 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21945 \$127389 i|z$36 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21951 AVDD|anode|cathode|pad|vdd \$127389 z$1 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21967 AVDD|anode|cathode|pad|vdd \$127554 i|z$106 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21969 AVDD|anode|cathode|pad|vdd i|z$28 \$127554 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21970 AVDD|anode|cathode|pad|vdd \$127556 i|z$24 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21972 AVDD|anode|cathode|pad|vdd i|z$12 \$127556 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21973 AVDD|anode|cathode|pad|vdd \$127557 i|z$15 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21975 AVDD|anode|cathode|pad|vdd i|z$29 \$127557 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21976 i|z|zn$6 i|zn$6 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21984 \$127392 i|zn$6 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21985 AVDD|anode|cathode|pad|vdd \$127114 \$127393 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21986 \$127114 \$127392 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21987 AVDD|anode|cathode|pad|vdd \$127393 i|z$8 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21988 i|z|zn$3 i|zn$4 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21996 VDD|pad|pin1|supply|vdd i|z$30 \$127394 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$21997 VDD|pad|pin1|supply|vdd \$127394 i|z$25 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$21998 VDD|pad|pin1|supply|vdd CLK|core|i|p2c \$127396 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$21999 VDD|pad|pin1|supply|vdd \$127396 i|z$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$22000 i|zn$4 i|z|zn$3 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22008 i|zn$5 i|z|zn AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22016 AVDD|anode|cathode|pad|vdd a2|z$5 \$128987 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22017 \$128987 a1|z$12 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=0.996p AD=0.996p PS=4.06u PD=4.06u
M$22020 AVDD|anode|cathode|pad|vdd \$128987 i|z$6 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$22024 AVDD|anode|cathode|pad|vdd \$128989 \$128990 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22025 \$128988 i|z$38 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22026 \$128989 \$128988 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22027 AVDD|anode|cathode|pad|vdd \$128990 i|z$27 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22028 AVDD|anode|cathode|pad|vdd \$129730 i|z$32 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22030 AVDD|anode|cathode|pad|vdd i|z$42 \$129730 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22031 AVDD|anode|cathode|pad|vdd i|z$43 \$128992 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22033 AVDD|anode|cathode|pad|vdd \$128992 a2|z$4 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$22037 AVDD|anode|cathode|pad|vdd \$128995 \$128996 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22038 \$128994 i|z|zn$8 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22039 \$128995 \$128994 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22040 AVDD|anode|cathode|pad|vdd \$128996 i|z$33 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22041 AVDD|anode|cathode|pad|vdd \$128999 \$129000 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22042 \$128998 i|z$39 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22043 \$128999 \$128998 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22044 AVDD|anode|cathode|pad|vdd \$129000 i|z$34 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22045 AVDD|anode|cathode|pad|vdd \$129733 i|z$35 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22047 AVDD|anode|cathode|pad|vdd i|z$44 \$129733 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22048 AVDD|anode|cathode|pad|vdd i|z$45 \$129003 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22054 AVDD|anode|cathode|pad|vdd \$129003 z$9 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22070 AVDD|anode|cathode|pad|vdd i|z$46 \$129004 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22076 AVDD|anode|cathode|pad|vdd \$129004 z AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22092 AVDD|anode|cathode|pad|vdd i|z|zn$1 \$129005 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=3.205u AS=1.569325p AD=1.389325p PS=7.59u PD=6.09u
M$22095 AVDD|anode|cathode|pad|vdd \$129005 i|z$36 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=3.984p AD=4.164p PS=16.24u PD=17.74u
M$22103 AVDD|anode|cathode|pad|vdd i|z$5 \$129007 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22109 AVDD|anode|cathode|pad|vdd \$129007 a1|z$11 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22125 AVDD|anode|cathode|pad|vdd i|z$48 \$129009 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22131 AVDD|anode|cathode|pad|vdd \$129009 z$13 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22147 AVDD|anode|cathode|pad|vdd \$129011 \$129012 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22148 \$129010 i|z$24 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22149 \$129011 \$129010 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22150 AVDD|anode|cathode|pad|vdd \$129012 i|z$29 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22151 i|z|zn$2 i|zn$8 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22159 AVDD|anode|cathode|pad|vdd i|z$49 \$129013 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22165 AVDD|anode|cathode|pad|vdd \$129013 z$14 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22181 AVDD|anode|cathode|pad|vdd \$129015 \$129016 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22182 \$129014 a2|i|z AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22183 \$129015 \$129014 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22184 AVDD|anode|cathode|pad|vdd \$129016 i|z$2 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22185 AVDD|anode|cathode|pad|vdd \$129018 \$129019 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22186 \$129017 i|z$113 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22187 \$129018 \$129017 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22188 AVDD|anode|cathode|pad|vdd \$129019 i|z$28 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22189 z$6 \$129970 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22190 i|zn$6 i|z|zn$6 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22198 i|z|zn$5 i|zn$3 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22206 i|zn$7 i|zn$2 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22214 AVDD|anode|cathode|pad|vdd \$129023 \$129024 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22215 \$129022 i|z$60 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22216 \$129023 \$129022 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22217 AVDD|anode|cathode|pad|vdd \$129024 i|z$37 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22218 AVDD|anode|cathode|pad|vdd \$129740 i|z$7 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22220 AVDD|anode|cathode|pad|vdd i|z$13 \$129740 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22221 AVDD|anode|cathode|pad|vdd RESULT[3]|c2p|core|i|q \$129026
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p
+ AD=2.8813375p PS=12.07u PD=12.18u
M$22227 AVDD|anode|cathode|pad|vdd \$129026 i|z|zn$7 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22243 a2|zn a1|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22244 VDD|pad|pin1|supply|vdd a1|a2|a3|z a2|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$22245 a2|zn a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22246 \$128890 cp|i|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.339p AD=0.4185p PS=2.33u PD=2.03u
M$22247 VDD|pad|pin1|supply|vdd \$128890 cp|z$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$22248 \$131483 a2$1 a1|c|i|zn AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$22252 AVDD|anode|cathode|pad|vdd a1|z$11 \$131483 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$22256 AVDD|anode|cathode|pad|vdd a2|b|z a1|c|i|zn AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=21.6u AS=9.144p AD=9.144p PS=38.04u PD=38.04u
M$22260 AVDD|anode|cathode|pad|vdd a1|c|i|zn$1 a1|c|i|zn
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=21.6u AS=8.964p AD=9.684p
+ PS=36.54u PD=42.54u
M$22264 \$131484 a2$1 a1|c|i|zn AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$22268 AVDD|anode|cathode|pad|vdd a1|z$11 \$131484 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$22280 \$131485 a2$1 a1|c|i|zn AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$22284 AVDD|anode|cathode|pad|vdd a1|z$11 \$131485 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$22296 \$131486 a2$1 a1|c|i|zn AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$22300 AVDD|anode|cathode|pad|vdd a1|z$11 \$131486 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$22312 AVDD|anode|cathode|pad|vdd a2|b|z a1|c|i|zn$1
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=21.6u AS=9.144p AD=9.144p
+ PS=38.04u PD=38.04u
M$22313 a1|c|i|zn$1 a1|c|i|zn AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=21.6u AS=8.964p AD=9.684p
+ PS=36.54u PD=42.54u
M$22316 AVDD|anode|cathode|pad|vdd \$130779 z$22 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22318 AVDD|anode|cathode|pad|vdd i|z$53 \$130779 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22319 \$130338 i|z$32 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22320 AVDD|anode|cathode|pad|vdd \$130277 \$130339 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22321 \$130277 \$130338 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22322 AVDD|anode|cathode|pad|vdd \$130339 i|z$26 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22323 \$130340 i|z$40 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22329 AVDD|anode|cathode|pad|vdd \$130340 z$23 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22345 \$130342 i|zn$11 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22346 AVDD|anode|cathode|pad|vdd \$130278 \$130343 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22347 \$130278 \$130342 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22348 AVDD|anode|cathode|pad|vdd \$130343 i|z$56 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22349 i|zn$8 i|z|zn$2 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22357 \$130346 i|z$47 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22363 AVDD|anode|cathode|pad|vdd \$130346 z$16 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22379 \$130347 i|z$52 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22380 AVDD|anode|cathode|pad|vdd \$130279 \$130348 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22381 \$130279 \$130347 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22382 AVDD|anode|cathode|pad|vdd \$130348 i|z$57 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22383 \$130350 i|z$36 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22389 AVDD|anode|cathode|pad|vdd \$130350 z$1 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22405 \$130351 i|z$35 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22406 AVDD|anode|cathode|pad|vdd \$130280 \$130352 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22407 \$130280 \$130351 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22408 AVDD|anode|cathode|pad|vdd \$130352 i|z$51 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22409 \$130353 i|z$54 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22410 AVDD|anode|cathode|pad|vdd \$130282 \$130354 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22411 \$130282 \$130353 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22412 AVDD|anode|cathode|pad|vdd \$130354 i|z$58 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22413 \$131062 VALID|a3|c2p|core|i|z AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=3.984p
+ PS=17.74u PD=16.24u
M$22421 \$131062 a2|i|z \$131488 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=9.6u AS=3.984p AD=4.164p PS=16.24u PD=17.74u
M$22429 \$131488 SAMPLE|a1|c2p|core|i|z i|zn$9 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22437 a1|i|z|zn i|zn AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=7.2u AS=3.168p AD=3.168p PS=13.68u PD=13.68u
M$22443 z$17 \$130283 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22444 i|zn$10 i|z|zn$7 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22452 \$130358 i|z|zn$2 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22453 AVDD|anode|cathode|pad|vdd \$130284 \$130359 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22454 \$130284 \$130358 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22455 AVDD|anode|cathode|pad|vdd \$130359 i|z$42 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22456 AVDD|anode|cathode|pad|vdd \$130780 i|z$59 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22458 AVDD|anode|cathode|pad|vdd i|z$34 \$130780 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22459 AVDD|anode|cathode|pad|vdd \$130781 i|z$60 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22461 AVDD|anode|cathode|pad|vdd i|z$1 \$130781 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22462 AVDD|anode|cathode|pad|vdd \$130782 i|z$49 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22464 AVDD|anode|cathode|pad|vdd i|z$58 \$130782 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22465 \$130362 i|z|zn$6 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22466 AVDD|anode|cathode|pad|vdd \$130285 \$130363 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22467 \$130285 \$130362 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22468 AVDD|anode|cathode|pad|vdd \$130363 i|z$114 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22469 \$130364 i|z$55 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22470 AVDD|anode|cathode|pad|vdd \$130287 \$130365 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22471 \$130287 \$130364 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22472 AVDD|anode|cathode|pad|vdd \$130365 i|z AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22473 \$130824 \$130824 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22474 \$130366 i|z$41 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22475 AVDD|anode|cathode|pad|vdd \$130288 \$130367 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22476 \$130288 \$130366 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22477 AVDD|anode|cathode|pad|vdd \$130367 i|z$61 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22478 \$130369 i|zn$9 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=3.205u AS=1.569325p AD=1.389325p PS=7.59u PD=6.09u
M$22481 AVDD|anode|cathode|pad|vdd \$130369 i|z$23 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=3.984p AD=4.164p PS=16.24u PD=17.74u
M$22489 AVDD|anode|cathode|pad|vdd \$130783 i|z$55 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22491 AVDD|anode|cathode|pad|vdd i|z$37 \$130783 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22492 i|zn$2 SAMPLE|a1|c2p|core|i|z AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p
+ PS=17.74u PD=17.74u
M$22500 AVDD|anode|cathode|pad|vdd i|z$11 \$130370 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22502 AVDD|anode|cathode|pad|vdd \$130370 i|z$18 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$22506 \$130371 i|z$25 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22512 AVDD|anode|cathode|pad|vdd \$130371 a2|i|z AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22528 VDD|pad|pin1|supply|vdd CLK|core|i|p2c \$130289 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$22529 VDD|pad|pin1|supply|vdd \$130289 i|z$62 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$22530 VDD|pad|pin1|supply|vdd i|z$62 \$130290 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$22531 VDD|pad|pin1|supply|vdd \$130290 i|z$30 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$22532 a2|z$1 \$130373 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22533 VDD|pad|pin1|supply|vdd b|q \$131489 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$22534 \$131489 a1|b|i|q$2 \$130373 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$22535 \$130373 a2|zn$5 \$131489 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22536 \$130374 \$130291 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22537 VDD|pad|pin1|supply|vdd cp|z$2 \$130291 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22538 RESULT[2]|c2p|core|i|q \$130375 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$22539 a2$1 z$7 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=3.6u
+ AS=2.034p AD=2.034p PS=13.98u PD=13.98u
M$22540 a2 z$4 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.8u
+ AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$22542 a2$1 z$4 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.8u
+ AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$22551 \$131967 a2 a1|c|i|zn$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$22555 AVDD|anode|cathode|pad|vdd a1|z$11 \$131967 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$22567 \$131969 a2 a1|c|i|zn$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$22571 AVDD|anode|cathode|pad|vdd a1|z$11 \$131969 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$22583 \$131970 a2 a1|c|i|zn$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$22587 AVDD|anode|cathode|pad|vdd a1|z$11 \$131970 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$22599 \$131971 a2 a1|c|i|zn$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$22603 AVDD|anode|cathode|pad|vdd a1|z$11 \$131971 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$22619 AVDD|anode|cathode|pad|vdd a1|c|i|zn$1 \$130275
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.36u AS=0.2129625p
+ AD=0.2034p PS=1.415u PD=1.85u
M$22620 AVDD|anode|cathode|pad|vdd \$130275 i|z$53 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.585u AS=0.2129625p AD=0.330525p PS=1.415u PD=2.3u
M$22621 \$131962 a1|c|i|zn AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.36u AS=0.2034p
+ AD=0.2129625p PS=1.85u PD=1.415u
M$22622 AVDD|anode|cathode|pad|vdd \$131962 i|z$65 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.585u AS=0.2129625p AD=0.330525p PS=1.415u PD=2.3u
M$22623 AVDD|anode|cathode|pad|vdd \$132660 a2|a3|z AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22625 AVDD|anode|cathode|pad|vdd i|z$65 \$132660 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22626 AVDD|anode|cathode|pad|vdd a2|z$4 \$131972 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22627 \$131972 a1|i|z|zn AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u AS=0.996p AD=0.996p
+ PS=4.06u PD=4.06u
M$22630 AVDD|anode|cathode|pad|vdd \$131972 i|z$66 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$22634 AVDD|anode|cathode|pad|vdd i|z$74 \$131974 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22640 AVDD|anode|cathode|pad|vdd \$131974 z$11 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22656 z$24 \$132944 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22657 i|z|zn$7 i|zn$10 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22665 AVDD|anode|cathode|pad|vdd i|z$75 \$131975 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22671 AVDD|anode|cathode|pad|vdd \$131975 z$25 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22687 AVDD|anode|cathode|pad|vdd i|z|zn \$131977 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=3.205u AS=1.569325p AD=1.389325p PS=7.59u PD=6.09u
M$22690 AVDD|anode|cathode|pad|vdd \$131977 i|z$67 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=3.984p AD=4.164p PS=16.24u PD=17.74u
M$22698 AVDD|anode|cathode|pad|vdd \$131980 \$131981 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22699 \$131979 i|z|zn$4 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22700 \$131980 \$131979 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22701 AVDD|anode|cathode|pad|vdd \$131981 i|z$63 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22702 AVDD|anode|cathode|pad|vdd i|z$76 \$131982 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22708 AVDD|anode|cathode|pad|vdd \$131982 z$10 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22724 AVDD|anode|cathode|pad|vdd i|z$59 \$131983 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22730 AVDD|anode|cathode|pad|vdd \$131983 z$19 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22746 AVDD|anode|cathode|pad|vdd \$132664 i|z$74 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22748 AVDD|anode|cathode|pad|vdd i|z$101 \$132664 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22749 AVDD|anode|cathode|pad|vdd \$131985 \$131986 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22750 \$131984 i|zn$10 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22751 \$131985 \$131984 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22752 AVDD|anode|cathode|pad|vdd \$131986 i|z$68 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22753 i|zn$11 i|z|zn$8 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22761 z$2 \$132946 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22762 AVDD|anode|cathode|pad|vdd b|i|q \$131989 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22768 AVDD|anode|cathode|pad|vdd \$131989 i|z|zn$8 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22784 AVDD|anode|cathode|pad|vdd \$132668 i|z$69 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22786 AVDD|anode|cathode|pad|vdd i|z$77 \$132668 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22787 AVDD|anode|cathode|pad|vdd \$131992 \$131993 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22788 \$131991 i|z$72 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22789 \$131992 \$131991 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22790 AVDD|anode|cathode|pad|vdd \$131993 i|z$64 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22791 AVDD|anode|cathode|pad|vdd \$131995 \$131996 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22792 \$131994 i|z$69 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22793 \$131995 \$131994 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22794 AVDD|anode|cathode|pad|vdd \$131996 i|z$70 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22795 AVDD|anode|cathode|pad|vdd \$132670 i|z$46 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22797 AVDD|anode|cathode|pad|vdd i|z$79 \$132670 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22798 AVDD|anode|cathode|pad|vdd \$131999 \$132000 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22799 \$131998 i|z$103 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22800 \$131999 \$131998 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22801 AVDD|anode|cathode|pad|vdd \$132000 i|z$111 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22802 AVDD|anode|cathode|pad|vdd \$132002 \$132003 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22803 \$132001 i|z$73 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22804 \$132002 \$132001 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22805 AVDD|anode|cathode|pad|vdd \$132003 i|z$71 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22806 AVDD|anode|cathode|pad|vdd \$132671 i|z$16 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22808 AVDD|anode|cathode|pad|vdd i|z$80 \$132671 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22809 AVDD|anode|cathode|pad|vdd b|i|q$1 \$132005 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22815 AVDD|anode|cathode|pad|vdd \$132005 i|z|zn$9 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22831 \$132007 \$131965 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22832 VDD|pad|pin1|supply|vdd cp|z$1 \$131965 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22833 \$131966 \$131965 \$132213 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22834 \$132213 \$132008 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$22835 \$132948 \$132007 \$132215 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$22836 \$132215 \$132009 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$22837 \$132223 d|zn$4 \$131966 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$22838 VDD|pad|pin1|supply|vdd \$131966 \$132008 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$22839 VDD|pad|pin1|supply|vdd \$132007 \$132223 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$22840 \$132008 \$131965 \$132948 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$22841 VDD|pad|pin1|supply|vdd \$132948 \$132009 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$22842 a1|i|q$1 \$132009 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22843 VDD|pad|pin1|supply|vdd \$130374 \$131585 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$22844 \$131585 d|zn$3 \$130292 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$22845 \$130292 \$130291 \$131586 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22846 VDD|pad|pin1|supply|vdd \$130293 \$131586 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22847 \$130293 \$130292 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$22848 \$130293 \$130291 \$130294 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$22849 \$130294 \$130374 \$131582 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$22850 VDD|pad|pin1|supply|vdd \$130375 \$131582 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$22851 VDD|pad|pin1|supply|vdd \$130294 \$130375 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$22852 AVDD|anode|cathode|pad|vdd i|zn$1 \$134936 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22858 AVDD|anode|cathode|pad|vdd \$134936 z$3 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22874 z$26 \$133281 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22875 \$133696 \$133696 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22876 i|z|zn i|zn$5 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22884 \$133345 i|z$66 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22890 AVDD|anode|cathode|pad|vdd \$133345 a2|b|z AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22906 \$133697 \$133697 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22907 AVDD|anode|cathode|pad|vdd \$134938 \$134875 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22908 \$134937 i|z$9 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22909 \$133346 i|z$83 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22910 AVDD|anode|cathode|pad|vdd \$133283 \$133347 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22911 \$134938 \$134937 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22912 AVDD|anode|cathode|pad|vdd \$134875 i|z$87 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22913 \$133283 \$133346 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22914 AVDD|anode|cathode|pad|vdd \$133347 i|z$86 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22915 AVDD|anode|cathode|pad|vdd \$135839 i|z$50 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22917 AVDD|anode|cathode|pad|vdd i|z$57 \$135839 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22918 \$133349 i|zn$7 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=3.205u AS=1.569325p AD=1.389325p PS=7.59u PD=6.09u
M$22921 AVDD|anode|cathode|pad|vdd \$133349 a1|z$12 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=3.984p AD=4.164p PS=16.24u PD=17.74u
M$22929 AVDD|anode|cathode|pad|vdd \$133351 i|z$83 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22931 AVDD|anode|cathode|pad|vdd i|z$87 \$133351 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22932 AVDD|anode|cathode|pad|vdd \$133353 i|z$88 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22934 AVDD|anode|cathode|pad|vdd i|z$102 \$133353 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22935 \$133355 a1|i|z|zn AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p
+ PS=3.53u PD=2.03u
M$22936 AVDD|anode|cathode|pad|vdd \$133284 \$133356 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22937 \$134939 \$134939 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22938 \$133284 \$133355 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22939 AVDD|anode|cathode|pad|vdd \$133356 i|z$43 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22940 AVDD|anode|cathode|pad|vdd i|zn$1 \$134940 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22946 AVDD|anode|cathode|pad|vdd \$134940 z$3 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22962 \$133358 i|z$89 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22968 AVDD|anode|cathode|pad|vdd \$133358 z$8 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22984 AVDD|anode|cathode|pad|vdd \$135840 i|z$22 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22986 AVDD|anode|cathode|pad|vdd i|z$86 \$135840 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22987 \$133359 i|z$84 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22988 AVDD|anode|cathode|pad|vdd \$133286 \$133360 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22989 AVDD|anode|cathode|pad|vdd \$134942 \$134876 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22990 \$134941 i|z|zn$9 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22991 \$133286 \$133359 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22992 AVDD|anode|cathode|pad|vdd \$133360 i|z$80 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22993 \$134942 \$134941 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22994 AVDD|anode|cathode|pad|vdd \$134876 i|z$99 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22995 \$133361 i|zn$3 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22996 AVDD|anode|cathode|pad|vdd \$133287 \$133362 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22997 \$133287 \$133361 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22998 AVDD|anode|cathode|pad|vdd \$133362 i|z$90 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22999 AVDD|anode|cathode|pad|vdd b|i|q$3 \$134943 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$23005 AVDD|anode|cathode|pad|vdd \$134943 i|z|zn$3 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$23021 AVDD|anode|cathode|pad|vdd \$133364 i|z$82 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23023 AVDD|anode|cathode|pad|vdd i|z$91 \$133364 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23024 i|zn$12 i|z|zn$4 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$23032 AVDD|anode|cathode|pad|vdd i|z$31 \$133367 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23034 AVDD|anode|cathode|pad|vdd \$133367 a2|z$5 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$23038 AVDD|anode|cathode|pad|vdd \$134945 \$134877 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23039 \$134944 i|z$20 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23040 \$134945 \$134944 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23041 AVDD|anode|cathode|pad|vdd \$134877 i|z$105 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23042 AVDD|anode|cathode|pad|vdd \$134949 \$134878 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23043 \$134947 i|z$106 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23044 i|zn a1|i|z|zn AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=7.2u AS=3.168p AD=3.168p PS=13.68u PD=13.68u
M$23050 \$134949 \$134947 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23051 AVDD|anode|cathode|pad|vdd \$134878 i|z$101 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23052 AVDD|anode|cathode|pad|vdd \$133368 i|z$17 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23054 AVDD|anode|cathode|pad|vdd i|z$81 \$133368 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23055 \$133369 i|z$50 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23056 AVDD|anode|cathode|pad|vdd \$133288 \$133370 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23057 AVDD|anode|cathode|pad|vdd \$135841 i|z$103 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23059 AVDD|anode|cathode|pad|vdd i|z$56 \$135841 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23060 \$133288 \$133369 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23061 AVDD|anode|cathode|pad|vdd \$133370 i|z$79 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23062 z$27 \$136067 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$23063 \$133371 i|z$88 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$23069 AVDD|anode|cathode|pad|vdd \$133371 z$18 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$23085 AVDD|anode|cathode|pad|vdd \$135842 i|z$38 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23087 AVDD|anode|cathode|pad|vdd i|z$90 \$135842 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23088 i|zn$13 i|z|zn$9 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$23096 AVDD|anode|cathode|pad|vdd \$135843 i|z$107 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23098 AVDD|anode|cathode|pad|vdd i|z$97 \$135843 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23099 \$134951 \$134951 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$23100 AVDD|anode|cathode|pad|vdd \$133372 i|z$39 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23102 AVDD|anode|cathode|pad|vdd i|z$19 \$133372 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23103 AVDD|anode|cathode|pad|vdd \$133373 i|z$41 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23105 AVDD|anode|cathode|pad|vdd i|z$33 \$133373 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23106 AVDD|anode|cathode|pad|vdd \$134954 \$134879 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23107 \$134952 i|z$108 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23108 \$134954 \$134952 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23109 AVDD|anode|cathode|pad|vdd \$134879 i|z$92 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23110 \$133374 i|z$78 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$23116 AVDD|anode|cathode|pad|vdd \$133374 z$5 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$23132 AVDD|anode|cathode|pad|vdd \$134957 \$134880 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23133 \$134955 i|z$109 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23134 \$134957 \$134955 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23135 AVDD|anode|cathode|pad|vdd \$134880 i|z$77 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23136 i|z|zn$4 i|zn$12 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$23144 AVDD|anode|cathode|pad|vdd \$135844 i|z$110 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23146 AVDD|anode|cathode|pad|vdd i|z$104 \$135844 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23147 AVDD|anode|cathode|pad|vdd \$133376 i|z$45 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23149 AVDD|anode|cathode|pad|vdd i|z$93 \$133376 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23150 i|z|zn$8 i|zn$11 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$23158 AVDD|anode|cathode|pad|vdd \$133378 i|z$94 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23160 AVDD|anode|cathode|pad|vdd i|z$95 \$133378 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23161 AVDD|anode|cathode|pad|vdd \$135845 i|z$73 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23163 AVDD|anode|cathode|pad|vdd i|z$68 \$135845 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23164 AVDD|anode|cathode|pad|vdd \$133381 i|z$89 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23166 AVDD|anode|cathode|pad|vdd i|z$92 \$133381 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23167 \$133383 b|i|q$2 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$23173 AVDD|anode|cathode|pad|vdd \$133383 i|z|zn$6 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$23189 AVDD|anode|cathode|pad|vdd \$135846 i|z$108 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23191 AVDD|anode|cathode|pad|vdd i|z$64 \$135846 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23192 AVDD|anode|cathode|pad|vdd \$134960 \$134881 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23193 \$134959 i|z$110 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23194 \$134960 \$134959 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23195 AVDD|anode|cathode|pad|vdd \$134881 i|z$95 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23196 AVDD|anode|cathode|pad|vdd \$134962 \$134882 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23197 \$134961 i|z$94 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23198 \$134962 \$134961 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23199 AVDD|anode|cathode|pad|vdd \$134882 i|z$93 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23200 AVDD|anode|cathode|pad|vdd \$135847 i|z$84 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23202 AVDD|anode|cathode|pad|vdd i|z$61 \$135847 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23203 \$133384 i|z|zn$7 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23204 AVDD|anode|cathode|pad|vdd \$133289 \$133385 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23205 \$133289 \$133384 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23206 AVDD|anode|cathode|pad|vdd \$133385 i|z$91 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23207 AVDD|anode|cathode|pad|vdd \$135848 i|z$40 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23209 AVDD|anode|cathode|pad|vdd i|z$105 \$135848 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23210 \$133386 i|z$85 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23211 AVDD|anode|cathode|pad|vdd \$133291 \$133387 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23212 AVDD|anode|cathode|pad|vdd \$135849 i|z$76 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23214 AVDD|anode|cathode|pad|vdd i|z$96 \$135849 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23215 \$133291 \$133386 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23216 AVDD|anode|cathode|pad|vdd \$133387 i|z$96 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23217 AVDD|anode|cathode|pad|vdd \$133389 i|z$47 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23219 AVDD|anode|cathode|pad|vdd i|z$70 \$133389 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23220 \$133390 i|z$82 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23221 AVDD|anode|cathode|pad|vdd \$133292 \$133391 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23222 \$133292 \$133390 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23223 AVDD|anode|cathode|pad|vdd \$133391 i|z$97 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23224 AVDD|anode|cathode|pad|vdd \$134964 \$134883 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23225 \$134963 i|z$21 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23226 AVDD|anode|cathode|pad|vdd \$133393 i|z$85 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23228 AVDD|anode|cathode|pad|vdd i|z$71 \$133393 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23229 \$134964 \$134963 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23230 AVDD|anode|cathode|pad|vdd \$134883 i|z$102 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23231 AVDD|anode|cathode|pad|vdd \$134966 \$134884 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23232 \$134965 i|z$112 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23233 i|z|zn$9 i|zn$13 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$23241 \$134966 \$134965 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23242 AVDD|anode|cathode|pad|vdd \$134884 i|z$44 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23243 AVDD|anode|cathode|pad|vdd \$135850 i|z$48 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23245 AVDD|anode|cathode|pad|vdd i|z$100 \$135850 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23246 \$133395 i|z$107 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23247 AVDD|anode|cathode|pad|vdd \$133293 \$133396 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23248 AVDD|anode|cathode|pad|vdd \$134968 \$134885 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23249 \$134967 i|zn$13 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23250 \$133293 \$133395 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23251 AVDD|anode|cathode|pad|vdd \$133396 i|z$100 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23252 \$134968 \$134967 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23253 AVDD|anode|cathode|pad|vdd \$134885 i|z$104 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23254 \$133397 i|zn$12 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23255 AVDD|anode|cathode|pad|vdd \$133294 \$133398 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23256 \$133294 \$133397 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23257 AVDD|anode|cathode|pad|vdd \$133398 i|z$98 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23258 AVDD|anode|cathode|pad|vdd \$133401 i|z$52 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23260 AVDD|anode|cathode|pad|vdd i|z$99 \$133401 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23261 AVDD|anode|cathode|pad|vdd \$135851 i|z$78 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23263 AVDD|anode|cathode|pad|vdd i|z$51 \$135851 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23264 AVDD|anode|cathode|pad|vdd \$133402 i|z$72 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23266 AVDD|anode|cathode|pad|vdd i|z$98 \$133402 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23267 \$134969 \$134735 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23268 VDD|pad|pin1|supply|vdd cp|z$2 \$134735 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23269 \$134736 \$134735 \$134922 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$23270 \$134922 \$134886 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$23271 \$136070 \$134969 \$134923 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$23272 \$134923 \$134970 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$23273 \$135763 d|zn$6 \$134736 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$23274 VDD|pad|pin1|supply|vdd \$134736 \$134886 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$23275 VDD|pad|pin1|supply|vdd \$134969 \$135763 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$23276 \$134886 \$134735 \$136070 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$23277 VDD|pad|pin1|supply|vdd \$136070 \$134970 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$23278 VDD|pad|pin1|supply|vdd a2|a3|zn \$134676 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23279 \$134676 RST|a1|b|cdn|core|i|p2c b|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$23280 b|zn$4 a1|b|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23281 VDD|pad|pin1|supply|vdd i|z$4 \$133305 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$23282 VDD|pad|pin1|supply|vdd \$133305 cp|i|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$23283 a1|b|i|q$2 \$134970 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$23284 \$134887 a2|zn$6 d|zn$2 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23285 d|zn$2 a1|z$13 \$134887 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$23286 \$134887 b|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23287 \$139964 \$140018 \$139964 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23299 \$137099 \$137099 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$23300 \$136386 i|zn$4 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$23301 AVDD|anode|cathode|pad|vdd \$136342 \$136387 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$23302 \$136342 \$136386 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23303 AVDD|anode|cathode|pad|vdd \$136387 i|z$14 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23304 \$136388 i|zn$5 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$23310 AVDD|anode|cathode|pad|vdd \$136388 z$7 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$23350 \$139965 \$140019 \$139965 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23386 \$139966 \$140020 \$139966 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23422 \$136389 i|z$67 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$23428 AVDD|anode|cathode|pad|vdd \$136389 z$4 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$23444 \$139967 \$140021 \$139967 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23468 AVDD|anode|cathode|pad|vdd \$136706 i|z$113 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23470 AVDD|anode|cathode|pad|vdd i|z$114 \$136706 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23483 \$139968 \$140022 \$139968 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23519 \$139969 \$140023 \$139969 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23543 AVDD|anode|cathode|pad|vdd \$136708 i|z$54 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23545 AVDD|anode|cathode|pad|vdd i|z$111 \$136708 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23558 \$139970 \$140024 \$139970 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23594 \$139971 \$140025 \$139971 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23630 AVDD|anode|cathode|pad|vdd \$136709 i|z$112 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$23632 AVDD|anode|cathode|pad|vdd i|z$63 \$136709 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23633 \$139972 \$140026 \$139972 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23669 \$139973 \$140027 \$139973 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23705 \$136391 \$136343 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23706 VDD|pad|pin1|supply|vdd cp|i|z \$136343 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23707 VDD|pad|pin1|supply|vdd \$136391 \$138029 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$23708 \$138029 d|zn$9 \$136344 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$23709 \$136344 \$136343 \$138008 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$23710 VDD|pad|pin1|supply|vdd \$136392 \$138008 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$23711 \$136392 \$136344 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$23712 \$136392 \$136343 \$136345 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$23713 \$136345 \$136391 \$138011 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$23714 VDD|pad|pin1|supply|vdd \$136393 \$138011 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$23715 VDD|pad|pin1|supply|vdd \$136345 \$136393 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$23716 a1|b|i|q$1 \$136393 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$23717 \$136394 \$136346 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23718 VDD|pad|pin1|supply|vdd cp|z$3 \$136346 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23719 VDD|pad|pin1|supply|vdd a1|z$3 \$140028 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23720 \$140028 a2|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$23721 VDD|pad|pin1|supply|vdd \$140028 d|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23722 a2|zn$6 a1|b|i|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23723 VDD|pad|pin1|supply|vdd a1|a2|a3|z a2|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$23724 a2|zn$6 a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23725 VDD|pad|pin1|supply|vdd \$136394 \$138006 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$23726 \$138006 d|zn$10 \$136347 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$23727 \$136347 \$136346 \$137985 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$23728 VDD|pad|pin1|supply|vdd \$136395 \$137985 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$23729 \$136395 \$136347 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$23730 \$136395 \$136346 \$136348 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$23731 \$136348 \$136394 \$137991 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$23732 VDD|pad|pin1|supply|vdd \$136396 \$137991 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$23733 VDD|pad|pin1|supply|vdd \$136348 \$136396 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$23734 a1|b|i|q \$136396 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$24095 \$141594 \$141285 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$24096 VDD|pad|pin1|supply|vdd cp|z$3 \$141285 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$24097 \$141286 \$141285 \$141943 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$24098 \$141943 \$141595 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$24099 \$142757 \$141594 \$141945 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$24100 \$141945 \$141596 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$24101 \$141952 d|zn$5 \$141286 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$24102 VDD|pad|pin1|supply|vdd \$141286 \$141595 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$24103 VDD|pad|pin1|supply|vdd \$141594 \$141952 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$24104 \$141595 \$141285 \$142757 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$24105 VDD|pad|pin1|supply|vdd \$142757 \$141596 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$24106 a2|i|q \$141596 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$24107 a2|z \$141598 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$24108 VDD|pad|pin1|supply|vdd b|i|q \$141597 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$24109 \$141597 a1|b|i|q \$141598 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$24110 \$141598 a2|zn$5 \$141597 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$24111 \$145293 \$145605 \$145293 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$24123 \$140018 z$26 \$143069 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24124 \$143069 zn$3 \$143069 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24126 \$140018 zn$3 \$140018 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24139 \$143070 z$26 \$140018 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24142 \$143070 zn$3 \$143070 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24155 \$143071 z$26 \$140018 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24158 \$143071 zn$3 \$143071 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24159 \$145294 \$145606 \$145294 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=1382.4u AS=590.976p AD=590.976p PS=2482.56u PD=2482.56u
M$24171 \$140019 z$26 \$143072 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24172 \$143072 zn$3 \$143072 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24174 \$140019 zn$3 \$140019 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24187 \$143073 z$26 \$140019 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24190 \$143073 zn$3 \$143073 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24203 \$143074 z$26 \$140019 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24206 \$143074 zn$3 \$143074 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24207 \$145295 \$145607 \$145295 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=691.2u AS=295.488p AD=295.488p PS=1241.28u PD=1241.28u
M$24219 \$140020 z$26 \$143075 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24220 \$143075 zn$3 \$143075 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24222 \$140020 zn$3 \$140020 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24235 \$143076 z$26 \$140020 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24238 \$143076 zn$3 \$143076 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24251 \$143077 z$26 \$140020 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24254 \$143077 zn$3 \$143077 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24255 \$145296 \$145608 \$145296 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=172.8u AS=73.872p AD=73.872p PS=310.32u PD=310.32u
M$24267 \$140021 z$26 \$143078 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24268 \$143078 zn$3 \$143078 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24270 \$140021 zn$3 \$140021 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24283 \$143079 z$26 \$140021 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24286 \$143079 zn$3 \$143079 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24299 \$143080 z$26 \$140021 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24302 \$143080 zn$3 \$143080 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24303 \$145297 \$145609 \$145297 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$24315 \$140022 z$26 \$143081 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24316 \$143081 zn$3 \$143081 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24318 \$140022 zn$3 \$140022 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24331 \$143082 z$26 \$140022 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24334 \$143082 zn$3 \$143082 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24347 \$143083 z$26 \$140022 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24350 \$143083 zn$3 \$143083 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24351 \$145298 \$145610 \$145298 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$24363 \$140023 z$26 \$143084 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24364 \$143084 zn$3 \$143084 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24366 \$140023 zn$3 \$140023 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24379 \$143085 z$26 \$140023 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24382 \$143085 zn$3 \$143085 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24395 \$143086 z$26 \$140023 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24398 \$143086 zn$3 \$143086 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24411 \$140024 z$26 \$143087 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24412 \$143087 zn$3 \$143087 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24414 \$140024 zn$3 \$140024 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24427 \$143088 z$26 \$140024 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24430 \$143088 zn$3 \$143088 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24443 \$143089 z$26 \$140024 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24446 \$143089 zn$3 \$143089 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24459 \$140025 z$26 \$143090 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24460 \$143090 zn$3 \$143090 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24462 \$140025 zn$3 \$140025 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24475 \$143091 z$26 \$140025 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24478 \$143091 zn$3 \$143091 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24491 \$143092 z$26 \$140025 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24494 \$143092 zn$3 \$143092 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24507 \$140026 z$26 \$143093 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24508 \$143093 zn$3 \$143093 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24510 \$140026 zn$3 \$140026 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24523 \$143094 z$26 \$140026 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24526 \$143094 zn$3 \$143094 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24539 \$143095 z$26 \$140026 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24542 \$143095 zn$3 \$143095 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24543 \$145299 \$145611 \$145299 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$24555 \$140027 z$26 \$143096 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24556 \$143096 zn$3 \$143096 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24558 \$140027 zn$3 \$140027 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24571 \$143097 z$26 \$140027 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24574 \$143097 zn$3 \$143097 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24587 \$143098 z$26 \$140027 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24590 \$143098 zn$3 \$143098 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24591 \$145049 \$144246 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$24592 VDD|pad|pin1|supply|vdd cp|z$3 \$144246 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$24593 \$144248 \$144246 \$144892 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$24594 \$144892 \$144249 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$24595 \$145612 \$145049 \$144908 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$24596 \$144908 \$145050 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$24597 \$145290 d|z$4 \$144248 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$24598 VDD|pad|pin1|supply|vdd \$144248 \$144249 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$24599 VDD|pad|pin1|supply|vdd \$145049 \$145290 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$24600 \$144249 \$144246 \$145612 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$24601 VDD|pad|pin1|supply|vdd \$145612 \$145050 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$24602 VDD|pad|pin1|supply|vdd a2|a3|zn \$144167 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$24603 \$144167 RST|a1|b|cdn|core|i|p2c b|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$24604 b|zn$5 a1|b|i|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$24605 b|i|q$2 \$145050 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$24966 \$150121 \$150578 \$150121 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$24978 \$145605 z$26 \$148728 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24979 \$148728 zn$3 \$148728 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24981 \$145605 zn$3 \$145605 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24994 \$148729 z$26 \$145605 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24997 \$148729 zn$3 \$148729 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25010 \$148730 z$26 \$145605 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25013 \$148730 zn$3 \$148730 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25026 \$145606 z$3 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=19.2u AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$25027 a2$1 z$1 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u
+ AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$25029 \$145606 z$1 \$145606 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$25042 VIN|core|padres z$7 \$145606 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=19.2u AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$25043 \$145606 z$4 \$145606 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$25045 VIN|core|padres z$4 VIN|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$25058 VIP|core|padres z$27 \$145606 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=19.2u AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$25059 \$145606 zn$5 \$145606 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$25061 VIP|core|padres zn$5 VIP|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$25074 \$145607 z$7 VREFL|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$25075 VREFL|core|padres z$4 VREFL|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$25077 \$145607 z$4 \$145607 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$25090 a2$1 z$9 \$145607 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$25091 \$145607 z \$145607 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$25093 a2$1 z a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$25106 a2 z$8 \$145607 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u
+ AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$25107 \$145607 z$5 \$145607 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$25109 a2 z$5 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$25110 \$150122 \$150579 \$150122 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=345.6u AS=147.744p AD=147.744p PS=620.64u PD=620.64u
M$25122 \$145608 z$7 VREFL|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$25125 \$145608 z$4 \$145608 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25138 a2$1 z$14 \$145608 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$25139 \$145608 z$15 \$145608 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25141 a2$1 z$15 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25154 a2 z$18 \$145608 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$25155 \$145608 z$19 \$145608 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25157 a2 z$19 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25170 \$145609 z$7 VREFL|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25173 \$145609 z$4 \$145609 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25186 a2$1 z$16 \$145609 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25187 \$145609 z$25 \$145609 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25189 a2$1 z$25 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25202 a2 z$21 \$145609 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25203 \$145609 z$23 \$145609 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25205 a2 z$23 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25218 \$145610 z$7 VREFL|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25221 \$145610 z$4 \$145610 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25234 a2$1 z$24 \$145610 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25235 \$145610 zn$4 \$145610 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25237 a2$1 zn$4 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25250 a2 z$24 \$145610 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25253 a2 zn$4 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25398 \$150123 \$150580 \$150123 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$25410 \$145611 z$26 \$148731 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25411 \$148731 zn$3 \$148731 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25413 \$145611 zn$3 \$145611 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$25426 \$148732 z$26 \$145611 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25429 \$148732 zn$3 \$148732 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25442 \$148733 z$26 \$145611 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25445 \$148733 zn$3 \$148733 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25446 a1|z$3 \$146514 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$25447 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$147109
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p
+ PS=2.03u PD=2.03u
M$25448 \$147109 a1|i|q \$146514 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25449 \$146514 a2|z$2 \$147109 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$25450 a2|z$6 \$149324 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$25451 VDD|pad|pin1|supply|vdd b|i|q$1 \$149869 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25452 \$149869 a1|i|q$1 \$149324 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25453 \$149324 a2|zn$5 \$149869 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$25454 VDD|pad|pin1|supply|vdd a2|zn$3 \$148240 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$25455 \$148240 a1|z$9 d|zn$9 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25456 d|zn$9 b|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$25457 VDD|pad|pin1|supply|vdd a1|z$3 \$150581 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$25458 \$150581 a2|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25459 VDD|pad|pin1|supply|vdd \$150581 d|z$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$25460 VDD|pad|pin1|supply|vdd a1|z$3 \$146314 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$25461 \$146314 a2|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25462 VDD|pad|pin1|supply|vdd \$146314 d|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$25463 VDD|pad|pin1|supply|vdd cp|i|z \$146315 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$25464 VDD|pad|pin1|supply|vdd \$146315 cp|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$25825 \$155172 \$155875 \$155172 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$25837 \$150578 z$26 \$153380 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25838 \$153380 zn$3 \$153380 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25840 \$150578 zn$3 \$150578 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$25853 \$153381 z$26 \$150578 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25856 \$153381 zn$3 \$153381 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25869 \$153382 z$26 \$150578 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25872 \$153382 zn$3 \$153382 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25981 \$150579 z$7 VREFL|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$25984 \$150579 z$4 \$150579 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$25997 a2$1 z$12 \$150579 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$25998 \$150579 z$11 \$150579 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$26000 a2$1 z$11 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$26013 a2 z$10 \$150579 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$26014 \$150579 z$13 \$150579 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$26016 a2 z$13 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$26257 \$155173 \$155876 \$155173 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$26269 \$150580 z$26 \$153383 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26270 \$153383 zn$3 \$153383 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26272 \$150580 zn$3 \$150580 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$26285 \$153384 z$26 \$150580 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26288 \$153384 zn$3 \$153384 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26301 \$153385 z$26 \$150580 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26304 \$153385 zn$3 \$153385 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26305 a1|z$13 RESULT[0]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$26306 a2|z$7 \$155174 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$26307 VDD|pad|pin1|supply|vdd b|i|q$3 \$156094 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$26308 \$156094 a1|b|i|q$3 \$155174 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$26309 \$155174 a2|zn$5 \$156094 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$26310 VDD|pad|pin1|supply|vdd a2|a3|zn \$153081 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$26311 \$153081 RST|a1|b|cdn|core|i|p2c b|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$26312 b|zn$6 a1|b|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$26313 VDD|pad|pin1|supply|vdd a2|zn$3 \$153738 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$26314 \$153738 a1|z$1 d|zn$10 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$26315 d|zn$10 b|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$26316 a1|z RESULT[4]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$26677 a2|zn$1 a1|b|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$26678 VDD|pad|pin1|supply|vdd a1|a2|a3|z a2|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$26679 a2|zn$1 a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$26680 \$160833 \$161529 \$160833 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$26692 \$155875 z$26 \$159177 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26693 \$159177 zn$3 \$159177 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26695 \$155875 zn$3 \$155875 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$26708 \$159178 z$26 \$155875 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26711 \$159178 zn$3 \$159178 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26724 \$159179 z$26 \$155875 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26727 \$159179 zn$3 \$159179 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27112 \$160834 \$161530 \$160834 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27124 \$155876 z$26 \$159180 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27125 \$159180 zn$3 \$159180 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27127 \$155876 zn$3 \$155876 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27140 \$159181 z$26 \$155876 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27143 \$159181 zn$3 \$159181 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27156 \$159182 z$26 \$155876 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27159 \$159182 zn$3 \$159182 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27160 \$158510 \$157993 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$27161 VDD|pad|pin1|supply|vdd cp|z$3 \$157993 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$27162 VDD|pad|pin1|supply|vdd \$158510 \$159281 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$27163 \$159281 a2|d|zn \$157994 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$27164 \$157994 \$157993 \$159282 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$27165 VDD|pad|pin1|supply|vdd \$158244 \$159282 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$27166 \$158244 \$157994 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$27167 \$158244 \$157993 \$157995 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$27168 \$157995 \$158510 \$159279 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$27169 VDD|pad|pin1|supply|vdd \$158511 \$159279 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$27170 VDD|pad|pin1|supply|vdd \$157995 \$158511 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$27171 a2|zn$2 a1|b|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$27172 VDD|pad|pin1|supply|vdd a1|a2|a3|z a2|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$27173 a2|zn$2 a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$27174 a1|i|q \$158511 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$27535 \$162671 a2|zn$4 d|zn$7 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$27536 d|zn$7 a1|z$8 \$162671 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$27537 \$162671 b|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$27538 VDD|pad|pin1|supply|vdd a2|a3|zn \$162768 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$27539 \$162768 RST|a1|b|cdn|core|i|p2c a2|d|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$27540 \$166600 \$167242 \$166600 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27552 \$161529 z$26 \$164854 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27553 \$164854 zn$3 \$164854 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27555 \$161529 zn$3 \$161529 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27568 \$164855 z$26 \$161529 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27571 \$164855 zn$3 \$164855 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27584 \$164856 z$26 \$161529 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27587 \$164856 zn$3 \$164856 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27588 \$166601 \$167243 \$166601 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27636 \$166602 \$167244 \$166602 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27684 \$166603 \$167245 \$166603 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27732 \$166604 \$167246 \$166604 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27780 \$166605 \$167247 \$166605 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27828 \$166606 \$167248 \$166606 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27876 \$166607 \$167249 \$166607 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27924 \$166608 \$167250 \$166608 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27972 \$166609 \$167251 \$166609 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27984 \$161530 z$26 \$164857 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27985 \$164857 zn$3 \$164857 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27987 \$161530 zn$3 \$161530 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28000 \$164858 z$26 \$161530 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28003 \$164858 zn$3 \$164858 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28016 \$164859 z$26 \$161530 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28019 \$164859 zn$3 \$164859 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28020 VDD|pad|pin1|supply|vdd a2|zn$3 \$163558 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$28021 \$163558 a1|z$2 d|zn$8 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$28022 d|zn$8 b|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$28023 VDD|pad|pin1|supply|vdd a2|a3|zn \$165877 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$28024 \$165877 RST|a1|b|cdn|core|i|p2c b|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$28025 b|zn$3 a1|b|i|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$28026 a2|zn$3 a1|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$28027 VDD|pad|pin1|supply|vdd a2|z$2 a2|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$28028 a2|zn$3 a1|a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$28029 a1|z$7 a1|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$28390 \$167242 z$26 \$169906 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28391 \$169906 zn$3 \$169906 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28393 \$167242 zn$3 \$167242 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28394 \$169907 z$26 \$167242 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28397 VDD|pad|pin1|supply|vdd a1|a2|q \$207273 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28398 \$207273 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28399 \$169907 zn$3 \$169907 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28400 d|z$5 \$207273 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28401 \$169908 z$26 \$167242 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28402 \$207275 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28403 VDD|pad|pin1|supply|vdd \$207275 \$207253 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28406 VDD|pad|pin1|supply|vdd \$207253 \$209048 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28407 \$209048 d|z$14 \$207276 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28408 \$207276 \$207275 \$208955 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28409 \$208955 \$207277 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28410 \$169908 zn$3 \$169908 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28411 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$208955
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28412 \$207277 \$207276 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28413 \$207277 \$207275 \$207254 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28414 \$207254 \$207253 \$209053 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28415 VDD|pad|pin1|supply|vdd \$207279 \$209053 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28416 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$207279
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28417 VDD|pad|pin1|supply|vdd \$207254 \$207279 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28418 VDD|pad|pin1|supply|vdd \$207279 a2|q$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28419 \$167243 z$26 \$169909 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28420 \$169909 zn$3 \$169909 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28422 VDD|pad|pin1|supply|vdd a2|i|q$1 \$207280 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28423 \$207280 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28424 \$167243 zn$3 \$167243 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28425 d|z$6 \$207280 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28426 \$169910 z$26 \$167243 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28429 \$207282 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28430 VDD|pad|pin1|supply|vdd \$207282 \$207255 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28431 \$169910 zn$3 \$169910 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28432 VDD|pad|pin1|supply|vdd \$207255 \$209065 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28433 \$209065 d|z$15 \$207283 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28434 \$207283 \$207282 \$208956 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28435 \$208956 \$207284 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28436 \$169911 z$26 \$167243 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28438 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$208956
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28439 \$207284 \$207283 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28440 \$207284 \$207282 \$207256 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28441 \$207256 \$207255 \$209068 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28442 VDD|pad|pin1|supply|vdd \$207286 \$209068 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28443 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$207286
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28444 VDD|pad|pin1|supply|vdd \$207256 \$207286 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28445 VDD|pad|pin1|supply|vdd \$207286 a2|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28447 \$169911 zn$3 \$169911 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28448 a3|zn a1|a2|q$1 \$209074 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$28449 \$209074 a2|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$28450 VDD|pad|pin1|supply|vdd a2|q$2 \$207287 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28451 \$207287 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28452 d|z$7 \$207287 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28453 \$167244 z$26 \$169912 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28454 \$169912 zn$3 \$169912 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28455 VDD|pad|pin1|supply|vdd a2|q$1 \$207289 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28456 \$207289 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28458 d|z$8 \$207289 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28459 \$167244 zn$3 \$167244 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28460 \$207291 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28461 VDD|pad|pin1|supply|vdd \$207291 \$207257 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28462 VDD|pad|pin1|supply|vdd \$207257 \$209075 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28463 \$209075 d|z$16 \$207292 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28464 \$207292 \$207291 \$208958 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28465 \$208958 \$207293 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28466 \$169913 z$26 \$167244 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28469 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$208958
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28470 \$207293 \$207292 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28471 \$207293 \$207291 \$207258 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28472 \$207258 \$207257 \$209076 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28473 VDD|pad|pin1|supply|vdd \$207295 \$209076 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28474 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$207295
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28475 VDD|pad|pin1|supply|vdd \$207258 \$207295 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28476 VDD|pad|pin1|supply|vdd \$207295 a1|a2|q$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28477 \$169913 zn$3 \$169913 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28478 \$169914 z$26 \$167244 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28480 VDD|pad|pin1|supply|vdd a1|a2|q$2 \$207296 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28481 \$207296 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28483 d|z$9 \$207296 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28484 \$169914 zn$3 \$169914 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28485 \$207299 \$207260 \$207298 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28486 \$207299 R[32]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28487 VDD|pad|pin1|supply|vdd i0|i1|q \$207300 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28488 \$207300 s|zn \$207298 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28489 VDD|pad|pin1|supply|vdd s|zn \$207260 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28490 VDD|pad|pin1|supply|vdd \$207298 d|z$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28491 \$207303 \$207262 \$207302 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28492 \$207303 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28493 VDD|pad|pin1|supply|vdd R[28]|i0|q \$207305 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28494 \$207305 s|z \$207302 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28495 \$167245 z$26 \$169915 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28496 \$169915 zn$3 \$169915 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28497 VDD|pad|pin1|supply|vdd s|z \$207262 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28498 VDD|pad|pin1|supply|vdd \$207302 d|z$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28500 \$207307 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28501 VDD|pad|pin1|supply|vdd \$207307 \$207263 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28502 \$167245 zn$3 \$167245 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28503 VDD|pad|pin1|supply|vdd \$207263 \$209085 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28504 \$209085 d|z$11 \$207308 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28505 \$207308 \$207307 \$208959 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28506 \$208959 \$207309 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28507 \$169916 z$26 \$167245 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28509 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$208959
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28510 \$207309 \$207308 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28511 \$207309 \$207307 \$207264 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28512 \$207264 \$207263 \$209084 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28513 VDD|pad|pin1|supply|vdd \$207311 \$209084 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28514 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$207311
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28515 VDD|pad|pin1|supply|vdd \$207264 \$207311 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28516 VDD|pad|pin1|supply|vdd \$207311 R[28]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28518 \$169916 zn$3 \$169916 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28519 \$169917 z$26 \$167245 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28522 \$207313 \$207265 \$207312 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28523 \$207313 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28524 VDD|pad|pin1|supply|vdd R[25]|i0|q \$207314 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28525 \$207314 s|z \$207312 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28526 \$169917 zn$3 \$169917 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28527 VDD|pad|pin1|supply|vdd s|z \$207265 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28528 VDD|pad|pin1|supply|vdd \$207312 d|z$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28529 \$167246 z$26 \$169918 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28530 \$207316 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28531 VDD|pad|pin1|supply|vdd \$207316 \$207266 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28532 \$169918 zn$3 \$169918 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28533 VDD|pad|pin1|supply|vdd \$207266 \$209096 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28534 \$209096 d|z$17 \$207317 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28535 \$207317 \$207316 \$208960 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28536 \$208960 \$207318 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28538 \$167246 zn$3 \$167246 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28539 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$208960
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28540 \$207318 \$207317 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28541 \$207318 \$207316 \$207267 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28542 \$207267 \$207266 \$209108 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28543 VDD|pad|pin1|supply|vdd \$207320 \$209108 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28544 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$207320
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28545 VDD|pad|pin1|supply|vdd \$207267 \$207320 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28546 VDD|pad|pin1|supply|vdd \$207320 R[27]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28547 \$169919 z$26 \$167246 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28550 \$169919 zn$3 \$169919 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28551 \$207321 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28552 VDD|pad|pin1|supply|vdd \$207321 \$207268 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28553 VDD|pad|pin1|supply|vdd \$207268 \$209121 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28554 \$209121 d|z$18 \$207322 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28555 \$207322 \$207321 \$208963 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28556 \$208963 \$207323 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28557 \$169920 z$26 \$167246 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28560 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$208963
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28561 \$207323 \$207322 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28562 \$207323 \$207321 \$207269 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28563 \$207269 \$207268 \$209137 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28564 VDD|pad|pin1|supply|vdd \$207325 \$209137 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28565 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$207325
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28566 VDD|pad|pin1|supply|vdd \$207269 \$207325 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28567 VDD|pad|pin1|supply|vdd \$207325 R[33]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28568 \$169920 zn$3 \$169920 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28569 \$167247 z$26 \$169921 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28570 \$169921 zn$3 \$169921 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28571 \$207326 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28572 VDD|pad|pin1|supply|vdd \$207326 \$207270 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28574 VDD|pad|pin1|supply|vdd \$207270 \$209142 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28575 \$209142 d|z$19 \$207327 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28576 \$207327 \$207326 \$208964 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28577 \$208964 \$207328 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28578 \$167247 zn$3 \$167247 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28579 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$208964
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28580 \$207328 \$207327 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28581 \$207328 \$207326 \$207271 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28582 \$207271 \$207270 \$209147 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28583 VDD|pad|pin1|supply|vdd \$207330 \$209147 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28584 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$207330
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28585 VDD|pad|pin1|supply|vdd \$207271 \$207330 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28586 VDD|pad|pin1|supply|vdd \$207330 i0|i1|q$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28587 \$169922 z$26 \$167247 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28590 \$169922 zn$3 \$169922 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28591 \$169923 z$26 \$167247 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28592 \$207332 \$207272 \$207331 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28593 \$207332 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28594 VDD|pad|pin1|supply|vdd i0|i1|q$5 \$207333 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28595 \$207333 s|zn$1 \$207331 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28598 VDD|pad|pin1|supply|vdd s|zn$1 \$207272 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28599 VDD|pad|pin1|supply|vdd \$207331 d|z$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28600 \$169923 zn$3 \$169923 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28601 \$167248 z$26 \$169924 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28602 \$169924 zn$3 \$169924 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28604 \$167248 zn$3 \$167248 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28605 \$169925 z$26 \$167248 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28608 \$169925 zn$3 \$169925 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28609 \$169926 z$26 \$167248 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28612 \$169926 zn$3 \$169926 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28613 \$167249 z$26 \$169927 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28614 \$169927 zn$3 \$169927 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28616 \$167249 zn$3 \$167249 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28617 \$169928 z$26 \$167249 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28620 \$169928 zn$3 \$169928 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28621 \$169929 z$26 \$167249 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28624 \$169929 zn$3 \$169929 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28625 VDD|pad|pin1|supply|vdd VALID|a3|c2p|core|i|z \$181364
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$28626 VDD|pad|pin1|supply|vdd \$181364 RD[8]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$28627 \$167250 z$26 \$169930 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28628 \$169930 zn$3 \$169930 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28630 \$167250 zn$3 \$167250 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28631 \$169931 z$26 \$167250 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28634 \$169931 zn$3 \$169931 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28635 \$169932 z$26 \$167250 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28638 \$169932 zn$3 \$169932 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28639 VDD|pad|pin1|supply|vdd SAMPLE|a1|c2p|core|i|z \$181365
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$28640 VDD|pad|pin1|supply|vdd \$181365 RD[9]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$28641 \$167251 z$26 \$169933 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28642 \$169933 zn$3 \$169933 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28644 \$167251 zn$3 \$167251 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$28645 \$169934 z$26 \$167251 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28648 \$169934 zn$3 \$169934 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28649 \$169935 z$26 \$167251 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$28652 \$169935 zn$3 \$169935 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$28653 a1|z$9 a1|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$28654 a1|z$10 a1|b|i|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$28655 VDD|pad|pin1|supply|vdd a2|a3|z \$169864 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$28656 \$169864 RST|a1|b|cdn|core|i|p2c a2|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$28657 a1|z$4 RESULT[3]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$28658 \$200224 DOUT_DAT|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$28659 \$198889 DOUT_DAT|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$28660 VDD|pad|pin1|supply|vdd cp|i|z$2 \$209535 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28661 VDD|pad|pin1|supply|vdd \$209535 \$209536 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28662 VDD|pad|pin1|supply|vdd \$209539 \$209538 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28663 \$209537 \$209535 \$209538 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28664 VDD|pad|pin1|supply|vdd \$209536 \$209931 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28665 \$209931 d|z$24 \$209537 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28666 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209538
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28667 \$209540 \$209536 \$209833 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28668 VDD|pad|pin1|supply|vdd \$210072 \$209833 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28669 VDD|pad|pin1|supply|vdd \$209537 \$209539 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28670 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210072
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28671 VDD|pad|pin1|supply|vdd \$209540 \$210072 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28672 \$209539 \$209535 \$209540 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28673 VDD|pad|pin1|supply|vdd \$210072 a1|a2|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28674 a2|zn$7 a1|a2|q$4 \$209932 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$28675 \$209932 a2|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$28676 VDD|pad|pin1|supply|vdd a2|q$3 \$209542 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28677 VDD|pad|pin1|supply|vdd a1|b|d|z \$209542 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28678 VDD|pad|pin1|supply|vdd \$209542 d|z$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28679 VDD|pad|pin1|supply|vdd cp|i|z$2 \$209544 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28680 VDD|pad|pin1|supply|vdd \$209544 \$209545 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28681 VDD|pad|pin1|supply|vdd \$209548 \$209547 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28682 \$209546 \$209544 \$209547 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28683 VDD|pad|pin1|supply|vdd \$209545 \$209933 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28684 \$209933 d|z$20 \$209546 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28685 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209547
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28686 \$209549 \$209545 \$209844 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28687 VDD|pad|pin1|supply|vdd \$210075 \$209844 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28688 VDD|pad|pin1|supply|vdd \$209546 \$209548 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28689 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210075
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28690 VDD|pad|pin1|supply|vdd \$209549 \$210075 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28691 \$209548 \$209544 \$209549 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28692 VDD|pad|pin1|supply|vdd \$210075 a2|i|q$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28693 VDD|pad|pin1|supply|vdd a1|a2|q$5 \$209550 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28694 VDD|pad|pin1|supply|vdd a1|b|d|z \$209550 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28695 VDD|pad|pin1|supply|vdd \$209550 d|z$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28696 VDD|pad|pin1|supply|vdd a2|q \$209552 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28697 VDD|pad|pin1|supply|vdd a1|b|d|z \$209552 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28698 VDD|pad|pin1|supply|vdd \$209552 d|z$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28699 VDD|pad|pin1|supply|vdd cp|i|z$3 \$209554 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28700 VDD|pad|pin1|supply|vdd \$209554 \$209555 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28701 VDD|pad|pin1|supply|vdd \$209558 \$209557 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28702 \$209556 \$209554 \$209557 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28703 VDD|pad|pin1|supply|vdd \$209555 \$209938 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28704 \$209938 d|z$22 \$209556 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28705 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209557
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28706 \$209559 \$209555 \$209855 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28707 VDD|pad|pin1|supply|vdd \$210077 \$209855 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28708 VDD|pad|pin1|supply|vdd \$209556 \$209558 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28709 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210077
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28710 VDD|pad|pin1|supply|vdd \$209559 \$210077 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28711 \$209558 \$209554 \$209559 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28712 VDD|pad|pin1|supply|vdd \$210077 a2|q$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28713 VDD|pad|pin1|supply|vdd cp|i|z$3 \$209561 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28714 VDD|pad|pin1|supply|vdd \$209561 \$209562 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28715 VDD|pad|pin1|supply|vdd \$209565 \$209564 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28716 \$209563 \$209561 \$209564 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28717 VDD|pad|pin1|supply|vdd \$209562 \$209940 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28718 \$209940 d|z$7 \$209563 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28719 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209564
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28720 \$209566 \$209562 \$209863 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28721 VDD|pad|pin1|supply|vdd \$210078 \$209863 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28722 VDD|pad|pin1|supply|vdd \$209563 \$209565 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28723 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210078
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28724 VDD|pad|pin1|supply|vdd \$209566 \$210078 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28725 \$209565 \$209561 \$209566 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28726 VDD|pad|pin1|supply|vdd \$210078 a1|a2|q$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28727 VDD|pad|pin1|supply|vdd cp|i|z$3 \$209568 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28728 VDD|pad|pin1|supply|vdd \$209568 \$209569 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28729 VDD|pad|pin1|supply|vdd \$209572 \$209571 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28730 \$209570 \$209568 \$209571 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28731 VDD|pad|pin1|supply|vdd \$209569 \$209942 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28732 \$209942 d|z$9 \$209570 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28733 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209571
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28734 \$209573 \$209569 \$209865 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28735 VDD|pad|pin1|supply|vdd \$210079 \$209865 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28736 VDD|pad|pin1|supply|vdd \$209570 \$209572 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28737 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210079
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28738 VDD|pad|pin1|supply|vdd \$209573 \$210079 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28739 \$209572 \$209568 \$209573 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28740 VDD|pad|pin1|supply|vdd \$210079 a2|q$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28741 VDD|pad|pin1|supply|vdd cp|i|z$3 \$209574 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28742 VDD|pad|pin1|supply|vdd \$209574 \$209575 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28743 VDD|pad|pin1|supply|vdd \$209578 \$209577 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28744 \$209576 \$209574 \$209577 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28745 VDD|pad|pin1|supply|vdd \$209575 \$209941 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28746 \$209941 d|z$10 \$209576 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28747 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209577
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28748 \$209579 \$209575 \$209869 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28749 VDD|pad|pin1|supply|vdd \$210080 \$209869 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28750 VDD|pad|pin1|supply|vdd \$209576 \$209578 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28751 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210080
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28752 VDD|pad|pin1|supply|vdd \$209579 \$210080 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28753 \$209578 \$209574 \$209579 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28754 VDD|pad|pin1|supply|vdd \$210080 R[32]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28755 \$209580 \$209149 \$209581 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28756 \$209582 s|z \$209580 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28757 VDD|pad|pin1|supply|vdd R[26]|i0|q \$209582 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28758 \$209581 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28759 \$209149 s|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28760 VDD|pad|pin1|supply|vdd \$209580 d|z$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28761 VDD|pad|pin1|supply|vdd cp|i|z$4 \$209584 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28762 VDD|pad|pin1|supply|vdd \$209584 \$209585 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28763 VDD|pad|pin1|supply|vdd \$209588 \$209587 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28764 \$209586 \$209584 \$209587 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28765 VDD|pad|pin1|supply|vdd \$209585 \$209939 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28766 \$209939 d|z$23 \$209586 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28767 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209587
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28768 \$209589 \$209585 \$209873 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28769 VDD|pad|pin1|supply|vdd \$210083 \$209873 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28770 VDD|pad|pin1|supply|vdd \$209586 \$209588 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28771 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210083
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28772 VDD|pad|pin1|supply|vdd \$209589 \$210083 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28773 \$209588 \$209584 \$209589 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28774 VDD|pad|pin1|supply|vdd \$210083 R[26]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28775 VDD|pad|pin1|supply|vdd cp|i|z$4 \$209590 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28776 VDD|pad|pin1|supply|vdd \$209590 \$209591 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28777 VDD|pad|pin1|supply|vdd \$209594 \$209593 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28778 \$209592 \$209590 \$209593 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28779 VDD|pad|pin1|supply|vdd \$209591 \$209937 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28780 \$209937 d|z$12 \$209592 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28781 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209593
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28782 \$209595 \$209591 \$209874 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28783 VDD|pad|pin1|supply|vdd \$210084 \$209874 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28784 VDD|pad|pin1|supply|vdd \$209592 \$209594 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28785 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210084
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28786 VDD|pad|pin1|supply|vdd \$209595 \$210084 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28787 \$209594 \$209590 \$209595 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28788 VDD|pad|pin1|supply|vdd \$210084 R[25]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28789 VDD|pad|pin1|supply|vdd cp|i|z$1 \$209596 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28790 VDD|pad|pin1|supply|vdd \$209596 \$209597 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28791 VDD|pad|pin1|supply|vdd \$209600 \$209599 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28792 \$209598 \$209596 \$209599 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28793 VDD|pad|pin1|supply|vdd \$209597 \$209936 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28794 \$209936 d|z$25 \$209598 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28795 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209599
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28796 \$209601 \$209597 \$209892 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28797 VDD|pad|pin1|supply|vdd \$210086 \$209892 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28798 VDD|pad|pin1|supply|vdd \$209598 \$209600 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28799 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210086
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28800 VDD|pad|pin1|supply|vdd \$209601 \$210086 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28801 \$209600 \$209596 \$209601 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28802 VDD|pad|pin1|supply|vdd \$210086 R[24]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28803 VDD|pad|pin1|supply|vdd cp|i|z$1 \$209603 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28804 VDD|pad|pin1|supply|vdd \$209603 \$209604 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28805 VDD|pad|pin1|supply|vdd \$209607 \$209606 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28806 \$209605 \$209603 \$209606 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28807 VDD|pad|pin1|supply|vdd \$209604 \$209935 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28808 \$209935 d|z$26 \$209605 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28809 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209606
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28810 \$209608 \$209604 \$209926 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28811 VDD|pad|pin1|supply|vdd \$210088 \$209926 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28812 VDD|pad|pin1|supply|vdd \$209605 \$209607 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28813 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210088
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28814 VDD|pad|pin1|supply|vdd \$209608 \$210088 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28815 \$209607 \$209603 \$209608 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28816 VDD|pad|pin1|supply|vdd \$210088 R[34]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28817 VDD|pad|pin1|supply|vdd cp|i|z$1 \$209610 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28818 VDD|pad|pin1|supply|vdd \$209610 \$209611 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28819 VDD|pad|pin1|supply|vdd \$209614 \$209613 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28820 \$209612 \$209610 \$209613 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28821 VDD|pad|pin1|supply|vdd \$209611 \$209934 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28822 \$209934 d|z$27 \$209612 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28823 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209613
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28824 \$209615 \$209611 \$209927 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28825 VDD|pad|pin1|supply|vdd \$210090 \$209927 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28826 VDD|pad|pin1|supply|vdd \$209612 \$209614 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28827 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210090
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28828 VDD|pad|pin1|supply|vdd \$209615 \$210090 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28829 \$209614 \$209610 \$209615 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28830 VDD|pad|pin1|supply|vdd \$210090 i0|i1|q$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28831 VDD|pad|pin1|supply|vdd cp|i|z$1 \$209616 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28832 VDD|pad|pin1|supply|vdd \$209616 \$209617 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28833 VDD|pad|pin1|supply|vdd \$209620 \$209619 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28834 \$209618 \$209616 \$209619 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28835 VDD|pad|pin1|supply|vdd \$209617 \$209930 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28836 \$209930 d|z$28 \$209618 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28837 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209619
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28838 \$209621 \$209617 \$209920 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28839 VDD|pad|pin1|supply|vdd \$210092 \$209920 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28840 VDD|pad|pin1|supply|vdd \$209618 \$209620 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28841 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210092
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28842 VDD|pad|pin1|supply|vdd \$209621 \$210092 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28843 \$209620 \$209616 \$209621 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28844 VDD|pad|pin1|supply|vdd \$210092 i0|i1|q$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28845 VDD|pad|pin1|supply|vdd cp|i|z$1 \$209622 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28846 VDD|pad|pin1|supply|vdd \$209622 \$209623 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28847 VDD|pad|pin1|supply|vdd \$209626 \$209625 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28848 \$209624 \$209622 \$209625 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28849 VDD|pad|pin1|supply|vdd \$209623 \$209929 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28850 \$209929 d|z$13 \$209624 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28851 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$209625
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28852 \$209627 \$209623 \$209919 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28853 VDD|pad|pin1|supply|vdd \$210093 \$209919 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28854 VDD|pad|pin1|supply|vdd \$209624 \$209626 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28855 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$210093
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28856 VDD|pad|pin1|supply|vdd \$209627 \$210093 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28857 \$209626 \$209622 \$209627 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28858 VDD|pad|pin1|supply|vdd \$210093 i0|i1|q$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28859 \$211694 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28860 VDD|pad|pin1|supply|vdd \$211694 \$211695 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28861 VDD|pad|pin1|supply|vdd \$211695 \$213572 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28862 \$213572 d|z$5 \$211696 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28863 \$211696 \$211694 \$213209 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28864 \$213209 \$211697 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28865 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213209
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28866 \$211697 \$211696 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28867 \$211697 \$211694 \$211698 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28868 \$211698 \$211695 \$213582 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28869 VDD|pad|pin1|supply|vdd \$211700 \$213582 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28870 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211700
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28871 VDD|pad|pin1|supply|vdd \$211698 \$211700 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28872 VDD|pad|pin1|supply|vdd \$211700 a2|q$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28873 \$211701 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28874 VDD|pad|pin1|supply|vdd \$211701 \$211702 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28875 VDD|pad|pin1|supply|vdd \$211702 \$213579 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28876 \$213579 d|z$29 \$211703 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28877 \$211703 \$211701 \$213211 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28878 \$213211 \$211704 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28879 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213211
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28880 \$211704 \$211703 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28881 \$211704 \$211701 \$211705 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28882 \$211705 \$211702 \$213584 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28883 VDD|pad|pin1|supply|vdd \$211707 \$213584 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28884 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211707
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28885 VDD|pad|pin1|supply|vdd \$211705 \$211707 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28886 VDD|pad|pin1|supply|vdd \$211707 a1|a2|q$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28887 cp|i|z$2 \$211708 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$28888 VDD|pad|pin1|supply|vdd i|z$115 \$211708 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$28889 \$211709 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28890 VDD|pad|pin1|supply|vdd \$211709 \$211710 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28891 VDD|pad|pin1|supply|vdd \$211710 \$213581 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28892 \$213581 d|z$6 \$211711 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28893 \$211711 \$211709 \$213212 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28894 \$213212 \$211712 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28895 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213212
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28896 \$211712 \$211711 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28897 \$211712 \$211709 \$211713 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28898 \$211713 \$211710 \$213567 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28899 VDD|pad|pin1|supply|vdd \$211715 \$213567 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28900 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211715
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28901 VDD|pad|pin1|supply|vdd \$211713 \$211715 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28902 VDD|pad|pin1|supply|vdd \$211715 a1|a2|q$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28903 \$211716 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28904 VDD|pad|pin1|supply|vdd \$211716 \$211717 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28905 VDD|pad|pin1|supply|vdd \$211717 \$213574 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28906 \$213574 d|z$21 \$211718 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28907 \$211718 \$211716 \$213213 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28908 \$213213 \$211719 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28909 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213213
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28910 \$211719 \$211718 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28911 \$211719 \$211716 \$211720 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28912 \$211720 \$211717 \$213562 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28913 VDD|pad|pin1|supply|vdd \$211722 \$213562 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28914 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211722
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28915 VDD|pad|pin1|supply|vdd \$211720 \$211722 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28916 VDD|pad|pin1|supply|vdd \$211722 a1|a2|q$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28917 a4|zn a1|a2|q$5 \$213566 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$28918 \$213566 a2|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$28919 VDD|pad|pin1|supply|vdd a3|zn a2|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28920 a2|zn$9 a2|zn$8 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$28921 VDD|pad|pin1|supply|vdd a1|zn a2|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28922 a2|zn$9 a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28923 VDD|pad|pin1|supply|vdd a1|a2|q$3 \$211725 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28924 \$211725 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28925 d|z$16 \$211725 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28926 \$211726 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28927 VDD|pad|pin1|supply|vdd \$211726 \$211727 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28928 VDD|pad|pin1|supply|vdd \$211727 \$213560 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28929 \$213560 d|z$8 \$211728 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28930 \$211728 \$211726 \$213214 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28931 \$213214 \$211729 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28932 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213214
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28933 \$211729 \$211728 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28934 \$211729 \$211726 \$211730 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28935 \$211730 \$211727 \$213556 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28936 VDD|pad|pin1|supply|vdd \$211732 \$213556 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28937 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211732
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28938 VDD|pad|pin1|supply|vdd \$211730 \$211732 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28939 VDD|pad|pin1|supply|vdd \$211732 a2|q$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28940 \$211733 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28941 VDD|pad|pin1|supply|vdd \$211733 \$211734 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28942 VDD|pad|pin1|supply|vdd \$211734 \$213557 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28943 \$213557 d|z$30 \$211735 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28944 \$211735 \$211733 \$213216 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28945 \$213216 \$211736 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28946 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213216
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28947 \$211736 \$211735 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28948 \$211736 \$211733 \$211737 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28949 \$211737 \$211734 \$213554 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28950 VDD|pad|pin1|supply|vdd \$211739 \$213554 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28951 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211739
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28952 VDD|pad|pin1|supply|vdd \$211737 \$211739 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28953 VDD|pad|pin1|supply|vdd \$211739 i0|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28954 \$211740 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28955 VDD|pad|pin1|supply|vdd \$211740 \$211741 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28956 VDD|pad|pin1|supply|vdd \$211741 \$213549 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28957 \$213549 d|z$31 \$211742 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28958 \$211742 \$211740 \$213217 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28959 \$213217 \$211743 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28960 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213217
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28961 \$211743 \$211742 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28962 \$211743 \$211740 \$211744 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28963 \$211744 \$211741 \$213550 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28964 VDD|pad|pin1|supply|vdd \$211746 \$213550 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28965 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211746
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28966 VDD|pad|pin1|supply|vdd \$211744 \$211746 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28967 VDD|pad|pin1|supply|vdd \$211746 R[29]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28968 \$211747 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28969 VDD|pad|pin1|supply|vdd \$211747 \$211748 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28970 VDD|pad|pin1|supply|vdd \$211748 \$213548 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28971 \$213548 d|z$32 \$211749 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28972 \$211749 \$211747 \$213219 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28973 \$213219 \$211750 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28974 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213219
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28975 \$211750 \$211749 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28976 \$211750 \$211747 \$211751 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28977 \$211751 \$211748 \$213540 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28978 VDD|pad|pin1|supply|vdd \$211753 \$213540 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28979 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211753
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28980 VDD|pad|pin1|supply|vdd \$211751 \$211753 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28981 VDD|pad|pin1|supply|vdd \$211753 R[36]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28982 \$211755 \$211757 \$211754 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28983 \$211755 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28984 VDD|pad|pin1|supply|vdd R[24]|i0|q \$211756 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28985 \$211756 s|z \$211754 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28986 VDD|pad|pin1|supply|vdd s|z \$211757 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28987 VDD|pad|pin1|supply|vdd \$211754 d|z$25 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28988 \$211758 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28989 VDD|pad|pin1|supply|vdd \$211758 \$211759 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28990 VDD|pad|pin1|supply|vdd \$211759 \$213539 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28991 \$213539 d|z$33 \$211760 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28992 \$211760 \$211758 \$213221 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28993 \$213221 \$211761 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28994 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213221
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28995 \$211761 \$211760 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28996 \$211761 \$211758 \$211762 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28997 \$211762 \$211759 \$213538 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28998 VDD|pad|pin1|supply|vdd \$211764 \$213538 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28999 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211764
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29000 VDD|pad|pin1|supply|vdd \$211762 \$211764 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29001 VDD|pad|pin1|supply|vdd \$211764 R[30]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29002 \$211766 \$211768 \$211765 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29003 \$211766 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29004 VDD|pad|pin1|supply|vdd R[27]|i0|q \$211767 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29005 \$211767 s|z \$211765 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29006 VDD|pad|pin1|supply|vdd s|z \$211768 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29007 VDD|pad|pin1|supply|vdd \$211765 d|z$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29008 \$211770 \$211772 \$211769 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29009 \$211770 R[34]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29010 VDD|pad|pin1|supply|vdd i0|i1|q$2 \$211771 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29011 \$211771 s|zn \$211769 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29012 VDD|pad|pin1|supply|vdd s|zn \$211772 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29013 VDD|pad|pin1|supply|vdd \$211769 d|z$26 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29014 \$211775 \$211777 \$211773 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29015 \$211775 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29016 VDD|pad|pin1|supply|vdd i0|i1|q$6 \$211776 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29017 \$211776 s|zn$1 \$211773 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29018 VDD|pad|pin1|supply|vdd s|zn$1 \$211777 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29019 VDD|pad|pin1|supply|vdd \$211773 d|z$27 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29020 \$211779 \$211781 \$211778 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29021 \$211779 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29022 VDD|pad|pin1|supply|vdd i0|i1|q$2 \$211780 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29023 \$211780 s|zn$1 \$211778 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29024 VDD|pad|pin1|supply|vdd s|zn$1 \$211781 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29025 VDD|pad|pin1|supply|vdd \$211778 d|z$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29026 cp|i|z$1 \$211782 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$29027 VDD|pad|pin1|supply|vdd i|z$115 \$211782 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$29028 z$28 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29029 \$211784 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29030 VDD|pad|pin1|supply|vdd \$211784 \$211785 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29031 VDD|pad|pin1|supply|vdd \$211785 \$213535 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29032 \$213535 d|z$34 \$211786 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29033 \$211786 \$211784 \$213223 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29034 \$213223 \$211787 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29035 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213223
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29036 \$211787 \$211786 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29037 \$211787 \$211784 \$211788 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29038 \$211788 \$211785 \$213531 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29039 VDD|pad|pin1|supply|vdd \$211790 \$213531 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29040 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211790
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29041 VDD|pad|pin1|supply|vdd \$211788 \$211790 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29042 VDD|pad|pin1|supply|vdd \$211790 i0|i1|q$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29043 \$211791 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29044 VDD|pad|pin1|supply|vdd \$211791 \$211792 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29045 VDD|pad|pin1|supply|vdd \$211792 \$213526 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29046 \$213526 d|z$35 \$211793 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29047 \$211793 \$211791 \$213224 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29048 \$213224 \$211794 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29049 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213224
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29050 \$211794 \$211793 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29051 \$211794 \$211791 \$211795 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29052 \$211795 \$211792 \$213528 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29053 VDD|pad|pin1|supply|vdd \$211797 \$213528 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29054 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$211797
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29055 VDD|pad|pin1|supply|vdd \$211795 \$211797 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29056 VDD|pad|pin1|supply|vdd \$211797 i0|i1|q$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29057 VDD|pad|pin1|supply|vdd a2|q$6 \$213634 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29058 VDD|pad|pin1|supply|vdd a1|b|d|z \$213634 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29059 VDD|pad|pin1|supply|vdd \$213634 d|z$24 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29060 VDD|pad|pin1|supply|vdd cp|i|z$2 \$213635 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29061 VDD|pad|pin1|supply|vdd \$213635 \$213636 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29062 VDD|pad|pin1|supply|vdd \$213639 \$213638 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29063 \$213637 \$213635 \$213638 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29064 VDD|pad|pin1|supply|vdd \$213636 \$214320 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29065 \$214320 d|z$38 \$213637 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29066 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213638
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29067 \$213640 \$213636 \$213842 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29068 VDD|pad|pin1|supply|vdd \$214361 \$213842 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29069 VDD|pad|pin1|supply|vdd \$213637 \$213639 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29070 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$214361
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29071 VDD|pad|pin1|supply|vdd \$213640 \$214361 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29072 \$213639 \$213635 \$213640 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29073 VDD|pad|pin1|supply|vdd \$214361 a2|q$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29074 VDD|pad|pin1|supply|vdd a2|q$4 \$215804 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29075 \$215804 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29076 VDD|pad|pin1|supply|vdd a1|a2|q$6 \$213642 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29077 VDD|pad|pin1|supply|vdd a1|b|d|z \$213642 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29078 d|z$29 \$215804 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29079 VDD|pad|pin1|supply|vdd \$213642 d|z$38 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29080 a3|zn$1 a1|a2|q$6 \$217241 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29081 \$217241 a2|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29082 VDD|pad|pin1|supply|vdd a1|a2|q$4 \$213643 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29083 VDD|pad|pin1|supply|vdd a1|b|d|z \$213643 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29084 a4|zn$1 a1|a2|q \$217253 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29085 \$217253 a2|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29086 VDD|pad|pin1|supply|vdd \$213643 d|z$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29087 VDD|pad|pin1|supply|vdd a3|zn$1 a2|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29088 VDD|pad|pin1|supply|vdd a2|zn$7 a2|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$29089 VDD|pad|pin1|supply|vdd a1|z$14 a2|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$29090 z$31 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29091 VDD|pad|pin1|supply|vdd a4|zn$1 a2|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29092 a1|z$14 a2|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29093 VDD|pad|pin1|supply|vdd a1|b|d|z s|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29094 s|zn$1 a1|zn$1 \$214326 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.4565p AD=0.4565p PS=1.93u PD=1.93u
M$29095 \$214326 a2|zn$10 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29096 VDD|pad|pin1|supply|vdd cp|i|z$2 \$213645 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29097 VDD|pad|pin1|supply|vdd \$213645 \$213646 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29098 VDD|pad|pin1|supply|vdd \$213649 \$213648 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29099 \$213647 \$213645 \$213648 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29100 VDD|pad|pin1|supply|vdd \$213646 \$214325 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29101 \$214325 d|z$41 \$213647 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29102 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213648
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29103 \$213650 \$213646 \$213855 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29104 VDD|pad|pin1|supply|vdd \$214362 \$213855 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29105 VDD|pad|pin1|supply|vdd \$213647 \$213649 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29106 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$214362
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29107 VDD|pad|pin1|supply|vdd \$213650 \$214362 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29108 \$213649 \$213645 \$213650 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29109 VDD|pad|pin1|supply|vdd \$214362 a1|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29110 VDD|pad|pin1|supply|vdd a2|i|q$2 \$215812 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29111 \$215812 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29112 d|s|z \$215812 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29113 \$215815 \$215509 \$215814 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29114 \$215815 DATA|core|i0|i1|p2c VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p
+ PS=1.93u PD=1.93u
M$29115 VDD|pad|pin1|supply|vdd a1|i0|q$1 \$215816 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29116 \$215816 d|s|zn \$215814 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29117 VDD|pad|pin1|supply|vdd a2|zn$9 a2|i|s|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29118 a2|i|s|zn a1|i0|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29119 VDD|pad|pin1|supply|vdd a1|a2|q$1 \$213652 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29120 VDD|pad|pin1|supply|vdd a1|b|d|z \$213652 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29121 VDD|pad|pin1|supply|vdd \$213652 d|z$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29122 VDD|pad|pin1|supply|vdd cp|i|z$3 \$213653 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29123 VDD|pad|pin1|supply|vdd \$213653 \$213654 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29124 \$215820 \$215510 \$215819 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29125 \$215820 a1|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29126 VDD|pad|pin1|supply|vdd i0|i1|q$4 \$215821 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29127 \$215821 s|zn$1 \$215819 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29128 VDD|pad|pin1|supply|vdd \$213657 \$213656 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29129 \$213655 \$213653 \$213656 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29130 VDD|pad|pin1|supply|vdd \$213654 \$214330 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29131 \$214330 d|z$42 \$213655 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29132 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213656
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29133 \$213658 \$213654 \$213863 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29134 VDD|pad|pin1|supply|vdd \$214363 \$213863 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29135 VDD|pad|pin1|supply|vdd \$213655 \$213657 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29136 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$214363
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29137 VDD|pad|pin1|supply|vdd \$213658 \$214363 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29138 \$213657 \$213653 \$213658 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29139 VDD|pad|pin1|supply|vdd \$214363 a1|i|i0|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29140 z$29 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29141 a2|zn$8 a1|a2|q$3 \$214331 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29142 \$214331 a2|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29143 VDD|pad|pin1|supply|vdd i|z$115 \$213661 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$29144 VDD|pad|pin1|supply|vdd \$213661 cp|i|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$29145 \$213662 \$213585 \$213663 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29146 \$213664 s|zn$1 \$213662 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29147 VDD|pad|pin1|supply|vdd DATA|core|i0|i1|p2c \$213664
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p
+ PS=1.93u PD=1.74u
M$29148 \$213663 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29149 a1|zn a1|a2|q$2 \$217293 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29150 \$217293 a2|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29151 \$213585 s|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29152 VDD|pad|pin1|supply|vdd \$213662 d|z$30 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29153 VDD|pad|pin1|supply|vdd cp|i|z$3 \$213665 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29154 VDD|pad|pin1|supply|vdd \$213665 \$213666 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29155 VDD|pad|pin1|supply|vdd \$213669 \$213668 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29156 \$213667 \$213665 \$213668 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29157 VDD|pad|pin1|supply|vdd \$213666 \$214333 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29158 \$214333 d|z$39 \$213667 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29159 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213668
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29160 \$213670 \$213666 \$213936 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29161 VDD|pad|pin1|supply|vdd \$214364 \$213936 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29162 VDD|pad|pin1|supply|vdd \$213667 \$213669 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29163 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$214364
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29164 VDD|pad|pin1|supply|vdd \$213670 \$214364 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29165 \$213669 \$213665 \$213670 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29166 VDD|pad|pin1|supply|vdd \$214364 R[21]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29167 \$213672 \$213586 \$213673 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29168 \$213674 s|z \$213672 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29169 VDD|pad|pin1|supply|vdd R[29]|i0|q \$213674 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29170 \$213673 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29171 \$213586 s|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29172 VDD|pad|pin1|supply|vdd \$213672 d|z$31 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29173 \$213675 \$213587 \$213676 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29174 \$213677 s|zn \$213675 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29175 VDD|pad|pin1|supply|vdd i0|i1|q$4 \$213677 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29176 \$213676 R[39]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29177 \$213587 s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29178 VDD|pad|pin1|supply|vdd \$213675 d|z$36 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29179 \$213679 \$213588 \$213680 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29180 \$213681 s|zn \$213679 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29181 VDD|pad|pin1|supply|vdd i0|i1|q$5 \$213681 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29182 \$213680 R[36]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29183 \$213588 s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29184 VDD|pad|pin1|supply|vdd \$213679 d|z$32 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29185 z$30 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29186 VDD|pad|pin1|supply|vdd i|z$115 \$213683 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$29187 VDD|pad|pin1|supply|vdd \$213683 cp|i|z$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$29188 \$213684 \$213589 \$213685 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29189 \$213686 s|z \$213684 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29190 VDD|pad|pin1|supply|vdd R[30]|i0|q \$213686 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29191 \$213685 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29192 \$215846 \$215519 \$215845 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29193 \$215846 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29194 VDD|pad|pin1|supply|vdd R[22]|i0|q \$215847 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29195 \$215847 s|zn$2 \$215845 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29196 \$213589 s|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29197 VDD|pad|pin1|supply|vdd \$213684 d|z$33 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29198 VDD|pad|pin1|supply|vdd cp|i|z$1 \$213687 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29199 VDD|pad|pin1|supply|vdd \$213687 \$213688 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29200 VDD|pad|pin1|supply|vdd \$213691 \$213690 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29201 \$213689 \$213687 \$213690 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29202 VDD|pad|pin1|supply|vdd \$213688 \$214359 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29203 \$214359 d|z$40 \$213689 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29204 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213690
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29205 \$213692 \$213688 \$214175 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29206 VDD|pad|pin1|supply|vdd \$214367 \$214175 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29207 VDD|pad|pin1|supply|vdd \$213689 \$213691 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29208 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$214367
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29209 VDD|pad|pin1|supply|vdd \$213692 \$214367 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29210 \$213691 \$213687 \$213692 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29211 VDD|pad|pin1|supply|vdd \$214367 R[20]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29212 \$213694 \$213590 \$213695 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29213 \$213696 s|zn \$213694 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29214 VDD|pad|pin1|supply|vdd i0|i1|q$6 \$213696 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29215 \$213695 R[33]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29216 \$213590 s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29217 VDD|pad|pin1|supply|vdd \$213694 d|z$18 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29218 \$213697 \$213591 \$213698 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29219 \$213699 s|zn \$213697 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29220 VDD|pad|pin1|supply|vdd i0|i1|q$7 \$213699 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29221 \$213698 R[37]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29222 \$215855 \$215522 \$215854 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29223 \$215855 R[35]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29224 VDD|pad|pin1|supply|vdd i0|i1|q$1 \$215856 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29225 \$215856 s|zn \$215854 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29226 \$213591 s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29227 VDD|pad|pin1|supply|vdd \$213697 d|z$37 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29228 VDD|pad|pin1|supply|vdd cp|z$4 \$213701 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29229 VDD|pad|pin1|supply|vdd \$213701 \$213702 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29230 VDD|pad|pin1|supply|vdd \$213705 \$213704 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29231 \$213703 \$213701 \$213704 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29232 VDD|pad|pin1|supply|vdd \$213702 \$214355 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29233 \$214355 d|z$37 \$213703 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29234 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213704
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29235 \$213706 \$213702 \$214182 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29236 VDD|pad|pin1|supply|vdd \$214369 \$214182 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29237 VDD|pad|pin1|supply|vdd \$213703 \$213705 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29238 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$214369
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29239 VDD|pad|pin1|supply|vdd \$213706 \$214369 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29240 \$213705 \$213701 \$213706 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29241 VDD|pad|pin1|supply|vdd \$214369 R[37]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29242 \$213708 \$213592 \$213709 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29243 \$213710 s|zn$1 \$213708 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29244 VDD|pad|pin1|supply|vdd i0|i1|q$1 \$213710 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29245 \$213709 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29246 \$213592 s|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29247 VDD|pad|pin1|supply|vdd \$213708 d|z$28 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29248 \$213711 \$213593 \$213712 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29249 \$213713 s|zn$1 \$213711 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29250 VDD|pad|pin1|supply|vdd i0|i1|q \$213713 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29251 \$213712 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29252 \$215863 \$215525 \$215862 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29253 \$215863 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29254 VDD|pad|pin1|supply|vdd i0|i1|q$7 \$215864 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29255 \$215864 s|zn$1 \$215862 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29256 \$213593 s|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29257 VDD|pad|pin1|supply|vdd \$213711 d|z$34 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29258 \$215866 \$215526 \$215865 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29259 \$215866 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29260 VDD|pad|pin1|supply|vdd i0|i1|q$3 \$215867 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29261 \$215867 s|zn$1 \$215865 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29262 VDD|pad|pin1|supply|vdd cp|z$4 \$213714 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29263 VDD|pad|pin1|supply|vdd \$213714 \$213715 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29264 VDD|pad|pin1|supply|vdd \$213718 \$213717 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29265 \$213716 \$213714 \$213717 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29266 VDD|pad|pin1|supply|vdd \$213715 \$214353 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29267 \$214353 d|z$43 \$213716 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29268 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$213717
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29269 \$213719 \$213715 \$214161 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29270 VDD|pad|pin1|supply|vdd \$214371 \$214161 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29271 VDD|pad|pin1|supply|vdd \$213716 \$213718 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29272 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$214371
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29273 VDD|pad|pin1|supply|vdd \$213719 \$214371 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29274 \$213718 \$213714 \$213719 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29275 VDD|pad|pin1|supply|vdd \$214371 i0|i1|q$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29276 VDD|pad|pin1|supply|vdd \$215504 \$217221 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29277 \$217221 d|z$50 \$215800 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29278 \$215800 \$215799 \$217080 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29279 \$217080 \$215801 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29280 VDD|pad|pin1|supply|vdd \$215506 \$217246 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29281 \$217246 a1|b|d|z \$215807 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29282 \$215807 \$215806 \$217081 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29283 \$217081 \$215808 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29284 VDD|pad|pin1|supply|vdd \$215511 \$217278 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29285 \$217278 d|z$46 \$215823 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29286 \$215823 \$215822 \$217082 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29287 \$217082 \$215824 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29288 VDD|pad|pin1|supply|vdd \$215513 \$217306 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29289 \$217306 d|z$47 \$215829 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29290 \$215829 \$215828 \$217083 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29291 \$217083 \$215830 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29292 VDD|pad|pin1|supply|vdd \$215515 \$217316 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29293 \$217316 d|z$36 \$215835 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29294 \$215835 \$215834 \$217084 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29295 \$217084 \$215836 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29296 VDD|pad|pin1|supply|vdd \$215517 \$217325 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29297 \$217325 d|z$48 \$215840 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29298 \$215840 \$215839 \$217085 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29299 \$217085 \$215841 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29300 VDD|pad|pin1|supply|vdd \$215520 \$217349 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29301 \$217349 d|z$45 \$215850 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29302 \$215850 \$215849 \$217086 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29303 \$217086 \$215851 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29304 VDD|pad|pin1|supply|vdd \$215523 \$217377 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29305 \$217377 d|z$49 \$215858 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29306 \$215858 \$215857 \$217087 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29307 \$217087 \$215859 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29308 VDD|pad|pin1|supply|vdd \$215527 \$217409 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29309 \$217409 d|z$51 \$215869 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29310 \$215869 \$215868 \$217088 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29311 \$217088 \$215870 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29312 \$215799 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29313 VDD|pad|pin1|supply|vdd \$215799 \$215504 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29314 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217080
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29315 \$215801 \$215800 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29316 \$215801 \$215799 \$215505 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29317 \$215505 \$215504 \$217235 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29318 VDD|pad|pin1|supply|vdd \$215803 \$217235 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29319 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$215803
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29320 VDD|pad|pin1|supply|vdd \$215505 \$215803 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29321 VDD|pad|pin1|supply|vdd \$215803 a1|a2|q$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29322 \$215806 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29323 VDD|pad|pin1|supply|vdd \$215806 \$215506 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29324 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217081
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29325 \$215808 \$215807 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29326 \$215808 \$215806 \$215507 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29327 \$215507 \$215506 \$217256 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29328 VDD|pad|pin1|supply|vdd \$215810 \$217256 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29329 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$215810
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29330 VDD|pad|pin1|supply|vdd \$215507 \$215810 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29331 VDD|pad|pin1|supply|vdd \$215810 a1|a2|q$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29332 VDD|pad|pin1|supply|vdd d|s|zn \$215509 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29333 VDD|pad|pin1|supply|vdd \$215814 d|z$44 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29334 VDD|pad|pin1|supply|vdd s|zn$1 \$215510 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29335 VDD|pad|pin1|supply|vdd \$215819 d|z$42 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29336 \$215822 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29337 VDD|pad|pin1|supply|vdd \$215822 \$215511 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29338 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217082
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29339 \$215824 \$215823 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29340 \$215824 \$215822 \$215512 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29341 \$215512 \$215511 \$217285 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29342 VDD|pad|pin1|supply|vdd \$215826 \$217285 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29343 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$215826
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29344 VDD|pad|pin1|supply|vdd \$215512 \$215826 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29345 VDD|pad|pin1|supply|vdd \$215826 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29346 \$215828 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29347 VDD|pad|pin1|supply|vdd \$215828 \$215513 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29348 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217083
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29349 \$215830 \$215829 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29350 \$215830 \$215828 \$215514 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29351 \$215514 \$215513 \$217315 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29352 VDD|pad|pin1|supply|vdd \$215832 \$217315 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29353 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$215832
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29354 VDD|pad|pin1|supply|vdd \$215514 \$215832 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29355 VDD|pad|pin1|supply|vdd \$215832 R[18]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29356 \$215834 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29357 VDD|pad|pin1|supply|vdd \$215834 \$215515 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29358 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217084
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29359 \$215836 \$215835 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29360 \$215836 \$215834 \$215516 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29361 \$215516 \$215515 \$217318 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29362 VDD|pad|pin1|supply|vdd \$215838 \$217318 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29363 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$215838
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29364 VDD|pad|pin1|supply|vdd \$215516 \$215838 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29365 VDD|pad|pin1|supply|vdd \$215838 R[39]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29366 \$215839 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29367 VDD|pad|pin1|supply|vdd \$215839 \$215517 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29368 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217085
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29369 \$215841 \$215840 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29370 \$215841 \$215839 \$215518 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29371 \$215518 \$215517 \$217319 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29372 VDD|pad|pin1|supply|vdd \$215843 \$217319 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29373 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$215843
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29374 VDD|pad|pin1|supply|vdd \$215518 \$215843 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29375 VDD|pad|pin1|supply|vdd \$215843 R[23]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29376 VDD|pad|pin1|supply|vdd s|zn$2 \$215519 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29377 VDD|pad|pin1|supply|vdd \$215845 d|z$45 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29378 \$215849 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29379 VDD|pad|pin1|supply|vdd \$215849 \$215520 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29380 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217086
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29381 \$215851 \$215850 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29382 \$215851 \$215849 \$215521 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29383 \$215521 \$215520 \$217342 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29384 VDD|pad|pin1|supply|vdd \$215853 \$217342 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29385 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$215853
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29386 VDD|pad|pin1|supply|vdd \$215521 \$215853 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29387 VDD|pad|pin1|supply|vdd \$215853 R[22]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29388 VDD|pad|pin1|supply|vdd s|zn \$215522 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29389 VDD|pad|pin1|supply|vdd \$215854 d|z$49 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29390 \$215857 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29391 VDD|pad|pin1|supply|vdd \$215857 \$215523 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29392 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217087
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29393 \$215859 \$215858 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29394 \$215859 \$215857 \$215524 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29395 \$215524 \$215523 \$217371 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29396 VDD|pad|pin1|supply|vdd \$215861 \$217371 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29397 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$215861
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29398 VDD|pad|pin1|supply|vdd \$215524 \$215861 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29399 VDD|pad|pin1|supply|vdd \$215861 R[35]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29400 VDD|pad|pin1|supply|vdd s|zn$1 \$215525 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29401 VDD|pad|pin1|supply|vdd \$215862 d|z$35 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29402 VDD|pad|pin1|supply|vdd s|zn$1 \$215526 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29403 VDD|pad|pin1|supply|vdd \$215865 d|z$43 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29404 \$215868 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29405 VDD|pad|pin1|supply|vdd \$215868 \$215527 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29406 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217088
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29407 \$215870 \$215869 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29408 \$215870 \$215868 \$215528 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29409 \$215528 \$215527 \$217424 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29410 VDD|pad|pin1|supply|vdd \$215872 \$217424 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29411 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$215872
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29412 VDD|pad|pin1|supply|vdd \$215528 \$215872 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29413 VDD|pad|pin1|supply|vdd \$215872 R[53]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29414 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$217719 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29415 VDD|pad|pin1|supply|vdd a1|b|d|z \$217719 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29416 VDD|pad|pin1|supply|vdd \$217719 d|z$50 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29417 VDD|pad|pin1|supply|vdd cp|i|z$5 \$217661 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29418 VDD|pad|pin1|supply|vdd \$217661 \$217720 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29419 VDD|pad|pin1|supply|vdd \$218407 \$217722 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29420 \$217721 \$217661 \$217722 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29421 VDD|pad|pin1|supply|vdd \$217720 \$218025 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29422 \$218025 d|s|z \$217721 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29423 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217722
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29424 \$217723 \$217720 \$218022 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29425 VDD|pad|pin1|supply|vdd \$218627 \$218022 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29426 VDD|pad|pin1|supply|vdd \$217721 \$218407 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29427 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$218627
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29428 VDD|pad|pin1|supply|vdd \$217723 \$218627 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29429 \$218407 \$217661 \$217723 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29430 VDD|pad|pin1|supply|vdd \$218627 a1|a2|q$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29431 VDD|pad|pin1|supply|vdd a2|q$7 \$217725 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29432 VDD|pad|pin1|supply|vdd a1|b|d|z \$217725 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29433 VDD|pad|pin1|supply|vdd \$217725 d|z$52 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29434 a2|z$8 a2|i|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29435 VDD|pad|pin1|supply|vdd a3|zn$2 a1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29436 VDD|pad|pin1|supply|vdd a2|z$8 a1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$29437 VDD|pad|pin1|supply|vdd a1|a2|q$7 a1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$29438 VDD|pad|pin1|supply|vdd a4|zn$2 a1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29439 VDD|pad|pin1|supply|vdd cp|i|z$6 \$217662 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29440 VDD|pad|pin1|supply|vdd \$217662 \$217729 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29441 VDD|pad|pin1|supply|vdd \$218408 \$217731 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29442 \$217730 \$217662 \$217731 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29443 VDD|pad|pin1|supply|vdd \$217729 \$218033 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29444 \$218033 d|s|zn \$217730 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29445 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217731
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29446 \$217732 \$217729 \$218035 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29447 VDD|pad|pin1|supply|vdd \$218628 \$218035 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29448 VDD|pad|pin1|supply|vdd \$217730 \$218408 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29449 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$218628
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29450 VDD|pad|pin1|supply|vdd \$217732 \$218628 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29451 \$218408 \$217662 \$217732 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29452 VDD|pad|pin1|supply|vdd \$218628 a2|i|q$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29453 VDD|pad|pin1|supply|vdd cp|i|z$6 \$217663 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29454 VDD|pad|pin1|supply|vdd \$217663 \$217733 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29455 VDD|pad|pin1|supply|vdd \$218409 \$217735 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29456 \$217734 \$217663 \$217735 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29457 VDD|pad|pin1|supply|vdd \$217733 \$218040 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29458 \$218040 d|z$44 \$217734 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29459 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217735
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29460 \$217736 \$217733 \$218046 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29461 VDD|pad|pin1|supply|vdd \$218629 \$218046 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29462 VDD|pad|pin1|supply|vdd \$217734 \$218409 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29463 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$218629
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29464 VDD|pad|pin1|supply|vdd \$217736 \$218629 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29465 \$218409 \$217663 \$217736 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29466 VDD|pad|pin1|supply|vdd \$218629 a1|i0|q$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29467 VDD|pad|pin1|supply|vdd cp|i|z$3 \$217664 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29468 VDD|pad|pin1|supply|vdd \$217664 \$217737 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29469 VDD|pad|pin1|supply|vdd \$218410 \$217739 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29470 \$217738 \$217664 \$217739 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29471 VDD|pad|pin1|supply|vdd \$217737 \$218050 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29472 \$218050 d|z$55 \$217738 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29473 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217739
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29474 \$217740 \$217737 \$218054 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29475 VDD|pad|pin1|supply|vdd \$218630 \$218054 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29476 VDD|pad|pin1|supply|vdd \$217738 \$218410 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29477 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$218630
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29478 VDD|pad|pin1|supply|vdd \$217740 \$218630 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29479 \$218410 \$217664 \$217740 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29480 VDD|pad|pin1|supply|vdd \$218630 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29481 VDD|pad|pin1|supply|vdd cp|i|z$3 \$217665 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29482 VDD|pad|pin1|supply|vdd \$217665 \$217742 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29483 VDD|pad|pin1|supply|vdd \$218411 \$217744 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29484 \$217743 \$217665 \$217744 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29485 VDD|pad|pin1|supply|vdd \$217742 \$218057 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29486 \$218057 d|z$56 \$217743 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29487 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217744
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29488 \$217746 \$217742 \$218062 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29489 VDD|pad|pin1|supply|vdd \$218631 \$218062 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29490 VDD|pad|pin1|supply|vdd \$217743 \$218411 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29491 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$218631
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29492 VDD|pad|pin1|supply|vdd \$217746 \$218631 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29493 \$218411 \$217665 \$217746 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29494 VDD|pad|pin1|supply|vdd \$218631 R[50]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29495 \$217747 \$217666 \$217748 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29496 \$217749 s|zn$2 \$217747 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29497 VDD|pad|pin1|supply|vdd R[18]|i0|q \$217749 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29498 \$217748 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29499 \$217666 s|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29500 VDD|pad|pin1|supply|vdd \$217747 d|z$47 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29501 \$217750 \$217668 \$217751 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29502 \$217752 s|zn$2 \$217750 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29503 VDD|pad|pin1|supply|vdd R[21]|i0|q \$217752 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29504 \$217751 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29505 \$217668 s|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29506 VDD|pad|pin1|supply|vdd \$217750 d|z$39 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29507 VDD|pad|pin1|supply|vdd cp|i|z$4 \$217669 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29508 VDD|pad|pin1|supply|vdd \$217669 \$217753 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29509 VDD|pad|pin1|supply|vdd \$218412 \$217755 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29510 \$217754 \$217669 \$217755 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29511 VDD|pad|pin1|supply|vdd \$217753 \$218067 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29512 \$218067 d|z$57 \$217754 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29513 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217755
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29514 \$217756 \$217753 \$218071 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29515 VDD|pad|pin1|supply|vdd \$218632 \$218071 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29516 VDD|pad|pin1|supply|vdd \$217754 \$218412 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29517 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$218632
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29518 VDD|pad|pin1|supply|vdd \$217756 \$218632 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29519 \$218412 \$217669 \$217756 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29520 VDD|pad|pin1|supply|vdd \$218632 R[31]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29521 VDD|pad|pin1|supply|vdd cp|i|z$4 \$217670 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29522 VDD|pad|pin1|supply|vdd \$217670 \$217758 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29523 VDD|pad|pin1|supply|vdd \$218413 \$217760 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29524 \$217759 \$217670 \$217760 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29525 VDD|pad|pin1|supply|vdd \$217758 \$218079 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29526 \$218079 d|z$58 \$217759 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29527 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217760
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29528 \$217761 \$217758 \$218107 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29529 VDD|pad|pin1|supply|vdd \$218633 \$218107 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29530 VDD|pad|pin1|supply|vdd \$217759 \$218413 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29531 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$218633
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29532 VDD|pad|pin1|supply|vdd \$217761 \$218633 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29533 \$218413 \$217670 \$217761 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29534 VDD|pad|pin1|supply|vdd \$218633 R[17]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29535 VDD|pad|pin1|supply|vdd cp|i|z$4 \$217671 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29536 VDD|pad|pin1|supply|vdd \$217671 \$217763 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29537 VDD|pad|pin1|supply|vdd \$218414 \$217765 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29538 \$217764 \$217671 \$217765 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29539 VDD|pad|pin1|supply|vdd \$217763 \$218122 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29540 \$218122 d|z$59 \$217764 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29541 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217765
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29542 \$217766 \$217763 \$218154 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29543 VDD|pad|pin1|supply|vdd \$218634 \$218154 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29544 VDD|pad|pin1|supply|vdd \$217764 \$218414 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29545 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$218634
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29546 VDD|pad|pin1|supply|vdd \$217766 \$218634 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29547 \$218414 \$217671 \$217766 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29548 VDD|pad|pin1|supply|vdd \$218634 R[19]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29549 \$217768 \$217672 \$217769 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29550 \$217770 s|zn$2 \$217768 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29551 VDD|pad|pin1|supply|vdd R[20]|i0|q \$217770 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29552 \$217769 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29553 \$217672 s|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29554 VDD|pad|pin1|supply|vdd \$217768 d|z$40 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29555 VDD|pad|pin1|supply|vdd cp|z$4 \$217673 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29556 VDD|pad|pin1|supply|vdd \$217673 \$217771 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29557 VDD|pad|pin1|supply|vdd \$218415 \$217773 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29558 \$217772 \$217673 \$217773 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29559 VDD|pad|pin1|supply|vdd \$217771 \$218198 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29560 \$218198 d|z$60 \$217772 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29561 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217773
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29562 \$217774 \$217771 \$218231 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29563 VDD|pad|pin1|supply|vdd \$218635 \$218231 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29564 VDD|pad|pin1|supply|vdd \$217772 \$218415 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29565 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$218635
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29566 VDD|pad|pin1|supply|vdd \$217774 \$218635 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29567 \$218415 \$217673 \$217774 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29568 VDD|pad|pin1|supply|vdd \$218635 R[38]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29569 \$217776 \$217674 \$217777 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29570 \$217778 s|zn$3 \$217776 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29571 VDD|pad|pin1|supply|vdd i0|i1|q$1 \$217778 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29572 \$217777 R[51]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29573 \$217674 s|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29574 VDD|pad|pin1|supply|vdd \$217776 d|z$53 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29575 \$217780 \$217676 \$217781 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29576 \$217782 s|zn$3 \$217780 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29577 VDD|pad|pin1|supply|vdd i0|i1|q$6 \$217782 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29578 \$217781 R[49]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29579 \$217676 s|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29580 VDD|pad|pin1|supply|vdd \$217780 d|z$54 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29581 VDD|pad|pin1|supply|vdd cp|z$4 \$217677 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29582 VDD|pad|pin1|supply|vdd \$217677 \$217784 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29583 VDD|pad|pin1|supply|vdd \$218416 \$217786 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29584 \$217785 \$217677 \$217786 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29585 VDD|pad|pin1|supply|vdd \$217784 \$218302 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29586 \$218302 d|z$54 \$217785 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29587 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$217786
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29588 \$217787 \$217784 \$218341 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29589 VDD|pad|pin1|supply|vdd \$218636 \$218341 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29590 VDD|pad|pin1|supply|vdd \$217785 \$218416 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29591 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$218636
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29592 VDD|pad|pin1|supply|vdd \$217787 \$218636 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29593 \$218416 \$217677 \$217787 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29594 VDD|pad|pin1|supply|vdd \$218636 R[49]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29595 \$219901 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29596 VDD|pad|pin1|supply|vdd \$219901 \$219614 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29597 VDD|pad|pin1|supply|vdd \$219614 \$221513 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29598 \$221513 d|z$63 \$219902 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29599 \$219902 \$219901 \$221249 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29600 \$221249 \$219903 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29601 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$221249
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29602 \$219903 \$219902 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29603 \$219903 \$219901 \$219615 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29604 \$219615 \$219614 \$221532 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29605 VDD|pad|pin1|supply|vdd \$219905 \$221532 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29606 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$219905
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29607 VDD|pad|pin1|supply|vdd \$219615 \$219905 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29608 VDD|pad|pin1|supply|vdd \$219905 a2|q$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29609 \$219906 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29610 VDD|pad|pin1|supply|vdd \$219906 \$219616 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29611 VDD|pad|pin1|supply|vdd \$219616 \$221541 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29612 \$221541 d|z$52 \$219907 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29613 \$219907 \$219906 \$221250 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29614 \$221250 \$219908 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29615 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$221250
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29616 \$219908 \$219907 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29617 \$219908 \$219906 \$219617 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29618 \$219617 \$219616 \$221552 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29619 VDD|pad|pin1|supply|vdd \$219910 \$221552 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29620 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$219910
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29621 VDD|pad|pin1|supply|vdd \$219617 \$219910 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29622 VDD|pad|pin1|supply|vdd \$219910 a1|a2|q$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29623 \$219912 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29624 VDD|pad|pin1|supply|vdd \$219912 \$219618 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29625 VDD|pad|pin1|supply|vdd \$219618 \$221561 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29626 \$221561 d|z$64 \$219913 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29627 \$219913 \$219912 \$221251 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29628 \$221251 \$219914 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29629 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$221251
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29630 \$219914 \$219913 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29631 \$219914 \$219912 \$219619 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29632 \$219619 \$219618 \$221553 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29633 VDD|pad|pin1|supply|vdd \$219916 \$221553 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29634 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$219916
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29635 VDD|pad|pin1|supply|vdd \$219619 \$219916 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29636 VDD|pad|pin1|supply|vdd \$219916 a1|a2|b|q|s VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29637 \$219919 \$219620 \$219918 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29638 \$219919 DATA|core|i0|i1|p2c VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p
+ PS=1.93u PD=1.93u
M$29639 VDD|pad|pin1|supply|vdd a1|i0|q \$219920 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29640 \$219920 d|s|z \$219918 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29641 VDD|pad|pin1|supply|vdd d|s|z \$219620 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29642 VDD|pad|pin1|supply|vdd \$219918 d|z$41 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29643 VDD|pad|pin1|supply|vdd a1|a2|q$5 \$219921 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29644 \$219921 a1|i0|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29645 a1|a2|a4|z \$219921 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29646 \$219923 \$219621 \$219922 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29647 \$219923 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29648 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q \$219924 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29649 \$219924 s|zn$1 \$219922 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29650 VDD|pad|pin1|supply|vdd s|zn$1 \$219621 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29651 VDD|pad|pin1|supply|vdd \$219922 d|z$46 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29652 \$219926 \$219622 \$219925 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29653 \$219926 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29654 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q \$219927 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29655 \$219927 s|zn$1 \$219925 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29656 VDD|pad|pin1|supply|vdd s|zn$1 \$219622 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29657 VDD|pad|pin1|supply|vdd \$219925 d|z$55 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29658 s|zn$4 a1|zn$2 \$221599 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29659 \$221599 a2|zn$11 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29660 a2|a3|zn$1 a1|i|i0|i1|q \$221598 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29661 \$221598 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29662 \$219929 \$219623 \$219928 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29663 \$219929 R[50]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29664 VDD|pad|pin1|supply|vdd i0|i1|q$2 \$219930 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29665 \$219930 s|zn$3 \$219928 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29666 VDD|pad|pin1|supply|vdd s|zn$3 \$219623 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29667 VDD|pad|pin1|supply|vdd \$219928 d|z$56 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29668 \$219931 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29669 VDD|pad|pin1|supply|vdd \$219931 \$219624 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29670 VDD|pad|pin1|supply|vdd \$219624 \$221607 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29671 \$221607 d|z$65 \$219932 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29672 \$219932 \$219931 \$221252 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29673 \$221252 \$219933 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29674 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$221252
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29675 \$219933 \$219932 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29676 \$219933 \$219931 \$219625 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29677 \$219625 \$219624 \$221612 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29678 VDD|pad|pin1|supply|vdd \$219935 \$221612 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29679 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$219935
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29680 VDD|pad|pin1|supply|vdd \$219625 \$219935 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29681 VDD|pad|pin1|supply|vdd \$219935 R[54]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29682 VDD|pad|pin1|supply|vdd a1|a2|a4|z s|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29683 s|zn a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29684 s|zn a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29685 VDD|pad|pin1|supply|vdd a2|z$9 \$219937 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29686 \$219937 a1|a2|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29687 s|z \$219937 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29688 \$219939 \$219627 \$219938 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29689 \$219939 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29690 VDD|pad|pin1|supply|vdd R[31]|i0|q \$219940 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29691 \$219940 s|z \$219938 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29692 VDD|pad|pin1|supply|vdd s|z \$219627 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29693 VDD|pad|pin1|supply|vdd \$219938 d|z$57 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29694 \$219942 \$219628 \$219941 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29695 \$219942 R[52]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29696 VDD|pad|pin1|supply|vdd i0|i1|q$5 \$219943 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29697 \$219943 s|zn$3 \$219941 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29698 VDD|pad|pin1|supply|vdd s|zn$3 \$219628 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29699 VDD|pad|pin1|supply|vdd \$219941 d|z$61 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29700 \$219946 \$219629 \$219945 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29701 \$219946 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29702 VDD|pad|pin1|supply|vdd R[23]|i0|q \$219947 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29703 \$219947 s|zn$2 \$219945 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29704 VDD|pad|pin1|supply|vdd s|zn$2 \$219629 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29705 VDD|pad|pin1|supply|vdd \$219945 d|z$48 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29706 \$219949 \$219630 \$219948 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29707 \$219949 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29708 VDD|pad|pin1|supply|vdd R[17]|i0|q \$219950 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29709 \$219950 s|zn$2 \$219948 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29710 VDD|pad|pin1|supply|vdd s|zn$2 \$219630 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29711 VDD|pad|pin1|supply|vdd \$219948 d|z$58 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29712 \$219952 \$219631 \$219951 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29713 \$219952 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29714 VDD|pad|pin1|supply|vdd R[16]|i0|q \$219953 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29715 \$219953 s|zn$2 \$219951 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29716 VDD|pad|pin1|supply|vdd s|zn$2 \$219631 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29717 VDD|pad|pin1|supply|vdd \$219951 d|z$62 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29718 \$219955 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29719 VDD|pad|pin1|supply|vdd \$219955 \$219632 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29720 VDD|pad|pin1|supply|vdd \$219632 \$221632 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29721 \$221632 d|z$62 \$219956 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29722 \$219956 \$219955 \$221253 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29723 \$221253 \$219957 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29724 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$221253
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29725 \$219957 \$219956 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29726 \$219957 \$219955 \$219633 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29727 \$219633 \$219632 \$221629 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29728 VDD|pad|pin1|supply|vdd \$219959 \$221629 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29729 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$219959
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29730 VDD|pad|pin1|supply|vdd \$219633 \$219959 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29731 VDD|pad|pin1|supply|vdd \$219959 R[16]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29732 \$219961 \$219634 \$219960 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29733 \$219961 R[38]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29734 VDD|pad|pin1|supply|vdd i0|i1|q$3 \$219962 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29735 \$219962 s|zn \$219960 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29736 VDD|pad|pin1|supply|vdd s|zn \$219634 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29737 VDD|pad|pin1|supply|vdd \$219960 d|z$60 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29738 \$219963 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29739 VDD|pad|pin1|supply|vdd \$219963 \$219635 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29740 VDD|pad|pin1|supply|vdd \$219635 \$221661 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29741 \$221661 d|z$66 \$219964 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29742 \$219964 \$219963 \$221254 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29743 \$221254 \$219965 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29744 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$221254
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29745 \$219965 \$219964 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29746 \$219965 \$219963 \$219636 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29747 \$219636 \$219635 \$221651 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29748 VDD|pad|pin1|supply|vdd \$219967 \$221651 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29749 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$219967
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29750 VDD|pad|pin1|supply|vdd \$219636 \$219967 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29751 VDD|pad|pin1|supply|vdd \$219967 R[48]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29752 \$219969 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29753 VDD|pad|pin1|supply|vdd \$219969 \$219637 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29754 VDD|pad|pin1|supply|vdd \$219637 \$221664 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29755 \$221664 d|z$53 \$219970 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29756 \$219970 \$219969 \$221255 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29757 \$221255 \$219971 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29758 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$221255
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29759 \$219971 \$219970 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29760 \$219971 \$219969 \$219638 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29761 \$219638 \$219637 \$221673 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29762 VDD|pad|pin1|supply|vdd \$219973 \$221673 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29763 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$219973
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29764 VDD|pad|pin1|supply|vdd \$219638 \$219973 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29765 VDD|pad|pin1|supply|vdd \$219973 R[51]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29766 \$219974 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29767 VDD|pad|pin1|supply|vdd \$219974 \$219639 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29768 VDD|pad|pin1|supply|vdd \$219639 \$221680 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29769 \$221680 d|z$67 \$219975 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29770 \$219975 \$219974 \$221256 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29771 \$221256 \$219976 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29772 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$221256
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29773 \$219976 \$219975 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29774 \$219976 \$219974 \$219640 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29775 \$219640 \$219639 \$221691 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29776 VDD|pad|pin1|supply|vdd \$219978 \$221691 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29777 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$219978
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29778 VDD|pad|pin1|supply|vdd \$219640 \$219978 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29779 VDD|pad|pin1|supply|vdd \$219978 R[55]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29780 \$219981 \$219641 \$219980 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29781 \$219981 R[53]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29782 VDD|pad|pin1|supply|vdd i0|i1|q$7 \$219982 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29783 \$219982 s|zn$3 \$219980 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29784 VDD|pad|pin1|supply|vdd s|zn$3 \$219641 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29785 VDD|pad|pin1|supply|vdd \$219980 d|z$51 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29786 \$223949 \$223834 \$223948 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29787 \$223949 i0|i1|q$9 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29788 VDD|pad|pin1|supply|vdd i0|i1|q$8 \$223951 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29789 \$223951 a2|i|s|zn \$223948 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29790 VDD|pad|pin1|supply|vdd a1|a2|q$8 \$222044 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29791 VDD|pad|pin1|supply|vdd a1|b|d|z \$222044 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29792 \$223954 \$223835 \$223953 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29793 \$223954 i1|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29794 VDD|pad|pin1|supply|vdd i0|z$1 \$223956 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29795 \$223956 a1|a2|b|q|s \$223953 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29796 VDD|pad|pin1|supply|vdd \$222044 d|z$63 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29797 a3|zn$2 a1|a2|q$8 \$222730 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29798 \$222730 a2|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29799 z$33 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29800 cp|i|z$5 \$223959 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$29801 VDD|pad|pin1|supply|vdd i|z$115 \$223959 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$29802 VDD|pad|pin1|supply|vdd a1|a2|q$9 \$222046 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29803 VDD|pad|pin1|supply|vdd a1|b|d|z \$222046 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29804 VDD|pad|pin1|supply|vdd \$222046 d|z$64 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29805 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$225348
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29806 \$223962 \$223961 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29807 \$223962 \$223960 \$223837 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29808 \$223837 \$223836 \$225508 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29809 VDD|pad|pin1|supply|vdd \$223964 \$225508 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29810 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$223964
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29811 VDD|pad|pin1|supply|vdd \$223837 \$223964 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29812 VDD|pad|pin1|supply|vdd \$223964 a2|q$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29813 \$222022 \$221966 \$222047 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29814 \$222048 a1|a2|b|q|s \$222022 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29815 VDD|pad|pin1|supply|vdd i0|z \$222048 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29816 \$222047 i1|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29817 \$221966 a1|a2|b|q|s VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29818 VDD|pad|pin1|supply|vdd \$222022 d|z$68 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29819 a4|zn$2 a1|a2|q$9 \$222734 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29820 \$222734 a1|a2|b|q|s VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29821 VDD|pad|pin1|supply|vdd a2|q$8 \$223966 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29822 \$223966 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29823 DOUT_EN|z \$223966 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29824 d|s|zn CEB|a1|core|i|p2c \$222733 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29825 \$222733 a1|a2|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29826 a1|b|d|z CEB|a1|core|i|p2c VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p
+ PS=3.33u PD=3.33u
M$29827 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$225349
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29828 \$223970 \$223969 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29829 \$223970 \$223968 \$223839 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29830 \$223839 \$223838 \$225552 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29831 VDD|pad|pin1|supply|vdd \$223972 \$225552 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29832 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$223972
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29833 VDD|pad|pin1|supply|vdd \$223839 \$223972 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29834 VDD|pad|pin1|supply|vdd \$223972 R[7]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29835 VDD|pad|pin1|supply|vdd a1|a2|q$5 a1|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29836 VDD|pad|pin1|supply|vdd a1|i0|q$1 a1|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29837 \$222023 \$221967 \$222051 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29838 \$222052 s|z$1 \$222023 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29839 VDD|pad|pin1|supply|vdd R[7]|i|i0|q \$222052 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29840 \$222051 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29841 \$221967 s|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29842 VDD|pad|pin1|supply|vdd \$222023 d|z$69 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29843 VDD|pad|pin1|supply|vdd i|z$115 \$222024 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$29844 VDD|pad|pin1|supply|vdd \$222024 cp|i|z$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$29845 \$222025 \$221969 \$222054 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29846 \$222055 s|zn$4 \$222025 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29847 VDD|pad|pin1|supply|vdd R[47]|i0|q \$222055 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29848 \$222054 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29849 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$225350
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29850 \$223975 \$223974 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29851 \$223975 \$223973 \$223841 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29852 \$223841 \$223840 \$225567 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29853 VDD|pad|pin1|supply|vdd \$223977 \$225567 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29854 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$223977
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29855 VDD|pad|pin1|supply|vdd \$223841 \$223977 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29856 VDD|pad|pin1|supply|vdd \$223977 R[47]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29857 \$221969 s|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29858 VDD|pad|pin1|supply|vdd \$222025 d|z$70 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29859 z$32 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29860 a2|z$12 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29861 \$222058 a1|zn$14 \$222736 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29862 VDD|pad|pin1|supply|vdd a2|zn$32 \$222736 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$29863 VDD|pad|pin1|supply|vdd \$222058 i1|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$29864 VDD|pad|pin1|supply|vdd a2|z$10 \$223978 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29865 \$223978 a1|a2|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29866 s|z$1 \$223978 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29867 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a2|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29868 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29869 VDD|pad|pin1|supply|vdd a2|a3|zn$1 \$223979 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29870 \$223979 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29871 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29872 a2|z$10 \$223979 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29873 s|zn$5 a1|zn$2 \$225590 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29874 \$225590 a2|zn$13 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29875 s|zn$2 a1|zn$2 \$222735 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29876 \$222735 a2|zn$12 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29877 a1|a3|z a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29878 \$222026 \$221971 \$222061 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29879 \$222062 s|zn$3 \$222026 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29880 VDD|pad|pin1|supply|vdd i0|i1|q$3 \$222062 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29881 \$222061 R[54]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29882 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$225351
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29883 \$223983 \$223982 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29884 \$223983 \$223980 \$223843 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29885 \$223843 \$223842 \$225653 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29886 VDD|pad|pin1|supply|vdd \$223985 \$225653 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29887 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$223985
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29888 VDD|pad|pin1|supply|vdd \$223843 \$223985 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29889 VDD|pad|pin1|supply|vdd \$223985 R[43]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29890 \$221971 s|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29891 VDD|pad|pin1|supply|vdd \$222026 d|z$65 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29892 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q s|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29893 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q s|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$29894 VDD|pad|pin1|supply|vdd a1|z$15 s|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$29895 VDD|pad|pin1|supply|vdd a1|a2|a4|z s|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29896 s|zn$6 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29897 VDD|pad|pin1|supply|vdd a1|a2|a4|z s|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29898 VDD|pad|pin1|supply|vdd a2|a3|z$1 \$222063 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29899 VDD|pad|pin1|supply|vdd a1|a3|z \$222063 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29900 s|zn$6 a2|a3|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29901 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q \$223986 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29902 \$223986 a1|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29903 VDD|pad|pin1|supply|vdd \$222063 a2|z$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29904 VDD|pad|pin1|supply|vdd CLK|core|i|p2c$1 \$222027
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$29905 VDD|pad|pin1|supply|vdd \$222027 i|z$115 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$29906 a2|a3|z$1 \$223986 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29907 VDD|pad|pin1|supply|vdd cp|i|z$7 \$222028 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29908 VDD|pad|pin1|supply|vdd \$222028 \$222029 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29909 VDD|pad|pin1|supply|vdd \$222726 \$222030 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29910 \$222064 \$222028 \$222030 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29911 VDD|pad|pin1|supply|vdd \$222029 \$222413 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29912 \$222413 d|z$61 \$222064 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29913 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$222030
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29914 \$222031 \$222029 \$222455 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29915 VDD|pad|pin1|supply|vdd \$222738 \$222455 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29916 VDD|pad|pin1|supply|vdd \$222064 \$222726 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29917 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$222738
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29918 VDD|pad|pin1|supply|vdd \$222031 \$222738 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29919 \$222726 \$222028 \$222031 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29920 VDD|pad|pin1|supply|vdd \$222738 R[52]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29921 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$225352
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29922 \$223989 \$223988 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29923 \$223989 \$223987 \$223846 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29924 \$223846 \$223845 \$225692 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29925 VDD|pad|pin1|supply|vdd \$223991 \$225692 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29926 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$223991
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29927 VDD|pad|pin1|supply|vdd \$223846 \$223991 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29928 VDD|pad|pin1|supply|vdd \$223991 R[46]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29929 \$222032 \$221972 \$222065 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29930 \$222066 s|zn$5 \$222032 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29931 VDD|pad|pin1|supply|vdd R[15]|i|i0|q \$222066 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29932 \$222065 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29933 \$221972 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29934 VDD|pad|pin1|supply|vdd \$222032 d|z$71 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29935 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$225353
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29936 \$223995 \$223994 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29937 \$223995 \$223993 \$223848 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29938 \$223848 \$223847 \$225764 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29939 VDD|pad|pin1|supply|vdd \$223997 \$225764 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29940 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$223997
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29941 VDD|pad|pin1|supply|vdd \$223848 \$223997 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29942 VDD|pad|pin1|supply|vdd \$223997 R[15]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29943 \$222033 \$221974 \$222068 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29944 \$222069 s|zn$2 \$222033 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29945 VDD|pad|pin1|supply|vdd R[19]|i0|q \$222069 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29946 \$222068 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29947 \$221974 s|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29948 VDD|pad|pin1|supply|vdd \$222033 d|z$59 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29949 \$222034 \$221975 \$222070 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29950 \$222071 s|zn$5 \$222034 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29951 VDD|pad|pin1|supply|vdd R[12]|i|i0|q \$222071 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29952 \$222070 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29953 \$221975 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29954 VDD|pad|pin1|supply|vdd \$222034 d|z$72 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29955 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$225354
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29956 \$224000 \$223999 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29957 \$224000 \$223998 \$223850 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29958 \$223850 \$223849 \$225810 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29959 VDD|pad|pin1|supply|vdd \$224002 \$225810 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29960 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$224002
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29961 VDD|pad|pin1|supply|vdd \$223850 \$224002 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29962 VDD|pad|pin1|supply|vdd \$224002 R[12]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29963 \$222035 \$221976 \$222073 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29964 \$222074 s|z$1 \$222035 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29965 VDD|pad|pin1|supply|vdd R[4]|i|i0|q \$222074 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29966 \$222073 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29967 \$221976 s|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29968 VDD|pad|pin1|supply|vdd \$222035 d|z$73 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29969 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$225355
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29970 \$224005 \$224004 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29971 \$224005 \$224003 \$223852 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29972 \$223852 \$223851 \$225818 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29973 VDD|pad|pin1|supply|vdd \$224007 \$225818 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29974 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$224007
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29975 VDD|pad|pin1|supply|vdd \$223852 \$224007 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29976 VDD|pad|pin1|supply|vdd \$224007 R[4]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29977 \$222036 \$221977 \$222076 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29978 \$222077 s|zn$3 \$222036 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29979 VDD|pad|pin1|supply|vdd i0|i1|q \$222077 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29980 \$222076 R[48]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29981 \$221977 s|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29982 VDD|pad|pin1|supply|vdd \$222036 d|z$66 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29983 \$222037 \$221978 \$222078 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29984 \$222079 s|zn$4 \$222037 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29985 VDD|pad|pin1|supply|vdd R[44]|i0|q \$222079 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29986 \$222078 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29987 \$221978 s|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29988 VDD|pad|pin1|supply|vdd \$222037 d|z$74 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29989 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$225356
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29990 \$224010 \$224009 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29991 \$224010 \$224008 \$223854 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29992 \$223854 \$223853 \$225878 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29993 VDD|pad|pin1|supply|vdd \$224012 \$225878 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29994 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$224012
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29995 VDD|pad|pin1|supply|vdd \$223854 \$224012 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29996 VDD|pad|pin1|supply|vdd \$224012 R[44]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29997 \$222038 \$221979 \$222081 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29998 \$222082 s|zn$3 \$222038 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29999 VDD|pad|pin1|supply|vdd i0|i1|q$4 \$222082 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30000 \$222081 R[55]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30001 cp|z$4 \$224013 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$30002 VDD|pad|pin1|supply|vdd i|z$115 \$224013 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$30003 \$221979 s|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30004 VDD|pad|pin1|supply|vdd \$222038 d|z$67 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30005 \$222039 \$221980 \$222083 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30006 \$222084 s|zn$6 \$222039 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30007 VDD|pad|pin1|supply|vdd i0|i1|q$4 \$222084 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30008 \$222083 R[63]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30009 \$224015 \$223855 \$224014 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30010 \$224015 R[60]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30011 VDD|pad|pin1|supply|vdd i0|i1|q$5 \$224016 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30012 \$224016 s|zn$6 \$224014 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30013 \$221980 s|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30014 VDD|pad|pin1|supply|vdd \$222039 d|z$75 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30015 VDD|pad|pin1|supply|vdd cp|z$4 \$222040 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30016 VDD|pad|pin1|supply|vdd \$222040 \$222041 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30017 VDD|pad|pin1|supply|vdd \$222729 \$222042 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30018 \$222086 \$222040 \$222042 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30019 VDD|pad|pin1|supply|vdd \$222041 \$222680 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30020 \$222680 d|z$75 \$222086 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30021 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$222042
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30022 \$222043 \$222041 \$222706 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30023 VDD|pad|pin1|supply|vdd \$222739 \$222706 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30024 VDD|pad|pin1|supply|vdd \$222086 \$222729 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30025 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$222739
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30026 VDD|pad|pin1|supply|vdd \$222043 \$222739 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30027 \$222729 \$222040 \$222043 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30028 VDD|pad|pin1|supply|vdd \$222739 R[63]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30029 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$225357
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30030 \$224020 \$224019 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30031 \$224020 \$224018 \$223857 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30032 \$223857 \$223856 \$225917 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30033 VDD|pad|pin1|supply|vdd \$224022 \$225917 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30034 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$224022
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30035 VDD|pad|pin1|supply|vdd \$223857 \$224022 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30036 VDD|pad|pin1|supply|vdd \$224022 R[60]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30037 VDD|pad|pin1|supply|vdd a2|i|s|zn \$223834 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30038 VDD|pad|pin1|supply|vdd \$223948 i0|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30039 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$223835 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30040 VDD|pad|pin1|supply|vdd \$223953 d|z$76 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30041 \$223960 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30042 VDD|pad|pin1|supply|vdd \$223960 \$223836 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30043 VDD|pad|pin1|supply|vdd \$223836 \$225481 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30044 \$225481 a2|d|z \$223961 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30045 \$223961 \$223960 \$225348 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30046 \$225348 \$223962 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30047 \$223968 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30048 VDD|pad|pin1|supply|vdd \$223968 \$223838 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30049 VDD|pad|pin1|supply|vdd \$223838 \$225524 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30050 \$225524 d|z$69 \$223969 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30051 \$223969 \$223968 \$225349 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30052 \$225349 \$223970 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30053 \$223973 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30054 VDD|pad|pin1|supply|vdd \$223973 \$223840 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30055 VDD|pad|pin1|supply|vdd \$223840 \$225581 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30056 \$225581 d|z$70 \$223974 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30057 \$223974 \$223973 \$225350 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30058 \$225350 \$223975 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30059 \$223980 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30060 VDD|pad|pin1|supply|vdd \$223980 \$223842 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30061 VDD|pad|pin1|supply|vdd \$223842 \$225620 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30062 \$225620 d|z$78 \$223982 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30063 \$223982 \$223980 \$225351 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30064 \$225351 \$223983 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30065 \$223987 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30066 VDD|pad|pin1|supply|vdd \$223987 \$223845 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30067 VDD|pad|pin1|supply|vdd \$223845 \$225706 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30068 \$225706 d|z$79 \$223988 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30069 \$223988 \$223987 \$225352 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30070 \$225352 \$223989 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30071 \$223993 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30072 VDD|pad|pin1|supply|vdd \$223993 \$223847 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30073 VDD|pad|pin1|supply|vdd \$223847 \$225721 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30074 \$225721 d|z$71 \$223994 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30075 \$223994 \$223993 \$225353 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30076 \$225353 \$223995 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30077 \$223998 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30078 VDD|pad|pin1|supply|vdd \$223998 \$223849 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30079 VDD|pad|pin1|supply|vdd \$223849 \$225778 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30080 \$225778 d|z$72 \$223999 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30081 \$223999 \$223998 \$225354 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30082 \$225354 \$224000 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30083 \$224003 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30084 VDD|pad|pin1|supply|vdd \$224003 \$223851 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30085 VDD|pad|pin1|supply|vdd \$223851 \$225832 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30086 \$225832 d|z$73 \$224004 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30087 \$224004 \$224003 \$225355 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30088 \$225355 \$224005 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30089 \$224008 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30090 VDD|pad|pin1|supply|vdd \$224008 \$223853 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30091 VDD|pad|pin1|supply|vdd \$223853 \$225845 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30092 \$225845 d|z$74 \$224009 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30093 \$224009 \$224008 \$225356 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30094 \$225356 \$224010 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30095 VDD|pad|pin1|supply|vdd s|zn$6 \$223855 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30096 VDD|pad|pin1|supply|vdd \$224014 d|z$77 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30097 \$224018 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30098 VDD|pad|pin1|supply|vdd \$224018 \$223856 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30099 VDD|pad|pin1|supply|vdd \$223856 \$225915 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30100 \$225915 d|z$77 \$224019 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30101 \$224019 \$224018 \$225357 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30102 \$225357 \$224020 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30103 VDD|pad|pin1|supply|vdd cp|i|z$5 \$226128 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30104 VDD|pad|pin1|supply|vdd \$226128 \$226129 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30105 VDD|pad|pin1|supply|vdd \$226405 \$226130 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30106 \$226203 \$226128 \$226130 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30107 VDD|pad|pin1|supply|vdd \$226129 \$226347 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30108 \$226347 d|z$76 \$226203 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30109 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226130
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30110 \$226131 \$226129 \$226345 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30111 VDD|pad|pin1|supply|vdd \$226406 \$226345 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30112 VDD|pad|pin1|supply|vdd \$226203 \$226405 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30113 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226406
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30114 VDD|pad|pin1|supply|vdd \$226131 \$226406 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30115 \$226405 \$226128 \$226131 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30116 VDD|pad|pin1|supply|vdd \$226406 i0|i1|q$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30117 VDD|pad|pin1|supply|vdd cp|i|z$5 \$226132 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30118 VDD|pad|pin1|supply|vdd \$226132 \$226133 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30119 VDD|pad|pin1|supply|vdd \$226407 \$226134 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30120 \$226204 \$226132 \$226134 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30121 VDD|pad|pin1|supply|vdd \$226133 \$226348 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30122 \$226348 d|z$68 \$226204 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30123 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226134
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30124 \$226135 \$226133 \$226349 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30125 VDD|pad|pin1|supply|vdd \$226408 \$226349 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30126 VDD|pad|pin1|supply|vdd \$226204 \$226407 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30127 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226408
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30128 VDD|pad|pin1|supply|vdd \$226135 \$226408 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30129 \$226407 \$226132 \$226135 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30130 VDD|pad|pin1|supply|vdd \$226408 i0|i1|q$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30131 VDD|pad|pin1|supply|vdd cp|i|z$6 \$226136 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30132 VDD|pad|pin1|supply|vdd \$226136 \$226137 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30133 VDD|pad|pin1|supply|vdd \$226409 \$226138 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30134 \$226205 \$226136 \$226138 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30135 VDD|pad|pin1|supply|vdd \$226137 \$226351 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30136 \$226351 d|z$84 \$226205 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30137 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226138
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30138 \$226139 \$226137 \$226352 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30139 VDD|pad|pin1|supply|vdd \$226410 \$226352 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30140 VDD|pad|pin1|supply|vdd \$226205 \$226409 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30141 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226410
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30142 VDD|pad|pin1|supply|vdd \$226139 \$226410 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30143 \$226409 \$226136 \$226139 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30144 VDD|pad|pin1|supply|vdd \$226410 i0|i1|q$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30145 VDD|pad|pin1|supply|vdd cp|i|z$6 \$226140 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30146 VDD|pad|pin1|supply|vdd \$226140 \$226141 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30147 VDD|pad|pin1|supply|vdd \$226411 \$226142 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30148 \$226207 \$226140 \$226142 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30149 VDD|pad|pin1|supply|vdd \$226141 \$226356 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30150 \$226356 d|z$80 \$226207 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30151 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226142
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30152 \$226143 \$226141 \$226354 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30153 VDD|pad|pin1|supply|vdd \$226412 \$226354 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30154 VDD|pad|pin1|supply|vdd \$226207 \$226411 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30155 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226412
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30156 VDD|pad|pin1|supply|vdd \$226143 \$226412 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30157 \$226411 \$226140 \$226143 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30158 VDD|pad|pin1|supply|vdd \$226412 DUT_Footer|R[10]|Vdn|i|i0|q
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p
+ PS=2.67u PD=3.33u
M$30159 \$226144 \$226113 \$226208 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30160 \$226209 s|zn$5 \$226144 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30161 VDD|pad|pin1|supply|vdd DUT_Footer|R[10]|Vdn|i|i0|q \$226209
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p
+ PS=1.93u PD=1.74u
M$30162 \$226208 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30163 \$226113 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30164 VDD|pad|pin1|supply|vdd \$226144 d|z$80 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30165 VDD|pad|pin1|supply|vdd a2|z$12 a2|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30166 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30167 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30168 \$226145 \$226114 \$226212 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30169 \$226213 s|z$1 \$226145 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30170 VDD|pad|pin1|supply|vdd DUT_Header|R[3]|Vup|i|i0|q \$226213
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p
+ PS=1.93u PD=1.74u
M$30171 \$226212 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30172 \$226114 s|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30173 VDD|pad|pin1|supply|vdd \$226145 d|z$81 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30174 \$226146 \$226115 \$226215 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30175 \$226216 s|zn$5 \$226146 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30176 VDD|pad|pin1|supply|vdd R[14]|i|i0|q \$226216 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30177 \$226215 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30178 \$226115 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30179 VDD|pad|pin1|supply|vdd \$226146 d|z$82 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30180 VDD|pad|pin1|supply|vdd cp|i|z$6 \$226147 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30181 VDD|pad|pin1|supply|vdd \$226147 \$226148 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30182 VDD|pad|pin1|supply|vdd \$226415 \$226149 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30183 \$226218 \$226147 \$226149 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30184 VDD|pad|pin1|supply|vdd \$226148 \$226360 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30185 \$226360 d|z$82 \$226218 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30186 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226149
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30187 \$226150 \$226148 \$226361 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30188 VDD|pad|pin1|supply|vdd \$226416 \$226361 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30189 VDD|pad|pin1|supply|vdd \$226218 \$226415 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30190 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226416
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30191 VDD|pad|pin1|supply|vdd \$226150 \$226416 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30192 \$226415 \$226147 \$226150 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30193 VDD|pad|pin1|supply|vdd \$226416 R[14]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30194 a1|z$15 a1|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$30195 \$226219 a1|zn$20 \$226676 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30196 VDD|pad|pin1|supply|vdd a2|zn$14 \$226676 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30197 VDD|pad|pin1|supply|vdd \$226219 i1|z$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30198 \$226151 \$226116 \$226221 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30199 \$226222 s|zn$4 \$226151 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30200 VDD|pad|pin1|supply|vdd R[46]|i0|q \$226222 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30201 \$226221 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30202 \$226116 s|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30203 VDD|pad|pin1|supply|vdd \$226151 d|z$79 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30204 VDD|pad|pin1|supply|vdd cp|i|z$7 \$226152 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30205 VDD|pad|pin1|supply|vdd \$226152 \$226153 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30206 VDD|pad|pin1|supply|vdd \$226417 \$226154 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30207 \$226223 \$226152 \$226154 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30208 VDD|pad|pin1|supply|vdd \$226153 \$226394 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30209 \$226394 d|z$85 \$226223 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30210 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226154
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30211 \$226155 \$226153 \$226397 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30212 VDD|pad|pin1|supply|vdd \$226418 \$226397 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30213 VDD|pad|pin1|supply|vdd \$226223 \$226417 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30214 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226418
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30215 VDD|pad|pin1|supply|vdd \$226155 \$226418 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30216 \$226417 \$226152 \$226155 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30217 VDD|pad|pin1|supply|vdd \$226418 RO_control|R[1]|i|i0|nclk|q
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p
+ PS=2.67u PD=3.33u
M$30218 VDD|pad|pin1|supply|vdd cp|i|z$7 \$226156 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30219 VDD|pad|pin1|supply|vdd \$226156 \$226157 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30220 VDD|pad|pin1|supply|vdd \$226419 \$226158 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30221 \$226225 \$226156 \$226158 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30222 VDD|pad|pin1|supply|vdd \$226157 \$226399 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30223 \$226399 d|z$86 \$226225 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30224 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226158
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30225 \$226159 \$226157 \$226403 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30226 VDD|pad|pin1|supply|vdd \$226420 \$226403 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30227 VDD|pad|pin1|supply|vdd \$226225 \$226419 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30228 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226420
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30229 VDD|pad|pin1|supply|vdd \$226159 \$226420 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30230 \$226419 \$226156 \$226159 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30231 VDD|pad|pin1|supply|vdd \$226420 DUT_Header|R[11]|Vup|i|i0|q
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p
+ PS=2.67u PD=3.33u
M$30232 \$226160 \$226117 \$226226 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30233 \$226227 s|z$1 \$226160 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30234 VDD|pad|pin1|supply|vdd R[0]|clk|i|i0|n_RO_control|q \$226227
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p
+ PS=1.93u PD=1.74u
M$30235 \$226226 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30236 \$226117 s|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30237 VDD|pad|pin1|supply|vdd \$226160 d|z$83 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30238 VDD|pad|pin1|supply|vdd cp|i|z$7 \$226161 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30239 VDD|pad|pin1|supply|vdd \$226161 \$226162 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30240 VDD|pad|pin1|supply|vdd \$226422 \$226163 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30241 \$226229 \$226161 \$226163 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30242 VDD|pad|pin1|supply|vdd \$226162 \$226401 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30243 \$226401 d|z$87 \$226229 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30244 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226163
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30245 \$226164 \$226162 \$226398 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30246 VDD|pad|pin1|supply|vdd \$226423 \$226398 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30247 VDD|pad|pin1|supply|vdd \$226229 \$226422 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30248 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226423
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30249 VDD|pad|pin1|supply|vdd \$226164 \$226423 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30250 \$226422 \$226161 \$226164 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30251 VDD|pad|pin1|supply|vdd \$226423 R[8]|clk|i|i0|n_RO_control|q
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p
+ PS=2.67u PD=3.33u
M$30252 VDD|pad|pin1|supply|vdd cp|z$4 \$226165 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30253 VDD|pad|pin1|supply|vdd \$226165 \$226166 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30254 VDD|pad|pin1|supply|vdd \$226424 \$226167 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30255 \$226230 \$226165 \$226167 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30256 VDD|pad|pin1|supply|vdd \$226166 \$226396 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30257 \$226396 d|z$88 \$226230 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30258 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226167
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30259 \$226168 \$226166 \$226395 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30260 VDD|pad|pin1|supply|vdd \$226425 \$226395 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30261 VDD|pad|pin1|supply|vdd \$226230 \$226424 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30262 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226425
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30263 VDD|pad|pin1|supply|vdd \$226168 \$226425 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30264 \$226424 \$226165 \$226168 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30265 VDD|pad|pin1|supply|vdd \$226425 R[40]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30266 VDD|pad|pin1|supply|vdd cp|z$4 \$226169 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30267 VDD|pad|pin1|supply|vdd \$226169 \$226170 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30268 VDD|pad|pin1|supply|vdd \$226426 \$226171 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30269 \$226231 \$226169 \$226171 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30270 VDD|pad|pin1|supply|vdd \$226170 \$226390 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30271 \$226390 d|z$89 \$226231 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30272 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226171
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30273 \$226172 \$226170 \$226393 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30274 VDD|pad|pin1|supply|vdd \$226427 \$226393 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30275 VDD|pad|pin1|supply|vdd \$226231 \$226426 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30276 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$226427
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30277 VDD|pad|pin1|supply|vdd \$226172 \$226427 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30278 \$226426 \$226169 \$226172 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30279 VDD|pad|pin1|supply|vdd \$226427 R[59]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30280 VDD|pad|pin1|supply|vdd \$226404 RESET_B|RSTB|core|p2c
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$30281 \$227910 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30282 VDD|pad|pin1|supply|vdd \$227910 \$227880 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30283 VDD|pad|pin1|supply|vdd \$227880 \$229270 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30284 \$229270 d|z$90 \$227911 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30285 \$227911 \$227910 \$229158 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30286 \$229158 \$227913 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30287 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$229158
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30288 \$227913 \$227911 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30289 \$227913 \$227910 \$227881 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30290 \$227881 \$227880 \$229285 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30291 VDD|pad|pin1|supply|vdd \$227915 \$229285 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30292 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$227915
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30293 VDD|pad|pin1|supply|vdd \$227881 \$227915 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30294 VDD|pad|pin1|supply|vdd \$227915 i0|i1|q$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30295 \$227918 \$227882 \$227917 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30296 \$227918 i0|i1|q$11 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30297 VDD|pad|pin1|supply|vdd i0|i1|q$9 \$227919 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30298 \$227919 a2|i|s|zn \$227917 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30299 VDD|pad|pin1|supply|vdd a2|i|s|zn \$227882 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30300 VDD|pad|pin1|supply|vdd \$227917 i0|z$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30301 \$227922 \$227883 \$227921 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30302 \$227922 i1|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30303 VDD|pad|pin1|supply|vdd i0|z$2 \$227923 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30304 \$227923 a1|a2|b|q|s \$227921 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30305 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$227883 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30306 VDD|pad|pin1|supply|vdd \$227921 d|z$90 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30307 \$227925 \$227884 \$227924 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30308 \$227925 i0|i1|q$8 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30309 VDD|pad|pin1|supply|vdd i0|i1|q$10 \$227926 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30310 \$227926 a2|i|s|zn \$227924 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30311 VDD|pad|pin1|supply|vdd a2|i|s|zn \$227884 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30312 VDD|pad|pin1|supply|vdd \$227924 i0|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30313 \$227928 \$227885 \$227927 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30314 \$227928 i0|i1|q$10 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30315 VDD|pad|pin1|supply|vdd a1|i0|q$2 \$227929 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30316 \$227929 a2|i|s|zn \$227927 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30317 VDD|pad|pin1|supply|vdd a2|i|s|zn \$227885 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30318 VDD|pad|pin1|supply|vdd \$227927 i0|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30319 \$227932 \$227886 \$227931 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30320 \$227932 i1|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30321 VDD|pad|pin1|supply|vdd i0|z$3 \$227933 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30322 \$227933 a1|a2|b|q|s \$227931 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30323 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$227886 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30324 VDD|pad|pin1|supply|vdd \$227931 d|z$84 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30325 \$227934 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30326 VDD|pad|pin1|supply|vdd \$227934 \$227887 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30327 VDD|pad|pin1|supply|vdd \$227887 \$229320 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30328 \$229320 d|z$91 \$227935 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30329 \$227935 \$227934 \$229159 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30330 \$229159 \$227936 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30331 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$229159
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30332 \$227936 \$227935 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30333 \$227936 \$227934 \$227888 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30334 \$227888 \$227887 \$229332 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30335 VDD|pad|pin1|supply|vdd \$227939 \$229332 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30336 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$227939
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30337 VDD|pad|pin1|supply|vdd \$227888 \$227939 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30338 VDD|pad|pin1|supply|vdd \$227939 R[58]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30339 VDD|pad|pin1|supply|vdd a2|zn$18 a1|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30340 a1|zn$3 a1|zn$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30341 VDD|pad|pin1|supply|vdd a2|z$12 a2|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30342 a2|zn$11 a1|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30343 a2|zn$11 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30344 VDD|pad|pin1|supply|vdd RD[39]|a2|z a1|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30345 a1|zn$4 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30346 a1|zn$4 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30347 VDD|pad|pin1|supply|vdd RD[28]|a2|z a2|zn$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30348 a2|zn$15 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30349 a2|zn$15 a2|a3|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30350 \$227944 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30351 VDD|pad|pin1|supply|vdd \$227944 \$227892 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30352 VDD|pad|pin1|supply|vdd \$227892 \$229348 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30353 \$229348 d|z$81 \$227945 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30354 \$227945 \$227944 \$229160 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30355 \$229160 \$227946 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30356 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$229160
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30357 \$227946 \$227945 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30358 \$227946 \$227944 \$227893 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30359 \$227893 \$227892 \$229352 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30360 VDD|pad|pin1|supply|vdd \$227948 \$229352 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30361 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$227948
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30362 VDD|pad|pin1|supply|vdd \$227893 \$227948 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30363 VDD|pad|pin1|supply|vdd \$227948 DUT_Header|R[3]|Vup|i|i0|q
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p
+ PS=2.67u PD=3.33u
M$30364 \$227949 a1|zn$18 \$229361 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30365 \$229361 a2|zn$19 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30366 VDD|pad|pin1|supply|vdd \$227949 i1|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30367 VDD|pad|pin1|supply|vdd RD[33]|a2|z a1|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30368 a1|zn$5 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30369 a1|zn$5 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30370 VDD|pad|pin1|supply|vdd a2|zn$22 \$227951 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30371 \$227951 a1|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30372 a2|z$11 \$227951 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30373 VDD|pad|pin1|supply|vdd a2|zn$16 \$227953 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30374 \$227953 a1|zn$8 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30375 a1|z$16 \$227953 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30376 VDD|pad|pin1|supply|vdd RD[1]|a2|z a2|zn$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30377 a2|zn$16 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30378 a2|zn$16 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30379 VDD|pad|pin1|supply|vdd RD[29]|a2|zn a2|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30380 a2|zn$17 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30381 a2|zn$17 a2|a3|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30382 VDD|pad|pin1|supply|vdd RD[36]|a2|z a3|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30383 a3|zn$4 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30384 a3|zn$4 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30385 VDD|pad|pin1|supply|vdd RD[35]|a2|z a3|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30386 a3|zn$3 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30387 a3|zn$3 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30388 \$227959 \$227899 \$227958 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30389 \$227959 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30390 VDD|pad|pin1|supply|vdd RO_control|R[1]|i|i0|nclk|q \$227960
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p
+ PS=1.93u PD=1.74u
M$30391 \$227960 s|z$1 \$227958 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30392 VDD|pad|pin1|supply|vdd s|z$1 \$227899 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30393 VDD|pad|pin1|supply|vdd \$227958 d|z$85 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30394 VDD|pad|pin1|supply|vdd a2|zn$27 \$227961 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30395 \$227961 a1|zn$23 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30396 a1|z$17 \$227961 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30397 VDD|pad|pin1|supply|vdd a2|zn$35 \$227963 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30398 \$227963 a1|zn$10 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30399 a4|z \$227963 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30400 \$227966 \$227900 \$227965 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30401 \$227966 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30402 VDD|pad|pin1|supply|vdd DUT_Header|R[11]|Vup|i|i0|q \$227967
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p
+ PS=1.93u PD=1.74u
M$30403 \$227967 s|zn$5 \$227965 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30404 VDD|pad|pin1|supply|vdd s|zn$5 \$227900 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30405 VDD|pad|pin1|supply|vdd \$227965 d|z$86 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30406 \$227968 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30407 VDD|pad|pin1|supply|vdd \$227968 \$227901 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30408 VDD|pad|pin1|supply|vdd \$227901 \$229390 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30409 \$229390 d|z$83 \$227969 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30410 \$227969 \$227968 \$229161 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30411 \$229161 \$227970 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30412 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$229161
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30413 \$227970 \$227969 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30414 \$227970 \$227968 \$227902 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30415 \$227902 \$227901 \$229395 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30416 VDD|pad|pin1|supply|vdd \$227972 \$229395 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30417 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$227972
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30418 VDD|pad|pin1|supply|vdd \$227902 \$227972 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30419 VDD|pad|pin1|supply|vdd \$227972 R[0]|clk|i|i0|n_RO_control|q
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p
+ PS=2.67u PD=3.33u
M$30420 \$227974 \$227903 \$227973 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30421 \$227974 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30422 VDD|pad|pin1|supply|vdd R[6]|i|i0|q \$227975 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30423 \$227975 s|z$1 \$227973 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30424 VDD|pad|pin1|supply|vdd s|z$1 \$227903 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30425 VDD|pad|pin1|supply|vdd \$227973 d|z$92 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30426 \$227978 \$227904 \$227977 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30427 \$227978 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30428 VDD|pad|pin1|supply|vdd R[8]|clk|i|i0|n_RO_control|q \$227979
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p
+ PS=1.93u PD=1.74u
M$30429 \$227979 s|zn$5 \$227977 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30430 VDD|pad|pin1|supply|vdd s|zn$5 \$227904 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30431 VDD|pad|pin1|supply|vdd \$227977 d|z$87 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30432 \$227981 \$227905 \$227980 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30433 \$227981 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30434 VDD|pad|pin1|supply|vdd RO_control|R[9]|i|i0|nclk|q \$227982
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p
+ PS=1.93u PD=1.74u
M$30435 \$227982 s|zn$5 \$227980 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30436 VDD|pad|pin1|supply|vdd s|zn$5 \$227905 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30437 VDD|pad|pin1|supply|vdd \$227980 d|z$93 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30438 \$227985 \$227906 \$227984 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30439 \$227985 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30440 VDD|pad|pin1|supply|vdd R[40]|i0|q \$227986 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30441 \$227986 s|zn$4 \$227984 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30442 VDD|pad|pin1|supply|vdd s|zn$4 \$227906 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30443 VDD|pad|pin1|supply|vdd \$227984 d|z$88 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30444 \$227988 \$227907 \$227987 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30445 \$227988 R[59]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30446 VDD|pad|pin1|supply|vdd i0|i1|q$1 \$227989 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30447 \$227989 s|zn$6 \$227987 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30448 VDD|pad|pin1|supply|vdd s|zn$6 \$227907 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30449 VDD|pad|pin1|supply|vdd \$227987 d|z$89 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30450 \$227991 \$227908 \$227990 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30451 \$227991 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30452 VDD|pad|pin1|supply|vdd R[45]|i0|q \$227992 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30453 \$227992 s|zn$4 \$227990 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30454 VDD|pad|pin1|supply|vdd s|zn$4 \$227908 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30455 VDD|pad|pin1|supply|vdd \$227990 d|z$94 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30456 \$227995 \$227909 \$227994 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30457 \$227995 R[57]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30458 VDD|pad|pin1|supply|vdd i0|i1|q$6 \$227996 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30459 \$227996 s|zn$6 \$227994 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30460 VDD|pad|pin1|supply|vdd s|zn$6 \$227909 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30461 VDD|pad|pin1|supply|vdd \$227994 d|z$95 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30462 DATA|core|i0|i1|p2c \$227998 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$30463 VDD|pad|pin1|supply|vdd cp|i|z$5 \$230227 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30464 VDD|pad|pin1|supply|vdd \$230227 \$230247 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30465 VDD|pad|pin1|supply|vdd \$230541 \$230249 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30466 \$230248 \$230227 \$230249 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30467 VDD|pad|pin1|supply|vdd \$230247 \$230526 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30468 \$230526 d|z$99 \$230248 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30469 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230249
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30470 \$230250 \$230247 \$230451 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30471 VDD|pad|pin1|supply|vdd \$230542 \$230451 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30472 VDD|pad|pin1|supply|vdd \$230248 \$230541 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30473 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230542
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30474 VDD|pad|pin1|supply|vdd \$230250 \$230542 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30475 \$230541 \$230227 \$230250 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30476 VDD|pad|pin1|supply|vdd \$230542 i0|i1|q$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30477 \$230252 \$230228 \$230253 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30478 \$230254 a1|a2|b|q|s \$230252 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30479 VDD|pad|pin1|supply|vdd i0|z$5 \$230254 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30480 \$230253 i1|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30481 \$230228 a1|a2|b|q|s VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30482 VDD|pad|pin1|supply|vdd \$230252 d|z$96 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30483 \$230256 \$230229 \$230257 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30484 \$230258 a2|i|s|zn \$230256 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30485 VDD|pad|pin1|supply|vdd i0|i1|q$13 \$230258 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30486 \$230257 i0|i1|q$12 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30487 \$230229 a2|i|s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30488 VDD|pad|pin1|supply|vdd \$230256 i0|z$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30489 a2|d|z a2|i|s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$30490 VDD|pad|pin1|supply|vdd cp|i|z$5 \$230230 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30491 VDD|pad|pin1|supply|vdd \$230230 \$230260 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30492 VDD|pad|pin1|supply|vdd \$230545 \$230262 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30493 \$230261 \$230230 \$230262 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30494 VDD|pad|pin1|supply|vdd \$230260 \$230529 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30495 \$230529 d|z$100 \$230261 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30496 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230262
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30497 \$230263 \$230260 \$230483 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30498 VDD|pad|pin1|supply|vdd \$230546 \$230483 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30499 VDD|pad|pin1|supply|vdd \$230261 \$230545 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30500 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230546
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30501 VDD|pad|pin1|supply|vdd \$230263 \$230546 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30502 \$230545 \$230230 \$230263 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30503 VDD|pad|pin1|supply|vdd \$230546 a1|i0|q$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30504 VDD|pad|pin1|supply|vdd cp|i|z$5 \$230231 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30505 VDD|pad|pin1|supply|vdd \$230231 \$230264 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30506 VDD|pad|pin1|supply|vdd \$230547 \$230266 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30507 \$230265 \$230231 \$230266 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30508 VDD|pad|pin1|supply|vdd \$230264 \$230530 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30509 \$230530 d|z$101 \$230265 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30510 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230266
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30511 \$230267 \$230264 \$230486 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30512 VDD|pad|pin1|supply|vdd \$230548 \$230486 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30513 VDD|pad|pin1|supply|vdd \$230265 \$230547 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30514 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230548
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30515 VDD|pad|pin1|supply|vdd \$230267 \$230548 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30516 \$230547 \$230231 \$230267 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30517 VDD|pad|pin1|supply|vdd \$230548 R[61]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30518 \$230269 a1|zn$3 \$230531 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30519 VDD|pad|pin1|supply|vdd a2|zn$20 \$230531 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30520 VDD|pad|pin1|supply|vdd \$230269 i1|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30521 \$230270 \$230232 \$230271 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30522 \$230272 s|zn$6 \$230270 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30523 VDD|pad|pin1|supply|vdd i0|i1|q$2 \$230272 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30524 \$230271 R[58]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30525 \$230232 s|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30526 VDD|pad|pin1|supply|vdd \$230270 d|z$91 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30527 VDD|pad|pin1|supply|vdd RD[4]|a2|z a1|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30528 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30529 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a1|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30530 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a4|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30531 VDD|pad|pin1|supply|vdd a2|z$12 a4|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30532 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a4|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30533 VDD|pad|pin1|supply|vdd RD[43]|a4|z a4|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30534 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30535 VDD|pad|pin1|supply|vdd a2|z$12 a1|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30536 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a1|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30537 VDD|pad|pin1|supply|vdd RD[12]|a4|zn a1|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30538 VDD|pad|pin1|supply|vdd a3|zn$4 a2|zn$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30539 VDD|pad|pin1|supply|vdd a2|zn$15 a2|zn$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30540 VDD|pad|pin1|supply|vdd a1|zn$6 a2|zn$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30541 VDD|pad|pin1|supply|vdd a4|zn$5 a2|zn$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30542 \$230277 \$230233 \$230278 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30543 \$230279 s|zn$4 \$230277 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30544 VDD|pad|pin1|supply|vdd R[43]|i0|q \$230279 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30545 \$230278 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30546 \$230233 s|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30547 VDD|pad|pin1|supply|vdd \$230277 d|z$78 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30548 VDD|pad|pin1|supply|vdd RD[25]|a2|zn a4|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30549 VDD|pad|pin1|supply|vdd a1|a3|z a4|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30550 VDD|pad|pin1|supply|vdd a2|a3|z$1 a4|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30551 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30552 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a2|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30553 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30554 VDD|pad|pin1|supply|vdd RD[19]|a4|z a2|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30555 VDD|pad|pin1|supply|vdd a3|zn$5 i1|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30556 VDD|pad|pin1|supply|vdd a2|z$11 i1|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30557 VDD|pad|pin1|supply|vdd a1|z$16 i1|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30558 VDD|pad|pin1|supply|vdd a4|zn$4 i1|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30559 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30560 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a1|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30561 VDD|pad|pin1|supply|vdd a1|z$15 a1|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30562 VDD|pad|pin1|supply|vdd RD[17]|a4|z a1|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30563 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30564 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a1|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30565 VDD|pad|pin1|supply|vdd a1|z$15 a1|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30566 VDD|pad|pin1|supply|vdd RD[23]|a4|z a1|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30567 VDD|pad|pin1|supply|vdd a2|zn$25 \$230285 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30568 VDD|pad|pin1|supply|vdd a1|zn$13 \$230285 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30569 VDD|pad|pin1|supply|vdd \$230285 a4|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30570 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a3|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30571 VDD|pad|pin1|supply|vdd a2|z$12 a3|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30572 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a3|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30573 VDD|pad|pin1|supply|vdd RD[41]|a4|z a3|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30574 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30575 VDD|pad|pin1|supply|vdd a2|z$12 a2|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30576 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30577 VDD|pad|pin1|supply|vdd RD[9]|a4|z a2|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30578 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a2|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30579 VDD|pad|pin1|supply|vdd a2|z$12 a2|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30580 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30581 VDD|pad|pin1|supply|vdd RD[46]|a4|z a2|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30582 VDD|pad|pin1|supply|vdd RD[38]|a2|z a1|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30583 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a1|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30584 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a1|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30585 VDD|pad|pin1|supply|vdd RD[7]|a2|zn a2|zn$24 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30586 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$24 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30587 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a2|zn$24 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30588 z$34 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$30589 VDD|pad|pin1|supply|vdd i|z$115 \$230293 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$30590 VDD|pad|pin1|supply|vdd \$230293 cp|i|z$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$30591 VDD|pad|pin1|supply|vdd cp|i|z$7 \$230234 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30592 VDD|pad|pin1|supply|vdd \$230234 \$230294 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30593 VDD|pad|pin1|supply|vdd \$230551 \$230296 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30594 \$230295 \$230234 \$230296 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30595 VDD|pad|pin1|supply|vdd \$230294 \$230540 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30596 \$230540 d|z$102 \$230295 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30597 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230296
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30598 \$230297 \$230294 \$230495 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30599 VDD|pad|pin1|supply|vdd \$230552 \$230495 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30600 VDD|pad|pin1|supply|vdd \$230295 \$230551 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30601 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230552
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30602 VDD|pad|pin1|supply|vdd \$230297 \$230552 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30603 \$230551 \$230234 \$230297 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30604 VDD|pad|pin1|supply|vdd \$230552 DUT_Footer|R[2]|Vdn|i|i0|q
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p
+ PS=2.67u PD=3.33u
M$30605 VDD|pad|pin1|supply|vdd cp|i|z$7 \$230235 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30606 VDD|pad|pin1|supply|vdd \$230235 \$230299 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30607 VDD|pad|pin1|supply|vdd \$230553 \$230301 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30608 \$230300 \$230235 \$230301 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30609 VDD|pad|pin1|supply|vdd \$230299 \$230539 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30610 \$230539 d|z$103 \$230300 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30611 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230301
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30612 \$230302 \$230299 \$230494 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30613 VDD|pad|pin1|supply|vdd \$230554 \$230494 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30614 VDD|pad|pin1|supply|vdd \$230300 \$230553 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30615 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230554
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30616 VDD|pad|pin1|supply|vdd \$230302 \$230554 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30617 \$230553 \$230235 \$230302 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30618 VDD|pad|pin1|supply|vdd \$230554 R[41]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30619 \$230304 \$230236 \$230305 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30620 \$230306 s|zn$6 \$230304 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30621 VDD|pad|pin1|supply|vdd i0|i1|q \$230306 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30622 \$230305 R[56]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30623 \$230236 s|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30624 VDD|pad|pin1|supply|vdd \$230304 d|z$97 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30625 VDD|pad|pin1|supply|vdd cp|z$4 \$230237 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30626 VDD|pad|pin1|supply|vdd \$230237 \$230308 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30627 VDD|pad|pin1|supply|vdd \$230555 \$230310 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30628 \$230309 \$230237 \$230310 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30629 VDD|pad|pin1|supply|vdd \$230308 \$230538 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30630 \$230538 d|z$97 \$230309 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30631 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230310
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30632 \$230311 \$230308 \$230488 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30633 VDD|pad|pin1|supply|vdd \$230556 \$230488 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30634 VDD|pad|pin1|supply|vdd \$230309 \$230555 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30635 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230556
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30636 VDD|pad|pin1|supply|vdd \$230311 \$230556 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30637 \$230555 \$230237 \$230311 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30638 VDD|pad|pin1|supply|vdd \$230556 R[56]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30639 \$230312 \$230238 \$230313 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30640 \$230314 s|zn$6 \$230312 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30641 VDD|pad|pin1|supply|vdd i0|i1|q$3 \$230314 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30642 \$230313 R[62]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30643 \$230238 s|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30644 VDD|pad|pin1|supply|vdd \$230312 d|z$98 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30645 \$232162 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30646 VDD|pad|pin1|supply|vdd \$232162 \$232070 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30647 VDD|pad|pin1|supply|vdd \$232070 \$233354 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30648 \$233354 d|z$104 \$232163 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30649 \$232163 \$232162 \$233239 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30650 \$233239 \$232164 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30651 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$233239
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30652 \$232164 \$232163 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30653 \$232164 \$232162 \$232071 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30654 \$232071 \$232070 \$233364 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30655 VDD|pad|pin1|supply|vdd \$232166 \$233364 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30656 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232166
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30657 VDD|pad|pin1|supply|vdd \$232071 \$232166 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30658 VDD|pad|pin1|supply|vdd \$232166 i0|i1|q$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30659 \$232167 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30660 VDD|pad|pin1|supply|vdd \$232167 \$232072 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30661 VDD|pad|pin1|supply|vdd \$232072 \$233370 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30662 \$233370 d|z$96 \$232168 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30663 \$232168 \$232167 \$233240 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30664 \$233240 \$232169 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30665 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$233240
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30666 \$232169 \$232168 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30667 \$232169 \$232167 \$232073 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30668 \$232073 \$232072 \$233366 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30669 VDD|pad|pin1|supply|vdd \$232171 \$233366 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30670 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232171
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30671 VDD|pad|pin1|supply|vdd \$232073 \$232171 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30672 VDD|pad|pin1|supply|vdd \$232171 a1|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30673 \$232173 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30674 VDD|pad|pin1|supply|vdd \$232173 \$232075 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30675 VDD|pad|pin1|supply|vdd \$232075 \$233373 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30676 \$233373 d|z$105 \$232174 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30677 \$232174 \$232173 \$233241 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30678 \$233241 \$232175 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30679 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$233241
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30680 \$232175 \$232174 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30681 \$232175 \$232173 \$232076 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30682 \$232076 \$232075 \$233380 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30683 VDD|pad|pin1|supply|vdd \$232177 \$233380 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30684 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232177
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30685 VDD|pad|pin1|supply|vdd \$232076 \$232177 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30686 VDD|pad|pin1|supply|vdd \$232177 DOUT_DAT|c2p|core|i|q
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p
+ PS=2.67u PD=3.33u
M$30687 \$233242 a1|zn$12 \$232178 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30688 \$232178 b|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30689 VDD|pad|pin1|supply|vdd \$232178 d|z$100 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30690 \$233242 a2|zn$29 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30691 \$232179 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30692 VDD|pad|pin1|supply|vdd \$232179 \$232078 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30693 VDD|pad|pin1|supply|vdd \$232078 \$233383 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30694 \$233383 d|z$106 \$232180 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30695 \$232180 \$232179 \$233243 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30696 \$233243 \$232181 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30697 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$233243
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30698 \$232181 \$232180 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30699 \$232181 \$232179 \$232079 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30700 \$232079 \$232078 \$233388 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30701 VDD|pad|pin1|supply|vdd \$232183 \$233388 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30702 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232183
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30703 VDD|pad|pin1|supply|vdd \$232079 \$232183 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30704 VDD|pad|pin1|supply|vdd \$232183 R[5]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30705 \$232186 \$232080 \$232185 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30706 \$232186 R[61]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30707 VDD|pad|pin1|supply|vdd i0|i1|q$7 \$232187 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30708 \$232187 s|zn$6 \$232185 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30709 VDD|pad|pin1|supply|vdd s|zn$6 \$232080 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30710 VDD|pad|pin1|supply|vdd \$232185 d|z$101 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30711 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a3|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30712 a3|zn$6 a2|z$12 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30713 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a3|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30714 a3|zn$6 RD[40]|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30715 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$18 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30716 a2|zn$18 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30717 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$18 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30718 a2|zn$18 RD[20]|a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30719 VDD|pad|pin1|supply|vdd a1|a3|z a3|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30720 a3|zn$7 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30721 VDD|pad|pin1|supply|vdd a1|z$15 a3|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30722 a3|zn$7 RD[16]|a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30723 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a4|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30724 a4|zn$5 a2|z$12 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30725 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a4|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30726 a4|zn$5 RD[44]|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30727 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$26 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30728 a2|zn$26 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30729 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$26 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30730 a2|zn$26 RD[18]|a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30731 VDD|pad|pin1|supply|vdd a3|zn$7 a1|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30732 a1|zn$12 a2|zn$28 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30733 VDD|pad|pin1|supply|vdd a1|zn$17 a1|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30734 a1|zn$12 a4|zn$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30735 VDD|pad|pin1|supply|vdd RD[0]|a2|z a2|zn$28 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30736 a2|zn$28 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30737 a2|zn$28 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30738 VDD|pad|pin1|supply|vdd a3|zn$3 a2|zn$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30739 a2|zn$19 a2|zn$21 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30740 VDD|pad|pin1|supply|vdd a1|zn$21 a2|zn$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30741 a2|zn$19 a4|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30742 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$27 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30743 a2|zn$27 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30744 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$27 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30745 a2|zn$27 RD[22]|a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30746 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30747 a1|zn$11 a2|z$12 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30748 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a1|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30749 a1|zn$11 RD[13]|a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30750 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30751 a1|zn$13 a2|z$12 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30752 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a1|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30753 a1|zn$13 RD[15]|a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30754 VDD|pad|pin1|supply|vdd a3|zn$10 a2|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30755 a2|zn$14 a2|zn$34 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30756 VDD|pad|pin1|supply|vdd a1|zn$22 a2|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30757 a2|zn$14 a4|zn$8 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30758 VDD|pad|pin1|supply|vdd a3|zn$11 i1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30759 i1|zn$1 a2|z$13 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30760 VDD|pad|pin1|supply|vdd a1|zn$4 i1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30761 i1|zn$1 a4|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30762 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a4|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30763 a4|zn$6 a2|z$12 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30764 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a4|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30765 a4|zn$6 RD[42]|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30766 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a4|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30767 a4|zn$8 a2|z$12 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30768 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a4|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30769 a4|zn$8 RD[45]|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30770 VDD|pad|pin1|supply|vdd a3|zn$8 i1|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30771 i1|zn$2 a2|zn$23 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30772 VDD|pad|pin1|supply|vdd a1|z$17 i1|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30773 i1|zn$2 a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30774 VDD|pad|pin1|supply|vdd RD[30]|a2|z a3|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30775 a3|zn$8 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30776 a3|zn$8 a2|a3|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30777 \$232197 \$232099 \$232196 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$30778 \$232197 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30779 VDD|pad|pin1|supply|vdd DUT_Footer|R[2]|Vdn|i|i0|q \$232198
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p
+ PS=1.93u PD=1.74u
M$30780 \$232198 s|z$1 \$232196 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30781 VDD|pad|pin1|supply|vdd s|z$1 \$232099 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$30782 VDD|pad|pin1|supply|vdd \$232196 d|z$102 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30783 \$232199 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30784 VDD|pad|pin1|supply|vdd \$232199 \$232100 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30785 VDD|pad|pin1|supply|vdd \$232100 \$233596 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30786 \$233596 d|z$107 \$232200 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30787 \$232200 \$232199 \$233244 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30788 \$233244 \$232201 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30789 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$233244
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30790 \$232201 \$232200 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30791 \$232201 \$232199 \$232101 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30792 \$232101 \$232100 \$233604 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30793 VDD|pad|pin1|supply|vdd \$232203 \$233604 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30794 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232203
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30795 VDD|pad|pin1|supply|vdd \$232101 \$232203 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30796 VDD|pad|pin1|supply|vdd \$232203 R[13]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30797 \$232205 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30798 VDD|pad|pin1|supply|vdd \$232205 \$232102 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30799 VDD|pad|pin1|supply|vdd \$232102 \$233611 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30800 \$233611 d|z$93 \$232206 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30801 \$232206 \$232205 \$233245 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30802 \$233245 \$232207 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30803 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$233245
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30804 \$232207 \$232206 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30805 \$232207 \$232205 \$232103 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30806 \$232103 \$232102 \$233625 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30807 VDD|pad|pin1|supply|vdd \$232209 \$233625 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30808 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232209
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30809 VDD|pad|pin1|supply|vdd \$232103 \$232209 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30810 VDD|pad|pin1|supply|vdd \$232209 RO_control|R[9]|i|i0|nclk|q
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p
+ PS=2.67u PD=3.33u
M$30811 \$232210 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30812 VDD|pad|pin1|supply|vdd \$232210 \$232104 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30813 VDD|pad|pin1|supply|vdd \$232104 \$233618 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30814 \$233618 d|z$108 \$232211 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30815 \$232211 \$232210 \$233246 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30816 \$233246 \$232212 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30817 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$233246
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30818 \$232212 \$232211 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30819 \$232212 \$232210 \$232105 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30820 \$232105 \$232104 \$233632 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30821 VDD|pad|pin1|supply|vdd \$232214 \$233632 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30822 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232214
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30823 VDD|pad|pin1|supply|vdd \$232105 \$232214 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30824 VDD|pad|pin1|supply|vdd \$232214 R[42]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30825 \$232216 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30826 VDD|pad|pin1|supply|vdd \$232216 \$232106 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30827 VDD|pad|pin1|supply|vdd \$232106 \$233643 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30828 \$233643 d|z$95 \$232217 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30829 \$232217 \$232216 \$233247 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30830 \$233247 \$232218 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30831 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$233247
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30832 \$232218 \$232217 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30833 \$232218 \$232216 \$232107 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30834 \$232107 \$232106 \$233637 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30835 VDD|pad|pin1|supply|vdd \$232220 \$233637 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30836 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232220
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30837 VDD|pad|pin1|supply|vdd \$232107 \$232220 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30838 VDD|pad|pin1|supply|vdd \$232220 R[57]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30839 \$234140 \$233988 \$234141 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30840 \$234142 a1|a2|b|q|s \$234140 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30841 VDD|pad|pin1|supply|vdd i0|z$6 \$234142 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30842 \$234141 i1|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30843 \$233988 a1|a2|b|q|s VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30844 VDD|pad|pin1|supply|vdd \$234140 d|z$104 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30845 \$234143 \$233989 \$234144 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30846 \$234145 a2|i|s|zn \$234143 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30847 VDD|pad|pin1|supply|vdd i0|i1|q$11 \$234145 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30848 \$234144 i0|i1|q$13 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30849 \$233989 a2|i|s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30850 VDD|pad|pin1|supply|vdd \$234143 i0|z$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30851 \$234146 \$233990 \$234147 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30852 \$234148 a2|i|s|zn \$234146 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30853 VDD|pad|pin1|supply|vdd i0|i1|q$12 \$234148 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30854 \$234147 a1|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30855 \$233990 a2|i|s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30856 VDD|pad|pin1|supply|vdd \$234146 i0|z$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30857 \$234149 \$233991 \$234150 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30858 \$234151 a1|a2|b|q|s \$234149 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30859 VDD|pad|pin1|supply|vdd i0|z$4 \$234151 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30860 \$234150 i1|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30861 \$233991 a1|a2|b|q|s VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30862 VDD|pad|pin1|supply|vdd \$234149 d|z$99 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30863 VDD|pad|pin1|supply|vdd a2|d|z \$234152 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30864 VDD|pad|pin1|supply|vdd a1|i1|q \$234152 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30865 VDD|pad|pin1|supply|vdd \$234152 d|z$105 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30866 \$234153 a1|i0|q$2 \$234415 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30867 \$234415 a2|i|s|zn \$234153 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.4565p AD=0.4565p PS=1.93u PD=1.93u
M$30868 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$234153 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30869 VDD|pad|pin1|supply|vdd \$234415 b|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30870 VDD|pad|pin1|supply|vdd a2|zn$30 a2|zn$29 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30871 VDD|pad|pin1|supply|vdd a1|a2|b|q|s a2|zn$29 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30872 VDD|pad|pin1|supply|vdd a3|zn$6 a2|zn$29 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30873 \$234156 \$233992 \$234157 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30874 \$234158 s|z$1 \$234156 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30875 VDD|pad|pin1|supply|vdd R[5]|i|i0|q \$234158 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30876 \$234157 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30877 \$233992 s|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30878 VDD|pad|pin1|supply|vdd \$234156 d|z$106 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30879 VDD|pad|pin1|supply|vdd a2|zn$31 a1|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30880 VDD|pad|pin1|supply|vdd a1|zn$15 a1|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30881 VDD|pad|pin1|supply|vdd RD[32]|a2|z a2|zn$30 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30882 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a2|zn$30 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30883 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a2|zn$30 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30884 VDD|pad|pin1|supply|vdd RD[34]|a2|z a1|zn$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30885 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a1|zn$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30886 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a1|zn$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30887 VDD|pad|pin1|supply|vdd RD[2]|a2|z a3|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30888 VDD|pad|pin1|supply|vdd a1|a3|z a3|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30889 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a3|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30890 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$31 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30891 VDD|pad|pin1|supply|vdd a2|z$12 a2|zn$31 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30892 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$31 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30893 VDD|pad|pin1|supply|vdd RD[10]|a4|zn a2|zn$31 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30894 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30895 VDD|pad|pin1|supply|vdd a2|z$12 a1|zn$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30896 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a1|zn$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30897 VDD|pad|pin1|supply|vdd RD[11]|a4|zn a1|zn$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30898 VDD|pad|pin1|supply|vdd a3|zn$9 a2|zn$32 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30899 VDD|pad|pin1|supply|vdd a2|zn$26 a2|zn$32 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30900 VDD|pad|pin1|supply|vdd a1|zn$19 a2|zn$32 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30901 VDD|pad|pin1|supply|vdd a4|zn$6 a2|zn$32 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30902 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30903 VDD|pad|pin1|supply|vdd a2|z$12 a1|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30904 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a1|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30905 VDD|pad|pin1|supply|vdd RD[8]|a4|z a1|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30906 VDD|pad|pin1|supply|vdd a2|zn$33 a1|zn$18 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30907 VDD|pad|pin1|supply|vdd a1|zn$16 a1|zn$18 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30908 VDD|pad|pin1|supply|vdd RD[24]|a2|z a4|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30909 VDD|pad|pin1|supply|vdd a1|a3|z a4|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30910 VDD|pad|pin1|supply|vdd a2|a3|z$1 a4|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30911 VDD|pad|pin1|supply|vdd RD[26]|a2|z a1|zn$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30912 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30913 VDD|pad|pin1|supply|vdd a2|a3|z$1 a1|zn$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30914 VDD|pad|pin1|supply|vdd RD[37]|a2|z a3|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30915 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a3|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30916 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a3|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30917 VDD|pad|pin1|supply|vdd RD[27]|a2|zn a2|zn$33 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30918 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$33 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30919 VDD|pad|pin1|supply|vdd a2|a3|z$1 a2|zn$33 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30920 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$34 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30921 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a2|zn$34 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30922 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$34 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30923 VDD|pad|pin1|supply|vdd RD[21]|a4|z a2|zn$34 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30924 VDD|pad|pin1|supply|vdd RD[31]|a2|zn a3|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30925 VDD|pad|pin1|supply|vdd a1|a3|z a3|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30926 VDD|pad|pin1|supply|vdd a2|a3|z$1 a3|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30927 VDD|pad|pin1|supply|vdd a2|zn$24 \$234173 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30928 VDD|pad|pin1|supply|vdd a1|zn$9 \$234173 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30929 VDD|pad|pin1|supply|vdd \$234173 a2|z$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30930 VDD|pad|pin1|supply|vdd a2|zn$17 a1|zn$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30931 VDD|pad|pin1|supply|vdd a1|zn$11 a1|zn$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30932 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a2|zn$25 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30933 VDD|pad|pin1|supply|vdd a2|z$12 a2|zn$25 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30934 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$25 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30935 VDD|pad|pin1|supply|vdd RD[47]|a4|z a2|zn$25 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30936 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$35 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30937 VDD|pad|pin1|supply|vdd a2|z$12 a2|zn$35 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$30938 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$35 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30939 VDD|pad|pin1|supply|vdd RD[14]|a4|zn a2|zn$35 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30940 VDD|pad|pin1|supply|vdd RD[3]|a2|z a1|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30941 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30942 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a1|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30943 VDD|pad|pin1|supply|vdd RD[5]|a2|zn a1|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30944 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30945 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a1|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30946 VDD|pad|pin1|supply|vdd RD[6]|a2|zn a1|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30947 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30948 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a1|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30949 \$234179 \$233993 \$234180 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30950 \$234181 s|zn$5 \$234179 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30951 VDD|pad|pin1|supply|vdd R[13]|i|i0|q \$234181 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30952 \$234180 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30953 \$233993 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30954 VDD|pad|pin1|supply|vdd \$234179 d|z$107 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30955 VDD|pad|pin1|supply|vdd cp|i|z$7 \$234182 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30956 VDD|pad|pin1|supply|vdd \$234182 \$234183 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30957 VDD|pad|pin1|supply|vdd \$234416 \$234185 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30958 \$234184 \$234182 \$234185 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30959 VDD|pad|pin1|supply|vdd \$234183 \$234398 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30960 \$234398 d|z$92 \$234184 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30961 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$234185
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30962 \$234186 \$234183 \$234368 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30963 VDD|pad|pin1|supply|vdd \$234417 \$234368 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30964 VDD|pad|pin1|supply|vdd \$234184 \$234416 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30965 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$234417
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30966 VDD|pad|pin1|supply|vdd \$234186 \$234417 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30967 \$234416 \$234182 \$234186 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30968 VDD|pad|pin1|supply|vdd \$234417 R[6]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30969 \$234187 \$233994 \$234188 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30970 \$234189 s|zn$4 \$234187 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30971 VDD|pad|pin1|supply|vdd R[41]|i0|q \$234189 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30972 \$234188 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30973 \$233994 s|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30974 VDD|pad|pin1|supply|vdd \$234187 d|z$103 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30975 \$234190 \$233995 \$234191 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$30976 \$234192 s|zn$4 \$234190 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$30977 VDD|pad|pin1|supply|vdd R[42]|i0|q \$234192 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$30978 \$234191 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$30979 \$233995 s|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$30980 VDD|pad|pin1|supply|vdd \$234190 d|z$108 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$30981 VDD|pad|pin1|supply|vdd cp|z$4 \$234193 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30982 VDD|pad|pin1|supply|vdd \$234193 \$234194 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30983 VDD|pad|pin1|supply|vdd \$234418 \$234196 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30984 \$234195 \$234193 \$234196 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30985 VDD|pad|pin1|supply|vdd \$234194 \$234411 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30986 \$234411 d|z$94 \$234195 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30987 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$234196
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30988 \$234197 \$234194 \$234360 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30989 VDD|pad|pin1|supply|vdd \$234419 \$234360 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30990 VDD|pad|pin1|supply|vdd \$234195 \$234418 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30991 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$234419
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30992 VDD|pad|pin1|supply|vdd \$234197 \$234419 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30993 \$234418 \$234193 \$234197 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30994 VDD|pad|pin1|supply|vdd \$234419 R[45]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30995 VDD|pad|pin1|supply|vdd cp|z$4 \$234198 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30996 VDD|pad|pin1|supply|vdd \$234198 \$234199 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30997 VDD|pad|pin1|supply|vdd \$234420 \$234201 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30998 \$234200 \$234198 \$234201 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30999 VDD|pad|pin1|supply|vdd \$234199 \$234413 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$31000 \$234413 d|z$98 \$234200 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$31001 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$234201
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$31002 \$234202 \$234199 \$234357 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$31003 VDD|pad|pin1|supply|vdd \$234421 \$234357 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$31004 VDD|pad|pin1|supply|vdd \$234200 \$234420 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$31005 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$234421
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$31006 VDD|pad|pin1|supply|vdd \$234202 \$234421 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$31007 \$234420 \$234198 \$234202 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$31008 VDD|pad|pin1|supply|vdd \$234421 R[62]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$31009 \$236468 \$235938 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3864p
+ AD=0.41165p PS=2.93u PD=2.12u
M$31010 RO2VDD|VDD|anode|cathode|nclk|pad IN|Vout \$235938
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.41165p
+ AD=0.4088p PS=2.12u PD=2.97u
M$31011 \$235941 \$235940 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3864p
+ AD=0.2128p PS=2.93u PD=1.5u
M$31012 RO2VDD|VDD|anode|cathode|nclk|pad \$235941 Q
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p
+ AD=0.3808p PS=1.5u PD=2.92u
M$31013 \$236469 \$235946 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3864p
+ AD=0.41165p PS=2.93u PD=2.12u
M$31014 RO2VDD|VDD|anode|cathode|nclk|pad Q \$235946
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.41165p
+ AD=0.4088p PS=2.12u PD=2.97u
M$31015 \$235949 \$235948 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3864p
+ AD=0.2128p PS=2.93u PD=1.5u
M$31016 RO2VDD|VDD|anode|cathode|nclk|pad \$235949 Q$1
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p
+ AD=0.3808p PS=1.5u PD=2.92u
M$31017 \$236470 \$235954 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3864p
+ AD=0.41165p PS=2.93u PD=2.12u
M$31018 RO2VDD|VDD|anode|cathode|nclk|pad Q$1 \$235954
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.41165p
+ AD=0.4088p PS=2.12u PD=2.97u
M$31019 \$235957 \$235956 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3864p
+ AD=0.2128p PS=2.93u PD=1.5u
M$31020 RO2VDD|VDD|anode|cathode|nclk|pad \$235957 Q$2
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p
+ AD=0.3808p PS=1.5u PD=2.92u
M$31021 \$236471 \$235962 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3864p
+ AD=0.41165p PS=2.93u PD=2.12u
M$31022 RO2VDD|VDD|anode|cathode|nclk|pad Q$2 \$235962
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.41165p
+ AD=0.4088p PS=2.12u PD=2.97u
M$31023 \$235965 \$235964 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3864p
+ AD=0.2128p PS=2.93u PD=1.5u
M$31024 RO2VDD|VDD|anode|cathode|nclk|pad \$235965 Q$3
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p
+ AD=0.3808p PS=1.5u PD=2.92u
M$31025 \$236472 \$235970 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3864p
+ AD=0.41165p PS=2.93u PD=2.12u
M$31026 RO2VDD|VDD|anode|cathode|nclk|pad Q$3 \$235970
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.41165p
+ AD=0.4088p PS=2.12u PD=2.97u
M$31027 \$235973 \$235972 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3864p
+ AD=0.2128p PS=2.93u PD=1.5u
M$31028 RO2VDD|VDD|anode|cathode|nclk|pad \$235973 OUT|Q|c2p|core|i
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p
+ AD=0.3808p PS=1.5u PD=2.92u
M$31029 RO2VDD|VDD|anode|cathode|nclk|pad D|Q_N \$235935
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$31030 RO2VDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$235935
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.3623875p
+ AD=0.0798p PS=2.605u PD=0.8u
M$31031 RO2VDD|VDD|anode|cathode|nclk|pad \$236455 \$235757
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1u AS=0.3623875p
+ AD=0.34p PS=2.605u PD=2.68u
M$31032 \$235940 \$236468 \$236517 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.2048p AD=0.09345p PS=1.63u PD=0.865u
M$31033 \$236517 \$236456 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.09345p
+ AD=0.204p PS=0.865u PD=1.835u
M$31034 RO2VDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$236456
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.204p
+ AD=0.0798p PS=1.835u PD=0.8u
M$31035 RO2VDD|VDD|anode|cathode|nclk|pad \$235940 \$236456
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.2639p
+ AD=0.0798p PS=1.81u PD=0.8u
M$31036 \$235757 \$235938 \$235940 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.2048p PS=2.68u PD=1.63u
M$31037 RO2VDD|VDD|anode|cathode|nclk|pad \$235940 D|Q_N
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2639p
+ AD=0.4312p PS=1.81u PD=3.01u
M$31038 RO2VDD|VDD|anode|cathode|nclk|pad D|Q_N$1 \$235943
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$31039 RO2VDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$235943
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.3623875p
+ AD=0.0798p PS=2.605u PD=0.8u
M$31040 RO2VDD|VDD|anode|cathode|nclk|pad \$236457 \$235758
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1u AS=0.3623875p
+ AD=0.34p PS=2.605u PD=2.68u
M$31041 \$235948 \$236469 \$236515 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.2048p AD=0.09345p PS=1.63u PD=0.865u
M$31042 \$236515 \$236458 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.09345p
+ AD=0.204p PS=0.865u PD=1.835u
M$31043 RO2VDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$236458
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.204p
+ AD=0.0798p PS=1.835u PD=0.8u
M$31044 RO2VDD|VDD|anode|cathode|nclk|pad \$235948 \$236458
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.2639p
+ AD=0.0798p PS=1.81u PD=0.8u
M$31045 \$235758 \$235946 \$235948 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.2048p PS=2.68u PD=1.63u
M$31046 RO2VDD|VDD|anode|cathode|nclk|pad \$235948 D|Q_N$1
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2639p
+ AD=0.4312p PS=1.81u PD=3.01u
M$31047 RO2VDD|VDD|anode|cathode|nclk|pad D|Q_N$2 \$235951
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$31048 RO2VDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$235951
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.3623875p
+ AD=0.0798p PS=2.605u PD=0.8u
M$31049 RO2VDD|VDD|anode|cathode|nclk|pad \$236459 \$235759
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1u AS=0.3623875p
+ AD=0.34p PS=2.605u PD=2.68u
M$31050 \$235956 \$236470 \$236513 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.2048p AD=0.09345p PS=1.63u PD=0.865u
M$31051 \$236513 \$236460 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.09345p
+ AD=0.204p PS=0.865u PD=1.835u
M$31052 RO2VDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$236460
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.204p
+ AD=0.0798p PS=1.835u PD=0.8u
M$31053 RO2VDD|VDD|anode|cathode|nclk|pad \$235956 \$236460
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.2639p
+ AD=0.0798p PS=1.81u PD=0.8u
M$31054 \$235759 \$235954 \$235956 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.2048p PS=2.68u PD=1.63u
M$31055 RO2VDD|VDD|anode|cathode|nclk|pad \$235956 D|Q_N$2
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2639p
+ AD=0.4312p PS=1.81u PD=3.01u
M$31056 RO2VDD|VDD|anode|cathode|nclk|pad D|Q_N$3 \$235959
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$31057 RO2VDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$235959
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.3623875p
+ AD=0.0798p PS=2.605u PD=0.8u
M$31058 RO2VDD|VDD|anode|cathode|nclk|pad \$236461 \$235760
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1u AS=0.3623875p
+ AD=0.34p PS=2.605u PD=2.68u
M$31059 \$235964 \$236471 \$236511 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.2048p AD=0.09345p PS=1.63u PD=0.865u
M$31060 \$236511 \$236462 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.09345p
+ AD=0.204p PS=0.865u PD=1.835u
M$31061 RO2VDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$236462
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.204p
+ AD=0.0798p PS=1.835u PD=0.8u
M$31062 RO2VDD|VDD|anode|cathode|nclk|pad \$235964 \$236462
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.2639p
+ AD=0.0798p PS=1.81u PD=0.8u
M$31063 \$235760 \$235962 \$235964 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.2048p PS=2.68u PD=1.63u
M$31064 RO2VDD|VDD|anode|cathode|nclk|pad \$235964 D|Q_N$3
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2639p
+ AD=0.4312p PS=1.81u PD=3.01u
M$31065 RO2VDD|VDD|anode|cathode|nclk|pad D|Q_N$4 \$235967
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$31066 RO2VDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$235967
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.3623875p
+ AD=0.0798p PS=2.605u PD=0.8u
M$31067 RO2VDD|VDD|anode|cathode|nclk|pad \$236463 \$235761
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1u AS=0.3623875p
+ AD=0.34p PS=2.605u PD=2.68u
M$31068 \$235972 \$236472 \$236509 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.2048p AD=0.09345p PS=1.63u PD=0.865u
M$31069 \$236509 \$236464 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.09345p
+ AD=0.204p PS=0.865u PD=1.835u
M$31070 RO2VDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$236464
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.204p
+ AD=0.0798p PS=1.835u PD=0.8u
M$31071 RO2VDD|VDD|anode|cathode|nclk|pad \$235972 \$236464
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.2639p
+ AD=0.0798p PS=1.81u PD=0.8u
M$31072 \$235761 \$235970 \$235972 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.2048p PS=2.68u PD=1.63u
M$31073 RO2VDD|VDD|anode|cathode|nclk|pad \$235972 D|Q_N$4
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2639p
+ AD=0.4312p PS=1.81u PD=3.01u
M$31074 \$236475 R[8]|clk|i|i0|n_RO_control|q RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=40.8u AS=13.872p
+ AD=13.872p PS=89.76u PD=89.76u
M$31086 \$236475 Vin|Vout Vin RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos
+ L=0.45u W=13.6u AS=4.624p AD=4.624p PS=29.92u PD=29.92u
M$31090 Vin RO_control|R[9]|i|i0|nclk|q \$235205
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31091 Vin RO_control|R[9]|i|i0|nclk|q DUT_gate|core|p2c$1
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31092 \$236476 DUT_Header|R[11]|Vup|i|i0|q RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=40.8u AS=13.872p
+ AD=13.872p PS=89.76u PD=89.76u
M$31104 \$236476 Vin Vin|Vout|core|extra_load|padres
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31108 Vin|Vout|core|extra_load|padres RO_control|R[9]|i|i0|nclk|q
+ Drain_Sense|Vout|core|padres RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos
+ L=0.45u W=3.4u AS=1.156p AD=1.156p PS=7.48u PD=7.48u
M$31109 Vin|Vout|core|extra_load|padres RO_control|R[9]|i|i0|nclk|q
+ Drain_Force|Vout|core|padres RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos
+ L=0.45u W=13.6u AS=4.624p AD=4.624p PS=29.92u PD=29.92u
M$31113 RO2VDD|VDD|anode|cathode|nclk|pad R[8]|clk|i|i0|n_RO_control|q \$236477
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=40.8u AS=13.872p
+ AD=13.872p PS=89.76u PD=89.76u
M$31125 \$236477 Vin|Vout|core|extra_load|padres Vout
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31129 \$235211 RO2VDD|VDD|anode|cathode|nclk|pad Vout
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31130 VSS|anode|cathode|clk|vss RO2VDD|VDD|anode|cathode|nclk|pad Vout
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31131 RO2VDD|VDD|anode|cathode|nclk|pad Vout IN|Vout
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31135 Vin$1 RO2VDD|VDD|anode|cathode|nclk|pad IN|Vout
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31136 Vin$2 RO2VDD|VDD|anode|cathode|nclk|pad IN|Vout
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31137 VDD|pad|pin1|supply|vdd i \$247856 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31138 VDD|pad|pin1|supply|vdd \$247856 RD[4]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31139 VDD|pad|pin1|supply|vdd \$248626 \$248626 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31140 VDD|pad|pin1|supply|vdd i$1 \$247857 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31141 VDD|pad|pin1|supply|vdd \$247857 RD[2]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31142 VDD|pad|pin1|supply|vdd R[7]|i|i0|q \$247858 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31143 VDD|pad|pin1|supply|vdd \$247858 RD[39]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31144 \$248627 \$248627 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31145 \$248628 \$248628 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31146 \$248629 \$248629 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31147 VDD|pad|pin1|supply|vdd \$248630 \$248630 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31148 VDD|pad|pin1|supply|vdd \$248631 \$248631 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31149 VDD|pad|pin1|supply|vdd \$249521 RD[26]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31150 VDD|pad|pin1|supply|vdd R[5]|i|i0|q \$247859 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31151 VDD|pad|pin1|supply|vdd \$247859 RD[37]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31152 VDD|pad|pin1|supply|vdd \$248632 \$248632 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31153 VDD|pad|pin1|supply|vdd \$249522 RD[19]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31154 VDD|pad|pin1|supply|vdd \$248633 \$248633 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31155 VDD|pad|pin1|supply|vdd \$248634 \$248634 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31156 VDD|pad|pin1|supply|vdd i$2 \$247860 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31157 VDD|pad|pin1|supply|vdd \$247860 RD[0]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31158 VDD|pad|pin1|supply|vdd \$248635 \$248635 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31159 VDD|pad|pin1|supply|vdd \$249523 RD[17]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31160 VDD|pad|pin1|supply|vdd \$249524 RD[21]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31161 VDD|pad|pin1|supply|vdd R[14]|i|i0|q \$247861 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31162 VDD|pad|pin1|supply|vdd \$247861 RD[46]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31163 VDD|pad|pin1|supply|vdd i$3 \$247862 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31164 VDD|pad|pin1|supply|vdd \$247862 RD[1]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31165 RD[24]|a2|z \$249525 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31166 VDD|pad|pin1|supply|vdd R[12]|i|i0|q \$247863 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31167 VDD|pad|pin1|supply|vdd \$247863 RD[44]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31168 \$248636 \$248636 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31169 RD[28]|a2|z \$249526 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31170 RD[30]|a2|z \$249527 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31171 \$248637 \$248637 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31172 VDD|pad|pin1|supply|vdd i$4 \$247864 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31173 VDD|pad|pin1|supply|vdd \$247864 RD[3]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31174 VDD|pad|pin1|supply|vdd R[15]|i|i0|q \$247865 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31175 VDD|pad|pin1|supply|vdd \$247865 RD[47]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31176 VDD|pad|pin1|supply|vdd \$248638 \$248638 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31177 \$248639 \$248639 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31178 \$248640 \$248640 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31179 VDD|pad|pin1|supply|vdd R[13]|i|i0|q \$247866 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31180 VDD|pad|pin1|supply|vdd \$247866 RD[45]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31181 VDD|pad|pin1|supply|vdd R[4]|i|i0|q \$247867 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31182 VDD|pad|pin1|supply|vdd \$247867 RD[36]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31183 VDD|pad|pin1|supply|vdd R[6]|i|i0|q \$247868 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$31184 VDD|pad|pin1|supply|vdd \$247868 RD[38]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31185 VDD|pad|pin1|supply|vdd DUT_Header|R[11]|Vup|i|i0|q \$247869
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$31186 VDD|pad|pin1|supply|vdd \$247869 RD[43]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31187 VDD|pad|pin1|supply|vdd DUT_Footer|R[2]|Vdn|i|i0|q \$247870
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$31188 VDD|pad|pin1|supply|vdd \$247870 RD[34]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31189 VDD|pad|pin1|supply|vdd DUT_Footer|R[10]|Vdn|i|i0|q \$247871
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$31190 VDD|pad|pin1|supply|vdd \$247871 RD[42]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31191 VDD|pad|pin1|supply|vdd RO_control|R[1]|i|i0|nclk|q \$247872
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$31192 VDD|pad|pin1|supply|vdd \$247872 RD[33]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31193 VDD|pad|pin1|supply|vdd DUT_Header|R[3]|Vup|i|i0|q \$247873
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$31194 VDD|pad|pin1|supply|vdd \$247873 RD[35]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31195 VDD|pad|pin1|supply|vdd R[8]|clk|i|i0|n_RO_control|q \$247874
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$31196 VDD|pad|pin1|supply|vdd \$247874 RD[40]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31197 VDD|pad|pin1|supply|vdd R[0]|clk|i|i0|n_RO_control|q \$247875
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$31198 VDD|pad|pin1|supply|vdd \$247875 RD[32]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31199 VDD|pad|pin1|supply|vdd RO_control|R[9]|i|i0|nclk|q \$247876
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$31200 VDD|pad|pin1|supply|vdd \$247876 RD[41]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$31201 Vin|Vout RO2VDD|VDD|anode|cathode|nclk|pad Vin$3
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31202 Vin|Vout RO2VDD|VDD|anode|cathode|nclk|pad Vin$4
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31203 Vin|Vout Vout$1 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31207 Vout$1 RO2VDD|VDD|anode|cathode|nclk|pad Vin$5
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31208 Vout$1 RO2VDD|VDD|anode|cathode|nclk|pad Vin$6
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31209 Vout$1 Vout$2 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31213 Vout$2 RO2VDD|VDD|anode|cathode|nclk|pad Vin$7
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31214 Vout$2 RO2VDD|VDD|anode|cathode|nclk|pad Vin$8
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31215 Vout$2 Vout$3 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31219 Vout$3 RO2VDD|VDD|anode|cathode|nclk|pad Vin$9
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31220 Vout$3 RO2VDD|VDD|anode|cathode|nclk|pad Vin$10
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31221 Vout$3 Vout$4 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31225 Vout$4 RO2VDD|VDD|anode|cathode|nclk|pad Vin$11
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31226 Vout$4 RO2VDD|VDD|anode|cathode|nclk|pad Vin$12
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31227 Vout$4 Vout$5 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31231 Vout$5 RO2VDD|VDD|anode|cathode|nclk|pad Vin$13
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31232 Vout$5 RO2VDD|VDD|anode|cathode|nclk|pad Vin$14
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31233 Vout$5 Vout$6 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31237 Vout$6 RO2VDD|VDD|anode|cathode|nclk|pad Vin$15
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31238 Vout$6 RO2VDD|VDD|anode|cathode|nclk|pad Vin$16
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31239 Vout$6 Vout$7 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31243 Vout$7 RO2VDD|VDD|anode|cathode|nclk|pad Vin$17
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31244 Vout$7 RO2VDD|VDD|anode|cathode|nclk|pad Vin$18
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31245 Vout$7 Vout$8 RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31249 Vout$8 RO2VDD|VDD|anode|cathode|nclk|pad Vin$19
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31250 Vout$8 RO2VDD|VDD|anode|cathode|nclk|pad Vin$20
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31251 Vout$8 IN|Vout RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31255 \$236455 RESET_B|RSTB|core|p2c RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.147p
+ AD=0.1563p PS=1.54u PD=1.22u
M$31256 RO2VDD|VDD|anode|cathode|nclk|pad \$235757 \$236518
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1563p
+ AD=0.063p PS=1.22u PD=0.72u
M$31257 \$236518 \$235938 \$236455 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.063p AD=0.0798p PS=0.72u PD=0.8u
M$31258 \$236455 \$236468 \$235935 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u PD=1.52u
M$31259 \$236457 RESET_B|RSTB|core|p2c RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.147p
+ AD=0.1563p PS=1.54u PD=1.22u
M$31260 RO2VDD|VDD|anode|cathode|nclk|pad \$235758 \$236516
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1563p
+ AD=0.063p PS=1.22u PD=0.72u
M$31261 \$236516 \$235946 \$236457 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.063p AD=0.0798p PS=0.72u PD=0.8u
M$31262 \$236457 \$236469 \$235943 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u PD=1.52u
M$31263 \$236459 RESET_B|RSTB|core|p2c RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.147p
+ AD=0.1563p PS=1.54u PD=1.22u
M$31264 RO2VDD|VDD|anode|cathode|nclk|pad \$235759 \$236514
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1563p
+ AD=0.063p PS=1.22u PD=0.72u
M$31265 \$236514 \$235954 \$236459 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.063p AD=0.0798p PS=0.72u PD=0.8u
M$31266 \$236459 \$236470 \$235951 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u PD=1.52u
M$31267 \$236461 RESET_B|RSTB|core|p2c RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.147p
+ AD=0.1563p PS=1.54u PD=1.22u
M$31268 RO2VDD|VDD|anode|cathode|nclk|pad \$235760 \$236512
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1563p
+ AD=0.063p PS=1.22u PD=0.72u
M$31269 \$236512 \$235962 \$236461 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.063p AD=0.0798p PS=0.72u PD=0.8u
M$31270 \$236461 \$236471 \$235959 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u PD=1.52u
M$31271 \$236463 RESET_B|RSTB|core|p2c RO2VDD|VDD|anode|cathode|nclk|pad
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.147p
+ AD=0.1563p PS=1.54u PD=1.22u
M$31272 RO2VDD|VDD|anode|cathode|nclk|pad \$235761 \$236510
+ RO2VDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1563p
+ AD=0.063p PS=1.22u PD=0.72u
M$31273 \$236510 \$235970 \$236463 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.063p AD=0.0798p PS=0.72u PD=0.8u
M$31274 \$236463 \$236472 \$235967 RO2VDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p PS=0.8u PD=1.52u
M$31275 VDD|pad|pin1|supply|vdd \$252776 DUT_gate|core|p2c
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$31276 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$1 Vin|Vout$2
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31280 Vin$21 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$2
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31281 Vin$22 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$2
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31282 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$2 Vin|Vout$3
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31286 Vin$23 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$3
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31287 Vin$24 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$3
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31288 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$3 Vin|Vout$4
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31292 Vin$25 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$4
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31293 Vin$26 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$4
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31294 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$4 Vin|Vout$5
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31298 Vin$27 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$5
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31299 Vin$28 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$5
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31300 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$5 Vin|Vout$6
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31304 Vin$29 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$6
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31305 Vin$30 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$6
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31306 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$6 Vin|Vout$7
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31310 Vin$31 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$7
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31311 Vin$32 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$7
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31312 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$7 Vin|Vout$8
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31316 Vin$33 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$8
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31317 Vin$34 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$8
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31318 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$8 Vin|Vout$9
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31322 Vin$35 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$9
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31323 Vin$36 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$9
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31324 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$9 Vin|Vout$10
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31328 Vin$37 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$10
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31329 Vin$38 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$10
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31330 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$10 Vin|Vout$11
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31334 Vin$39 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$11
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31335 Vin$40 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$11
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31336 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$11 Vin|Vout$12
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31340 Vin$41 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$12
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31341 Vin$42 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$12
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31342 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$12 Vin|Vout$13
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31346 Vin$43 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$13
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31347 Vin$44 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$13
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31348 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$13 Vin|Vout$14
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31352 Vin$45 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$14
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31353 Vin$46 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$14
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31354 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$14 Vin|Vout$15
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31358 Vin$47 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$15
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31359 Vin$48 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$15
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31360 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$15 Vin|Vout$16
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31364 Vin$49 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$16
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31365 VDD|pad|pin1|supply|vdd \$250730 \$250730 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31366 Vin$50 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$16
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31367 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$16 Vin|Vout$17
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31371 VDD|pad|pin1|supply|vdd \$250731 \$250731 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31372 Vin$51 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$17
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31373 Vin$52 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$17
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31374 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$17 Vin|Vout$18
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31377 RD[23]|a4|z \$249966 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$31379 Vin$53 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$18
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31380 Vin$54 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$18
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31381 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$18 Vin|Vout$19
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31385 Vin$55 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$19
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31386 Vin$56 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$19
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31387 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$19 Vin|Vout$20
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31391 Vin$57 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$20
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31392 Vin$58 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$20
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31393 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$20 Vin|Vout$21
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31397 Vin$59 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$21
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31398 Vin$60 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$21
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31399 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$21 Vin|Vout$22
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31403 Vin$61 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$22
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31404 Vin$62 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$22
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31405 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$22 Vin|Vout$23
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31409 Vin$63 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$23
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31410 Vin$64 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$23
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31411 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$23 Vin|Vout$24
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31415 Vin$65 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$24
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31416 Vin$66 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$24
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31417 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$24 Vin|Vout$25
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31421 Vin$67 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$25
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31422 Vin$68 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$25
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31423 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$25 Vin|Vout$26
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31427 Vin$69 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$26
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31428 Vin$70 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$26
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31429 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$26 Vin|Vout$27
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31433 Vin$71 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$27
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31434 Vin$72 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$27
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31435 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$27 Vin|Vout$28
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31439 Vin$73 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$28
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31440 Vin$74 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$28
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31441 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$28 Vin|Vout$29
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31445 Vin$75 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$29
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31446 Vin$76 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$29
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31447 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$29 Vin|Vout$30
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31451 Vin$77 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$30
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31452 Vin$78 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$30
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31453 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$30 Vin|Vout$31
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31457 Vin$79 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$31
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31458 Vin$80 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$31
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31459 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$31 Vin|Vout$32
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31463 Vin$81 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$32
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31464 Vin$82 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$32
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31465 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$32 Vin|Vout$33
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31469 Vin$83 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$33
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31470 Vin$84 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$33
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31471 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$33 Vin|Vout$34
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31475 Vin$85 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$34
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31476 Vin$86 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$34
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31477 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$34 Vin|Vout$35
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31481 Vin$87 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$35
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31482 Vin$88 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$35
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31483 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$35 Vin|Vout$36
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31487 Vin$89 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$36
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31488 Vin$90 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$36
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31489 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$36 Vin|Vout$37
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31493 Vin$91 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$37
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31494 Vin$92 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$37
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31495 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$37 Vin|Vout$38
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31499 Vin$93 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$38
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31500 Vin$94 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$38
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31501 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$38 Vin|Vout$39
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31505 Vin$95 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$39
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31506 Vin$96 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$39
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31507 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$39 Vin|Vout$40
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31511 Vin$97 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$40
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31512 Vin$98 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$40
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31513 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$40 Vin|Vout$41
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31517 Vin$99 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$41
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31518 Vin$100 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$41
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31519 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$41 Vin|Vout$42
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31523 Vin$101 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$42
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31524 Vin$102 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$42
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31525 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$42 Vin|Vout$43
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31529 Vin$103 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$43
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31530 Vin$104 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$43
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31531 ROVDD|VDD|anode|cathode|nclk|pad Vin|Vout$43 Vout$9
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31535 Vin$105 ROVDD|VDD|anode|cathode|nclk|pad Vout$9
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31536 Vin$106 ROVDD|VDD|anode|cathode|nclk|pad Vout$9
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31537 \$271052 R[0]|clk|i|i0|n_RO_control|q ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=40.8u AS=13.872p
+ AD=13.872p PS=89.76u PD=89.76u
M$31549 \$271052 Vout$9 Vin$107 ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos
+ L=0.45u W=13.6u AS=4.624p AD=4.624p PS=29.92u PD=29.92u
M$31553 Vin$107 RO_control|R[1]|i|i0|nclk|q \$270153
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31554 Vin$107 RO_control|R[1]|i|i0|nclk|q DUT_gate|core|p2c
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31555 \$271053 DUT_Header|R[3]|Vup|i|i0|q ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=40.8u AS=13.872p
+ AD=13.872p PS=89.76u PD=89.76u
M$31567 \$271053 Vin$107 Vin|Vout|core|extra_load|padres$1
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31571 Vin|Vout|core|extra_load|padres$1 RO_control|R[1]|i|i0|nclk|q
+ Drain_Sense|Vout|core|padres$1 ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos
+ L=0.45u W=3.4u AS=1.156p AD=1.156p PS=7.48u PD=7.48u
M$31572 Vin|Vout|core|extra_load|padres$1 RO_control|R[1]|i|i0|nclk|q
+ Drain_Force|Vout|core|padres$1 ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos
+ L=0.45u W=13.6u AS=4.624p AD=4.624p PS=29.92u PD=29.92u
M$31576 ROVDD|VDD|anode|cathode|nclk|pad R[0]|clk|i|i0|n_RO_control|q \$271054
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=40.8u AS=13.872p
+ AD=13.872p PS=89.76u PD=89.76u
M$31588 \$271054 Vin|Vout|core|extra_load|padres$1 Vin$110
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31592 \$270157 ROVDD|VDD|anode|cathode|nclk|pad Vin$110
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31593 VSS|anode|cathode|clk|vss ROVDD|VDD|anode|cathode|nclk|pad Vin$110
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31594 ROVDD|VDD|anode|cathode|nclk|pad Vin$110 IN|Vin|Vout
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31598 Vin$108 ROVDD|VDD|anode|cathode|nclk|pad IN|Vin|Vout
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31599 Vin$109 ROVDD|VDD|anode|cathode|nclk|pad IN|Vin|Vout
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31600 CLK|core|i|p2c$1 \$254718 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$31601 Vin|Vout$1 ROVDD|VDD|anode|cathode|nclk|pad Vin$111
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31602 Vin|Vout$1 ROVDD|VDD|anode|cathode|nclk|pad Vin$112
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31603 Vin|Vout$1 Vin|Vout$44 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31607 Vin|Vout$44 ROVDD|VDD|anode|cathode|nclk|pad Vin$113
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31608 Vin|Vout$44 ROVDD|VDD|anode|cathode|nclk|pad Vin$114
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31609 Vin|Vout$44 Vin|Vout$45 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31613 Vin|Vout$45 ROVDD|VDD|anode|cathode|nclk|pad Vin$115
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31614 Vin|Vout$45 ROVDD|VDD|anode|cathode|nclk|pad Vin$116
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31615 Vin|Vout$45 Vin|Vout$46 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31619 Vin|Vout$46 ROVDD|VDD|anode|cathode|nclk|pad Vin$117
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31620 Vin|Vout$46 ROVDD|VDD|anode|cathode|nclk|pad Vin$118
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31621 Vin|Vout$46 Vin|Vout$47 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31625 Vin|Vout$47 ROVDD|VDD|anode|cathode|nclk|pad Vin$119
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31626 Vin|Vout$47 ROVDD|VDD|anode|cathode|nclk|pad Vin$120
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31627 Vin|Vout$47 Vin|Vout$48 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31631 Vin|Vout$48 ROVDD|VDD|anode|cathode|nclk|pad Vin$121
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31632 Vin|Vout$48 ROVDD|VDD|anode|cathode|nclk|pad Vin$122
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31633 Vin|Vout$48 Vin|Vout$49 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31637 Vin|Vout$49 ROVDD|VDD|anode|cathode|nclk|pad Vin$123
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31638 Vin|Vout$49 ROVDD|VDD|anode|cathode|nclk|pad Vin$124
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31639 Vin|Vout$49 Vin|Vout$50 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31643 Vin|Vout$50 ROVDD|VDD|anode|cathode|nclk|pad Vin$125
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31644 Vin|Vout$50 ROVDD|VDD|anode|cathode|nclk|pad Vin$126
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31645 Vin|Vout$50 Vin|Vout$51 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31649 Vin|Vout$51 ROVDD|VDD|anode|cathode|nclk|pad Vin$127
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31650 Vin|Vout$51 ROVDD|VDD|anode|cathode|nclk|pad Vin$128
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31651 Vin|Vout$51 Vin|Vout$52 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31655 Vin|Vout$52 ROVDD|VDD|anode|cathode|nclk|pad Vin$129
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31656 Vin|Vout$52 ROVDD|VDD|anode|cathode|nclk|pad Vin$130
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31657 Vin|Vout$52 Vin|Vout$53 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31661 Vin|Vout$53 ROVDD|VDD|anode|cathode|nclk|pad Vin$131
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31662 Vin|Vout$53 ROVDD|VDD|anode|cathode|nclk|pad Vin$132
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31663 Vin|Vout$53 Vin|Vout$54 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31667 Vin|Vout$54 ROVDD|VDD|anode|cathode|nclk|pad Vin$133
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31668 Vin|Vout$54 ROVDD|VDD|anode|cathode|nclk|pad Vin$134
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31669 Vin|Vout$54 Vin|Vout$55 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31673 Vin|Vout$55 ROVDD|VDD|anode|cathode|nclk|pad Vin$135
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31674 Vin|Vout$55 ROVDD|VDD|anode|cathode|nclk|pad Vin$136
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31675 Vin|Vout$55 Vin|Vout$56 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31679 Vin|Vout$56 ROVDD|VDD|anode|cathode|nclk|pad Vin$137
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31680 Vin|Vout$56 ROVDD|VDD|anode|cathode|nclk|pad Vin$138
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31681 Vin|Vout$56 Vin|Vout$57 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31685 Vin|Vout$57 ROVDD|VDD|anode|cathode|nclk|pad Vin$139
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31686 Vin|Vout$57 ROVDD|VDD|anode|cathode|nclk|pad Vin$140
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31687 Vin|Vout$57 Vin|Vout$58 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31691 Vin|Vout$58 ROVDD|VDD|anode|cathode|nclk|pad Vin$141
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31692 Vin|Vout$58 ROVDD|VDD|anode|cathode|nclk|pad Vin$142
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31693 Vin|Vout$58 Vin|Vout$59 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31697 Vin|Vout$59 ROVDD|VDD|anode|cathode|nclk|pad Vin$143
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31698 Vin|Vout$59 ROVDD|VDD|anode|cathode|nclk|pad Vin$144
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31699 Vin|Vout$59 Vin|Vout$60 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31703 Vin|Vout$60 ROVDD|VDD|anode|cathode|nclk|pad Vin$145
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31704 Vin|Vout$60 ROVDD|VDD|anode|cathode|nclk|pad Vin$146
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31705 Vin|Vout$60 Vin|Vout$61 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31709 Vin|Vout$61 ROVDD|VDD|anode|cathode|nclk|pad Vin$147
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31710 Vin|Vout$61 ROVDD|VDD|anode|cathode|nclk|pad Vin$148
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31711 Vin|Vout$61 Vin|Vout$62 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31715 Vin|Vout$62 ROVDD|VDD|anode|cathode|nclk|pad Vin$149
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31716 Vin|Vout$62 ROVDD|VDD|anode|cathode|nclk|pad Vin$150
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31717 Vin|Vout$62 Vin|Vout$63 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31721 Vin|Vout$63 ROVDD|VDD|anode|cathode|nclk|pad Vin$151
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31722 Vin|Vout$63 ROVDD|VDD|anode|cathode|nclk|pad Vin$152
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31723 Vin|Vout$63 Vin|Vout$64 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31727 Vin|Vout$64 ROVDD|VDD|anode|cathode|nclk|pad Vin$153
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31728 Vin|Vout$64 ROVDD|VDD|anode|cathode|nclk|pad Vin$154
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31729 Vin|Vout$64 Vin|Vout$65 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31733 Vin|Vout$65 ROVDD|VDD|anode|cathode|nclk|pad Vin$155
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31734 Vin|Vout$65 ROVDD|VDD|anode|cathode|nclk|pad Vin$156
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31735 Vin|Vout$65 Vin|Vout$66 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31739 Vin|Vout$66 ROVDD|VDD|anode|cathode|nclk|pad Vin$157
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31740 Vin|Vout$66 ROVDD|VDD|anode|cathode|nclk|pad Vin$158
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31741 Vin|Vout$66 Vin|Vout$67 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31745 Vin|Vout$67 ROVDD|VDD|anode|cathode|nclk|pad Vin$159
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31746 Vin|Vout$67 ROVDD|VDD|anode|cathode|nclk|pad Vin$160
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31747 Vin|Vout$67 Vin|Vout$68 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31751 Vin|Vout$68 ROVDD|VDD|anode|cathode|nclk|pad Vin$161
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31752 Vin|Vout$68 ROVDD|VDD|anode|cathode|nclk|pad Vin$162
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31753 Vin|Vout$68 Vin|Vout$69 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31757 Vin|Vout$69 ROVDD|VDD|anode|cathode|nclk|pad Vin$163
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31758 Vin|Vout$69 ROVDD|VDD|anode|cathode|nclk|pad Vin$164
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31759 Vin|Vout$69 Vin|Vout$70 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31763 Vin|Vout$70 ROVDD|VDD|anode|cathode|nclk|pad Vin$165
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31764 Vin|Vout$70 ROVDD|VDD|anode|cathode|nclk|pad Vin$166
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31765 Vin|Vout$70 Vin|Vout$71 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31769 Vin|Vout$71 ROVDD|VDD|anode|cathode|nclk|pad Vin$167
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31770 Vin|Vout$71 ROVDD|VDD|anode|cathode|nclk|pad Vin$168
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31771 Vin|Vout$71 Vin|Vout$72 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31775 Vin|Vout$72 ROVDD|VDD|anode|cathode|nclk|pad Vin$169
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31776 Vin|Vout$72 ROVDD|VDD|anode|cathode|nclk|pad Vin$170
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31777 Vin|Vout$72 Vin|Vout$73 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31781 Vin|Vout$73 ROVDD|VDD|anode|cathode|nclk|pad Vin$171
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31782 Vin|Vout$73 ROVDD|VDD|anode|cathode|nclk|pad Vin$172
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31783 Vin|Vout$73 Vin|Vout$74 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31787 Vin|Vout$74 ROVDD|VDD|anode|cathode|nclk|pad Vin$173
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31788 Vin|Vout$74 ROVDD|VDD|anode|cathode|nclk|pad Vin$174
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31789 Vin|Vout$74 Vin|Vout$75 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31793 Vin|Vout$75 ROVDD|VDD|anode|cathode|nclk|pad Vin$175
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31794 Vin|Vout$75 ROVDD|VDD|anode|cathode|nclk|pad Vin$176
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31795 Vin|Vout$75 Vin|Vout$76 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31799 Vin|Vout$76 ROVDD|VDD|anode|cathode|nclk|pad Vin$177
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31800 Vin|Vout$76 ROVDD|VDD|anode|cathode|nclk|pad Vin$178
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31801 Vin|Vout$76 Vin|Vout$77 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31805 Vin|Vout$77 ROVDD|VDD|anode|cathode|nclk|pad Vin$179
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31806 Vin|Vout$77 ROVDD|VDD|anode|cathode|nclk|pad Vin$180
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31807 Vin|Vout$77 Vin|Vout$78 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31811 Vin|Vout$78 ROVDD|VDD|anode|cathode|nclk|pad Vin$181
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31812 Vin|Vout$78 ROVDD|VDD|anode|cathode|nclk|pad Vin$182
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31813 Vin|Vout$78 Vin|Vout$79 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31817 Vin|Vout$79 ROVDD|VDD|anode|cathode|nclk|pad Vin$183
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31818 Vin|Vout$79 ROVDD|VDD|anode|cathode|nclk|pad Vin$184
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31819 Vin|Vout$79 Vin|Vout$80 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31823 Vin|Vout$80 ROVDD|VDD|anode|cathode|nclk|pad Vin$185
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31824 Vin|Vout$80 ROVDD|VDD|anode|cathode|nclk|pad Vin$186
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31825 Vin|Vout$80 Vin|Vout$81 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31829 Vin|Vout$81 ROVDD|VDD|anode|cathode|nclk|pad Vin$187
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31830 Vin|Vout$81 ROVDD|VDD|anode|cathode|nclk|pad Vin$188
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31831 Vin|Vout$81 Vin|Vout$82 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31835 Vin|Vout$82 ROVDD|VDD|anode|cathode|nclk|pad Vin$189
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31836 Vin|Vout$82 ROVDD|VDD|anode|cathode|nclk|pad Vin$190
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31837 Vin|Vout$82 Vin|Vout$83 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31841 Vin|Vout$83 ROVDD|VDD|anode|cathode|nclk|pad Vin$191
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31842 Vin|Vout$83 ROVDD|VDD|anode|cathode|nclk|pad Vin$192
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31843 Vin|Vout$83 Vin|Vout$84 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31847 Vin|Vout$84 ROVDD|VDD|anode|cathode|nclk|pad Vin$193
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31848 Vin|Vout$84 ROVDD|VDD|anode|cathode|nclk|pad Vin$194
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31849 Vin|Vout$84 Vin|Vout$85 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31853 Vin|Vout$85 ROVDD|VDD|anode|cathode|nclk|pad Vin$195
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31854 Vin|Vout$85 ROVDD|VDD|anode|cathode|nclk|pad Vin$196
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31855 Vin|Vout$85 Vin|Vout$86 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31859 Vin|Vout$86 ROVDD|VDD|anode|cathode|nclk|pad Vin$197
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31860 Vin|Vout$86 ROVDD|VDD|anode|cathode|nclk|pad Vin$198
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31861 Vin|Vout$86 Vin|Vout$87 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31865 Vin|Vout$87 ROVDD|VDD|anode|cathode|nclk|pad Vin$199
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31866 Vin|Vout$87 ROVDD|VDD|anode|cathode|nclk|pad Vin$200
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31867 Vin|Vout$87 Vin|Vout$88 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31871 Vin|Vout$88 ROVDD|VDD|anode|cathode|nclk|pad Vin$201
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31872 Vin|Vout$88 ROVDD|VDD|anode|cathode|nclk|pad Vin$202
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31873 Vin|Vout$88 Vin|Vout$89 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31877 Vin|Vout$89 ROVDD|VDD|anode|cathode|nclk|pad Vin$203
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31878 Vin|Vout$89 ROVDD|VDD|anode|cathode|nclk|pad Vin$204
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31879 Vin|Vout$89 Vin|Vout$90 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31883 Vin|Vout$90 ROVDD|VDD|anode|cathode|nclk|pad Vin$205
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31884 Vin|Vout$90 ROVDD|VDD|anode|cathode|nclk|pad Vin$206
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31885 Vin|Vout$90 Vin|Vout$91 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31889 Vin|Vout$91 ROVDD|VDD|anode|cathode|nclk|pad Vin$207
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31890 Vin|Vout$91 ROVDD|VDD|anode|cathode|nclk|pad Vin$208
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31891 Vin|Vout$91 Vin|Vout$92 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31895 Vin|Vout$92 ROVDD|VDD|anode|cathode|nclk|pad Vin$209
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31896 Vin|Vout$92 ROVDD|VDD|anode|cathode|nclk|pad Vin$210
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31897 Vin|Vout$92 Vin|Vout$93 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31901 Vin|Vout$93 ROVDD|VDD|anode|cathode|nclk|pad Vin$211
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31902 Vin|Vout$93 ROVDD|VDD|anode|cathode|nclk|pad Vin$212
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31903 Vin|Vout$93 Vin|Vout$94 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31907 Vin|Vout$94 ROVDD|VDD|anode|cathode|nclk|pad Vin$213
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31908 Vin|Vout$94 ROVDD|VDD|anode|cathode|nclk|pad Vin$214
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31909 Vin|Vout$94 Vin|Vout$95 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31913 Vin|Vout$95 ROVDD|VDD|anode|cathode|nclk|pad Vin$215
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31914 Vin|Vout$95 ROVDD|VDD|anode|cathode|nclk|pad Vin$216
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31915 Vin|Vout$95 Vin|Vout$96 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31919 Vin|Vout$96 ROVDD|VDD|anode|cathode|nclk|pad Vin$217
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31920 Vin|Vout$96 ROVDD|VDD|anode|cathode|nclk|pad Vin$218
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=3.4u AS=1.156p
+ AD=1.156p PS=7.48u PD=7.48u
M$31921 Vin|Vout$96 IN|Vin|Vout ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.45u W=13.6u AS=4.624p
+ AD=4.624p PS=29.92u PD=29.92u
M$31925 VDD|pad|pin1|supply|vdd \$278874 DUT_gate|core|p2c$1
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$31926 VDD|pad|pin1|supply|vdd OUT|Q|c2p|core|i$1 \$304122
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$31927 OUT|Q|c2p|core|i$1 \$279336 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p
+ AD=0.2128p PS=2.92u PD=1.5u
M$31928 ROVDD|VDD|anode|cathode|nclk|pad \$279856 \$279336
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p
+ AD=0.3864p PS=1.5u PD=2.93u
M$31929 ROVDD|VDD|anode|cathode|nclk|pad \$279856 \$279338
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.2639p
+ AD=0.0798p PS=1.81u PD=0.8u
M$31930 \$279338 RESET_B|RSTB|core|p2c ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p
+ AD=0.204p PS=0.8u PD=1.835u
M$31931 ROVDD|VDD|anode|cathode|nclk|pad \$279338 \$280132
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.204p
+ AD=0.09345p PS=1.835u PD=0.865u
M$31932 \$280132 \$279857 \$279856 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.09345p AD=0.2048p PS=0.865u PD=1.63u
M$31933 \$279856 \$279562 \$279340 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=1u AS=0.2048p AD=0.34p PS=1.63u PD=2.68u
M$31934 D|Q_N$5 \$279856 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.4312p
+ AD=0.2639p PS=3.01u PD=1.81u
M$31935 VDD|pad|pin1|supply|vdd OUT|Q|c2p|core|i$1 \$304123
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$31936 \$279562 Q$4 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.4088p
+ AD=0.41165p PS=2.97u PD=2.12u
M$31937 ROVDD|VDD|anode|cathode|nclk|pad \$279562 \$279857
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.41165p
+ AD=0.3864p PS=2.12u PD=2.93u
M$31938 \$279563 \$279857 \$279859 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u PD=0.8u
M$31939 \$279859 \$279562 \$280658 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.063p PS=0.8u PD=0.72u
M$31940 \$280658 \$279340 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.063p
+ AD=0.1563p PS=0.72u PD=1.22u
M$31941 ROVDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$279859
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1563p
+ AD=0.147p PS=1.22u PD=1.54u
M$31942 ROVDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$279563
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.3623875p
+ AD=0.0798p PS=2.605u PD=0.8u
M$31943 \$279563 D|Q_N$5 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$31944 \$279340 \$279859 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1u AS=0.34p
+ AD=0.3623875p PS=2.68u PD=2.605u
M$31945 Q$4 \$279341 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p
+ AD=0.2128p PS=2.92u PD=1.5u
M$31946 ROVDD|VDD|anode|cathode|nclk|pad \$279860 \$279341
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p
+ AD=0.3864p PS=1.5u PD=2.93u
M$31947 ROVDD|VDD|anode|cathode|nclk|pad \$279860 \$279343
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.2639p
+ AD=0.0798p PS=1.81u PD=0.8u
M$31948 \$279343 RESET_B|RSTB|core|p2c ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p
+ AD=0.204p PS=0.8u PD=1.835u
M$31949 ROVDD|VDD|anode|cathode|nclk|pad \$279343 \$280124
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.204p
+ AD=0.09345p PS=1.835u PD=0.865u
M$31950 \$280124 \$279861 \$279860 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.09345p AD=0.2048p PS=0.865u PD=1.63u
M$31951 \$279860 \$279565 \$279345 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=1u AS=0.2048p AD=0.34p PS=1.63u PD=2.68u
M$31952 D|Q_N$6 \$279860 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.4312p
+ AD=0.2639p PS=3.01u PD=1.81u
M$31953 \$279565 Q$5 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.4088p
+ AD=0.41165p PS=2.97u PD=2.12u
M$31954 ROVDD|VDD|anode|cathode|nclk|pad \$279565 \$279861
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.41165p
+ AD=0.3864p PS=2.12u PD=2.93u
M$31955 \$279566 \$279861 \$279863 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u PD=0.8u
M$31956 \$279863 \$279565 \$280667 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.063p PS=0.8u PD=0.72u
M$31957 \$280667 \$279345 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.063p
+ AD=0.1563p PS=0.72u PD=1.22u
M$31958 ROVDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$279863
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1563p
+ AD=0.147p PS=1.22u PD=1.54u
M$31959 ROVDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$279566
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.3623875p
+ AD=0.0798p PS=2.605u PD=0.8u
M$31960 \$279566 D|Q_N$6 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$31961 \$279345 \$279863 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1u AS=0.34p
+ AD=0.3623875p PS=2.68u PD=2.605u
M$31962 Q$5 \$279346 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p
+ AD=0.2128p PS=2.92u PD=1.5u
M$31963 ROVDD|VDD|anode|cathode|nclk|pad \$279864 \$279346
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p
+ AD=0.3864p PS=1.5u PD=2.93u
M$31964 ROVDD|VDD|anode|cathode|nclk|pad \$279864 \$279348
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.2639p
+ AD=0.0798p PS=1.81u PD=0.8u
M$31965 \$279348 RESET_B|RSTB|core|p2c ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p
+ AD=0.204p PS=0.8u PD=1.835u
M$31966 ROVDD|VDD|anode|cathode|nclk|pad \$279348 \$280117
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.204p
+ AD=0.09345p PS=1.835u PD=0.865u
M$31967 \$280117 \$279865 \$279864 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.09345p AD=0.2048p PS=0.865u PD=1.63u
M$31968 \$279864 \$279568 \$279350 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=1u AS=0.2048p AD=0.34p PS=1.63u PD=2.68u
M$31969 D|Q_N$7 \$279864 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.4312p
+ AD=0.2639p PS=3.01u PD=1.81u
M$31970 \$279568 Q$6 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.4088p
+ AD=0.41165p PS=2.97u PD=2.12u
M$31971 ROVDD|VDD|anode|cathode|nclk|pad \$279568 \$279865
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.41165p
+ AD=0.3864p PS=2.12u PD=2.93u
M$31972 \$279569 \$279865 \$279867 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u PD=0.8u
M$31973 \$279867 \$279568 \$280673 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.063p PS=0.8u PD=0.72u
M$31974 \$280673 \$279350 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.063p
+ AD=0.1563p PS=0.72u PD=1.22u
M$31975 ROVDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$279867
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1563p
+ AD=0.147p PS=1.22u PD=1.54u
M$31976 ROVDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$279569
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.3623875p
+ AD=0.0798p PS=2.605u PD=0.8u
M$31977 \$279569 D|Q_N$7 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$31978 \$279350 \$279867 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1u AS=0.34p
+ AD=0.3623875p PS=2.68u PD=2.605u
M$31979 Q$6 \$279351 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p
+ AD=0.2128p PS=2.92u PD=1.5u
M$31980 ROVDD|VDD|anode|cathode|nclk|pad \$279868 \$279351
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p
+ AD=0.3864p PS=1.5u PD=2.93u
M$31981 ROVDD|VDD|anode|cathode|nclk|pad \$279868 \$279353
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.2639p
+ AD=0.0798p PS=1.81u PD=0.8u
M$31982 \$279353 RESET_B|RSTB|core|p2c ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p
+ AD=0.204p PS=0.8u PD=1.835u
M$31983 ROVDD|VDD|anode|cathode|nclk|pad \$279353 \$280109
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.204p
+ AD=0.09345p PS=1.835u PD=0.865u
M$31984 \$280109 \$279869 \$279868 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.09345p AD=0.2048p PS=0.865u PD=1.63u
M$31985 \$279868 \$279571 \$279355 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=1u AS=0.2048p AD=0.34p PS=1.63u PD=2.68u
M$31986 D|Q_N$8 \$279868 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.4312p
+ AD=0.2639p PS=3.01u PD=1.81u
M$31987 \$279571 Q$7 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.4088p
+ AD=0.41165p PS=2.97u PD=2.12u
M$31988 ROVDD|VDD|anode|cathode|nclk|pad \$279571 \$279869
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.41165p
+ AD=0.3864p PS=2.12u PD=2.93u
M$31989 \$279572 \$279869 \$279871 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u PD=0.8u
M$31990 \$279871 \$279571 \$280681 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.063p PS=0.8u PD=0.72u
M$31991 \$280681 \$279355 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.063p
+ AD=0.1563p PS=0.72u PD=1.22u
M$31992 ROVDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$279871
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1563p
+ AD=0.147p PS=1.22u PD=1.54u
M$31993 ROVDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$279572
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.3623875p
+ AD=0.0798p PS=2.605u PD=0.8u
M$31994 \$279572 D|Q_N$8 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$31995 \$279355 \$279871 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1u AS=0.34p
+ AD=0.3623875p PS=2.68u PD=2.605u
M$31996 Q$7 \$279356 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p
+ AD=0.2128p PS=2.92u PD=1.5u
M$31997 ROVDD|VDD|anode|cathode|nclk|pad \$279872 \$279356
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p
+ AD=0.3864p PS=1.5u PD=2.93u
M$31998 ROVDD|VDD|anode|cathode|nclk|pad \$279872 \$279358
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.2639p
+ AD=0.0798p PS=1.81u PD=0.8u
M$31999 \$279358 RESET_B|RSTB|core|p2c ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p
+ AD=0.204p PS=0.8u PD=1.835u
M$32000 ROVDD|VDD|anode|cathode|nclk|pad \$279358 \$280098
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.204p
+ AD=0.09345p PS=1.835u PD=0.865u
M$32001 \$280098 \$279873 \$279872 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.09345p AD=0.2048p PS=0.865u PD=1.63u
M$32002 \$279872 \$279574 \$279360 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=1u AS=0.2048p AD=0.34p PS=1.63u PD=2.68u
M$32003 D|Q_N$9 \$279872 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.4312p
+ AD=0.2639p PS=3.01u PD=1.81u
M$32004 \$279574 IN|Vin|Vout ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.4088p
+ AD=0.41165p PS=2.97u PD=2.12u
M$32005 ROVDD|VDD|anode|cathode|nclk|pad \$279574 \$279873
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1.12u AS=0.41165p
+ AD=0.3864p PS=2.12u PD=2.93u
M$32006 \$279575 \$279873 \$279874 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u PD=0.8u
M$32007 \$279874 \$279574 \$280692 ROVDD|VDD|anode|cathode|nclk|pad
+ sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.063p PS=0.8u PD=0.72u
M$32008 \$280692 \$279360 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.063p
+ AD=0.1563p PS=0.72u PD=1.22u
M$32009 ROVDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$279874
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.1563p
+ AD=0.147p PS=1.22u PD=1.54u
M$32010 ROVDD|VDD|anode|cathode|nclk|pad RESET_B|RSTB|core|p2c \$279575
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.3623875p
+ AD=0.0798p PS=2.605u PD=0.8u
M$32011 \$279575 D|Q_N$9 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$32012 \$279360 \$279874 ROVDD|VDD|anode|cathode|nclk|pad
+ ROVDD|VDD|anode|cathode|nclk|pad sg13_lv_pmos L=0.13u W=1u AS=0.34p
+ AD=0.3623875p PS=2.68u PD=2.605u
M$32013 VDD|pad|pin1|supply|vdd OUT|Q|c2p|core|i \$304124
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$32014 VDD|pad|pin1|supply|vdd OUT|Q|c2p|core|i \$304125
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$32015 CEB|a1|core|i|p2c \$280694 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$32016 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$50381
+ AVDD|anode|cathode|pad|vdd VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32036 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate
+ anode|cathode|pad|pad_adc_result_0_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$32044 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$1
+ anode|cathode|pad|pad_adc_result_1_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$32052 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$2
+ anode|cathode|pad|pad_adc_result_2_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$32060 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$3
+ anode|cathode|pad|pad_adc_result_3_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$32068 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$4
+ anode|cathode|pad|pad_adc_result_4_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$32076 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$5
+ anode|cathode|pad|pad_adc_valid_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=106.56u AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$32084 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$6
+ anode|cathode|pad|pad_adc_sample_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$32168 VDD|pad|pin1|supply|vdd core \$64422 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$32169 VDD|pad|pin1|supply|vdd core$1 \$64424 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$32170 \$63424 \$63425 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32171 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63424 \$63425
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32172 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63425 gate|ngate|o
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32173 \$63426 \$63427 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32174 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63426 \$63427
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32175 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63427 gate|o|pgate
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32176 \$63428 \$63429 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32177 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63428 \$63429
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32178 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63429 gate|ngate|o$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32179 \$63430 \$63431 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32180 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63430 \$63431
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32181 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63431 gate|o|pgate$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32182 \$63432 \$63433 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32183 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63432 \$63433
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32184 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63433 gate|ngate|o$2
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32185 \$63434 \$63435 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32186 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63434 \$63435
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32187 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63435 gate|o|pgate$2
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32188 \$63436 \$63437 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32189 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63436 \$63437
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32190 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63437 gate|ngate|o$3
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32191 \$63438 \$63439 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32192 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63438 \$63439
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32193 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63439 gate|o|pgate$3
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32194 \$63440 \$63441 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32195 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63440 \$63441
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32196 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63441 gate|ngate|o$4
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32197 \$63442 \$63443 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32198 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63442 \$63443
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32199 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63443 gate|o|pgate$4
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32200 \$63444 \$63445 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32201 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63444 \$63445
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32202 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63445 gate|ngate|o$5
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32203 \$63446 \$63447 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32204 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63446 \$63447
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32205 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63447 gate|o|pgate$5
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32206 \$63448 \$63449 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32207 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63448 \$63449
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32208 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63449 gate|ngate|o$6
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32209 \$63450 \$63451 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32210 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63450 \$63451
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32211 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63451 gate|o|pgate$6
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32212 VDD|pad|pin1|supply|vdd core$2 \$90525 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$32213 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$106976
+ anode|cathode|pad|pad_adc_vrefp_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32253 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$127370
+ anode|cathode|pad|pad_adc_vrefn_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32293 VDD|pad|pin1|supply|vdd in|pin2 gate|out VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.5u W=350u AS=67.55p AD=67.55p PS=376.3u PD=376.3u
M$32343 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$144245
+ anode|cathode|pad|pad_adc_vin_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32383 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$168331
+ anode|cathode|pad|pad_adc_vip_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32423 VDDIO|cathode|guard|iovdd|pad|pin1|supply in|pin2$1 gate|out$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.5u W=350u
+ AS=67.55p AD=67.55p PS=376.3u PD=376.3u
M$32473 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$7
+ anode|cathode|pad|pad_miso_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=106.56u AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$32489 \$198890 \$199478 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32490 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$198890 \$199478
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32491 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$199478 gate|ngate|o$7
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32492 \$200225 \$200540 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32493 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$200225 \$200540
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32494 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$200540 gate|o|pgate$7
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32495 \$226404 core$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$32496 VDD|pad|pin1|supply|vdd core$4 \$227998 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$32497 \$252776 core$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$32498 VDD|pad|pin1|supply|vdd core$6 \$254718 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$32499 \$278874 core$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$32500 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$317767
+ anode|cathode|pad|pad_RO_101_Drain_Force_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32540 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$317768
+ anode|cathode|pad|pad_RO_101_Drain_Sense_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32580 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$317769
+ anode|cathode|pad|pad_RO_101_extra_load_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32620 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$317770
+ anode|cathode|pad|pad_RO_13_Drain_Force_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32660 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$317771
+ anode|cathode|pad|pad_RO_13_Drain_Sense_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32700 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$317772
+ anode|cathode|pad|pad_RO_13_extra_load_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32740 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$317773
+ ROVDD|VDD|anode|cathode|nclk|pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32780 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$317774
+ RO2VDD|VDD|anode|cathode|nclk|pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$32820 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$8
+ anode|cathode|pad|pad_RO_101_Vout_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$32836 gate|o|pgate$8 \$306590 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32837 \$306590 \$306591 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32838 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$306590 \$306591
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32839 gate|ngate|o$8 \$306593 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32840 \$306593 \$306594 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32841 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$306593 \$306594
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32842 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$9
+ anode|cathode|pad|pad_RO_13_Vout_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$32858 gate|o|pgate$9 \$306596 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32859 \$306596 \$306597 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32860 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$306596 \$306597
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32861 gate|ngate|o$9 \$306599 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$32862 \$306599 \$306600 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$32863 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$306599 \$306600
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$32864 VDD|pad|pin1|supply|vdd core$8 \$280694 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
D$32865 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_rst_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32867 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_clk_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32869 VSS|anode|cathode|clk|vss gate|ngate|o dantenna A=0.6084p P=3.12u m=1
D$32870 VSS|anode|cathode|clk|vss gate|ngate|o$1 dantenna A=0.6084p P=3.12u m=1
D$32871 VSS|anode|cathode|clk|vss gate|ngate|o$2 dantenna A=0.6084p P=3.12u m=1
D$32872 VSS|anode|cathode|clk|vss gate|ngate|o$3 dantenna A=0.6084p P=3.12u m=1
D$32873 VSS|anode|cathode|clk|vss gate|ngate|o$4 dantenna A=0.6084p P=3.12u m=1
D$32874 VSS|anode|cathode|clk|vss gate|ngate|o$5 dantenna A=0.6084p P=3.12u m=1
D$32875 VSS|anode|cathode|clk|vss gate|ngate|o$6 dantenna A=0.6084p P=3.12u m=1
D$32876 VSS|anode|cathode|clk|vss AVDD|anode|cathode|pad|vdd dantenna
+ A=35.0028p P=58.08u m=2
D$32877 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_result_0_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32878 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_result_1_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32879 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_result_2_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32880 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_result_3_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32881 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_result_4_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32882 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_valid_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32883 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_sample_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32885 VSS|anode|cathode|clk|vss core|padres dantenna A=1.984p P=7.48u m=1
D$32886 VSS|anode|cathode|clk|vss core dantenna A=1.984p P=7.48u m=1
D$32887 VSS|anode|cathode|clk|vss core$1 dantenna A=1.984p P=7.48u m=1
D$32895 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_go_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32897 VSS|anode|cathode|clk|vss core$2 dantenna A=1.984p P=7.48u m=1
D$32898 VSS|anode|cathode|clk|vss VSS|anode|cathode|clk|vss dantenna A=35.0028p
+ P=58.08u m=6
D$32902 VSS|anode|cathode|clk|vss VREFH|core|padres dantenna A=1.984p P=7.48u
+ m=1
D$32903 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_vrefp_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32905 VSS|anode|cathode|clk|vss VREFL|core|padres dantenna A=1.984p P=7.48u
+ m=1
D$32906 VSS|anode|cathode|clk|vss gate|out dantenna A=0.2304p P=1.92u m=1
D$32907 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_vrefn_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32909 VSS|anode|cathode|clk|vss VSSIO|anode|cathode|guard|iovss dantenna
+ A=35.0028p P=58.08u m=2
D$32911 VSS|anode|cathode|clk|vss VIN|core|padres dantenna A=1.984p P=7.48u m=1
D$32912 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_vin_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32914 VSS|anode|cathode|clk|vss VIP|core|padres dantenna A=1.984p P=7.48u m=1
D$32915 VSS|anode|cathode|clk|vss gate|out$1 dantenna A=0.2304p P=1.92u m=1
D$32916 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_adc_vip_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32918 VSS|anode|cathode|clk|vss SAMPLE|a1|c2p|core|i|z dantenna A=1.44045p
+ P=4.91u m=2
D$32920 VSS|anode|cathode|clk|vss gate|ngate|o$7 dantenna A=0.6084p P=3.12u m=1
D$32921 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_miso_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32925 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_mosi_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32927 VSS|anode|cathode|clk|vss core$3 dantenna A=1.984p P=7.48u m=1
D$32928 VSS|anode|cathode|clk|vss core$4 dantenna A=1.984p P=7.48u m=1
D$32929 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_RST_B_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32931 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_sclk_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32933 VSS|anode|cathode|clk|vss core$5 dantenna A=1.984p P=7.48u m=1
D$32934 VSS|anode|cathode|clk|vss core$6 dantenna A=1.984p P=7.48u m=1
D$32935 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_101_DUT_gate_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32937 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_cs_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32939 VSS|anode|cathode|clk|vss core$7 dantenna A=1.984p P=7.48u m=1
D$32940 VSS|anode|cathode|clk|vss core$8 dantenna A=1.984p P=7.48u m=1
D$32941 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_13_DUT_gate_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32943 VSS|anode|cathode|clk|vss Drain_Force|Vout|core|padres$1 dantenna
+ A=1.984p P=7.48u m=1
D$32944 VSS|anode|cathode|clk|vss Drain_Sense|Vout|core|padres$1 dantenna
+ A=1.984p P=7.48u m=1
D$32945 VSS|anode|cathode|clk|vss Vin|Vout|core|extra_load|padres$1 dantenna
+ A=1.984p P=7.48u m=1
D$32946 VSS|anode|cathode|clk|vss Drain_Force|Vout|core|padres dantenna
+ A=1.984p P=7.48u m=1
D$32947 VSS|anode|cathode|clk|vss Drain_Sense|Vout|core|padres dantenna
+ A=1.984p P=7.48u m=1
D$32948 VSS|anode|cathode|clk|vss Vin|Vout|core|extra_load|padres dantenna
+ A=1.984p P=7.48u m=1
D$32949 VSS|anode|cathode|clk|vss core|padres$1 dantenna A=1.984p P=7.48u m=1
D$32950 VSS|anode|cathode|clk|vss core|padres$2 dantenna A=1.984p P=7.48u m=1
D$32951 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_101_Drain_Force_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32952 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_101_Drain_Sense_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32953 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_101_extra_load_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32954 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_13_Drain_Force_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32955 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_13_Drain_Sense_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32956 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_13_extra_load_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32957 VSS|anode|cathode|clk|vss ROVDD|VDD|anode|cathode|nclk|pad dantenna
+ A=35.0028p P=58.08u m=2
D$32958 VSS|anode|cathode|clk|vss RO2VDD|VDD|anode|cathode|nclk|pad dantenna
+ A=35.0028p P=58.08u m=2
D$32959 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_101_Vout_pad
+ dantenna A=35.0028p P=58.08u m=2
D$32960 VSS|anode|cathode|clk|vss anode|cathode|pad|pad_RO_13_Vout_pad dantenna
+ A=35.0028p P=58.08u m=2
D$32971 VSS|anode|cathode|clk|vss gate|ngate|o$8 dantenna A=0.6084p P=3.12u m=1
D$32972 VSS|anode|cathode|clk|vss gate|ngate|o$9 dantenna A=0.6084p P=3.12u m=1
D$32973 AVDD|anode|cathode|pad|vdd VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=35.0028p P=58.08u m=2
D$32974 anode|cathode|pad|pad_adc_result_0_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$32975 anode|cathode|pad|pad_adc_result_1_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$32976 anode|cathode|pad|pad_adc_result_2_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$32977 anode|cathode|pad|pad_adc_result_3_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$32978 anode|cathode|pad|pad_adc_result_4_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$32979 anode|cathode|pad|pad_adc_valid_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$32980 anode|cathode|pad|pad_adc_sample_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$32989 anode|cathode|pad|pad_adc_rst_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$32991 anode|cathode|pad|pad_adc_clk_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$32993 gate|o|pgate VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$32994 gate|o|pgate$1 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$32995 gate|o|pgate$2 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$32996 gate|o|pgate$3 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$32997 gate|o|pgate$4 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$32998 gate|o|pgate$5 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$32999 gate|o|pgate$6 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$33000 VSS|anode|cathode|clk|vss VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=35.0028p P=58.08u m=6
D$33002 VREFH|core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$33003 core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$33004 core VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$33005 core$1 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$33006 core$2 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$33007 anode|cathode|pad|pad_adc_go_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33011 anode|cathode|pad|pad_adc_vrefp_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33013 anode|cathode|pad|pad_adc_vrefn_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33015 VREFL|core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$33016 VIN|core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$33017 VSSIO|anode|cathode|guard|iovss
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33019 anode|cathode|pad|pad_adc_vin_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33021 anode|cathode|pad|pad_adc_vip_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33023 VIP|core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$33024 SAMPLE|a1|c2p|core|i|z VDD|pad|pin1|supply|vdd dpantenna A=1.44045p
+ P=4.91u m=2
D$33026 gate|o|pgate$7 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$33027 anode|cathode|pad|pad_miso_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33031 anode|cathode|pad|pad_mosi_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33033 core$3 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$33034 core$4 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$33035 anode|cathode|pad|pad_RO_RST_B_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33037 anode|cathode|pad|pad_sclk_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33039 core$5 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$33040 core$6 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$33041 anode|cathode|pad|pad_RO_101_DUT_gate_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33043 anode|cathode|pad|pad_cs_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=35.0028p P=58.08u m=2
D$33045 core$7 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$33046 core$8 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$33047 anode|cathode|pad|pad_RO_13_DUT_gate_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33049 Drain_Force|Vout|core|padres$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p P=11.24u m=1
D$33050 Drain_Sense|Vout|core|padres$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p P=11.24u m=1
D$33051 Vin|Vout|core|extra_load|padres$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p P=11.24u m=1
D$33052 Drain_Force|Vout|core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=3.1872p P=11.24u m=1
D$33053 Drain_Sense|Vout|core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=3.1872p P=11.24u m=1
D$33054 Vin|Vout|core|extra_load|padres
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p P=11.24u m=1
D$33055 core|padres$1 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$33056 core|padres$2 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$33057 anode|cathode|pad|pad_RO_101_Drain_Force_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33058 anode|cathode|pad|pad_RO_101_Drain_Sense_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33059 anode|cathode|pad|pad_RO_101_extra_load_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33060 anode|cathode|pad|pad_RO_13_Drain_Force_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33061 anode|cathode|pad|pad_RO_13_Drain_Sense_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33062 anode|cathode|pad|pad_RO_13_extra_load_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33063 ROVDD|VDD|anode|cathode|nclk|pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33064 RO2VDD|VDD|anode|cathode|nclk|pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33065 anode|cathode|pad|pad_RO_101_Vout_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33066 gate|o|pgate$8 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$33067 anode|cathode|pad|pad_RO_13_Vout_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$33068 gate|o|pgate$9 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
R$33079 VSSIO|anode|cathode|guard|iovss \$40710 rppd w=0.5u l=3.54u ps=0 b=0 m=1
R$33080 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$50381 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33081 AVDD|anode|cathode|pad|vdd core|padres rppd w=1u l=2u ps=0 b=0 m=1
R$33082 anode|cathode|pad|pad_adc_rst_pad core rppd w=1u l=2u ps=0 b=0 m=1
R$33083 anode|cathode|pad|pad_adc_clk_pad core$1 rppd w=1u l=2u ps=0 b=0 m=1
R$33084 VSSIO|anode|cathode|guard|iovss \$104012 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33085 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$106976 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33086 core$2 anode|cathode|pad|pad_adc_go_pad rppd w=1u l=2u ps=0 b=0 m=1
R$33087 VSSIO|anode|cathode|guard|iovss \$123933 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33088 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$127370 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33089 anode|cathode|pad|pad_adc_vrefp_pad VREFH|core|padres rppd w=1u l=2u
+ ps=0 b=0 m=1
R$33095 anode|cathode|pad|pad_adc_vrefn_pad VREFL|core|padres rppd w=1u l=2u
+ ps=0 b=0 m=1
R$33116 in|pin2 VDD|pad|pin1|supply|vdd rppd w=1u l=520u ps=0 b=0 m=1
R$33117 VSSIO|anode|cathode|guard|iovss \$144244 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33118 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$144245 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33119 VSSIO|anode|cathode|guard|iovss \$165240 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33120 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$168331 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33121 anode|cathode|pad|pad_adc_vin_pad VIN|core|padres rppd w=1u l=2u ps=0
+ b=0 m=1
R$33127 anode|cathode|pad|pad_adc_vip_pad VIP|core|padres rppd w=1u l=2u ps=0
+ b=0 m=1
R$33148 in|pin2$1 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=1u l=520u
+ ps=0 b=0 m=1
R$33149 anode|cathode|pad|pad_RO_RST_B_pad core$3 rppd w=1u l=2u ps=0 b=0 m=1
R$33150 core$4 anode|cathode|pad|pad_mosi_pad rppd w=1u l=2u ps=0 b=0 m=1
R$33151 anode|cathode|pad|pad_RO_101_DUT_gate_pad core$5 rppd w=1u l=2u ps=0
+ b=0 m=1
R$33152 core$6 anode|cathode|pad|pad_sclk_pad rppd w=1u l=2u ps=0 b=0 m=1
R$33153 anode|cathode|pad|pad_RO_13_DUT_gate_pad core$7 rppd w=1u l=2u ps=0 b=0
+ m=1
R$33154 core$8 anode|cathode|pad|pad_cs_pad rppd w=1u l=2u ps=0 b=0 m=1
R$33155 Drain_Force|Vout|core|padres$1
+ anode|cathode|pad|pad_RO_101_Drain_Force_pad rppd w=1u l=2u ps=0 b=0 m=1
R$33156 Drain_Sense|Vout|core|padres$1
+ anode|cathode|pad|pad_RO_101_Drain_Sense_pad rppd w=1u l=2u ps=0 b=0 m=1
R$33157 Vin|Vout|core|extra_load|padres$1
+ anode|cathode|pad|pad_RO_101_extra_load_pad rppd w=1u l=2u ps=0 b=0 m=1
R$33158 Drain_Force|Vout|core|padres
+ anode|cathode|pad|pad_RO_13_Drain_Force_pad rppd w=1u l=2u ps=0 b=0 m=1
R$33159 Drain_Sense|Vout|core|padres
+ anode|cathode|pad|pad_RO_13_Drain_Sense_pad rppd w=1u l=2u ps=0 b=0 m=1
R$33160 Vin|Vout|core|extra_load|padres
+ anode|cathode|pad|pad_RO_13_extra_load_pad rppd w=1u l=2u ps=0 b=0 m=1
R$33161 core|padres$1 ROVDD|VDD|anode|cathode|nclk|pad rppd w=1u l=2u ps=0 b=0
+ m=1
R$33162 core|padres$2 RO2VDD|VDD|anode|cathode|nclk|pad rppd w=1u l=2u ps=0 b=0
+ m=1
R$33163 \$317767 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33164 \$317768 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33165 \$317769 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33166 \$317770 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33167 \$317771 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33168 \$317772 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33169 \$317773 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33170 \$317774 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$33171 \$329246 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33172 \$329247 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33173 \$329248 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33174 \$329249 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33175 \$329250 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33176 \$329251 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33177 \$329252 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$33178 \$329253 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
.ENDS asicone_202508
