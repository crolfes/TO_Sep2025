magic
tech ihp-sg13g2
timestamp 1756304713
<< nwell >>
rect -62 -62 3368 1088
<< pwell >>
rect -179 1145 3485 1205
rect -179 -119 -119 1145
rect 3425 -119 3485 1145
rect -179 -179 3485 -119
<< psubdiff >>
rect -166 1183 3472 1192
rect -166 1167 -157 1183
rect -141 1167 -123 1183
rect -107 1167 -89 1183
rect -73 1167 -55 1183
rect -39 1167 -21 1183
rect -5 1167 13 1183
rect 29 1167 47 1183
rect 63 1167 81 1183
rect 97 1167 115 1183
rect 131 1167 149 1183
rect 165 1167 183 1183
rect 199 1167 217 1183
rect 233 1167 251 1183
rect 267 1167 285 1183
rect 301 1167 319 1183
rect 335 1167 353 1183
rect 369 1167 387 1183
rect 403 1167 421 1183
rect 437 1167 455 1183
rect 471 1167 489 1183
rect 505 1167 523 1183
rect 539 1167 557 1183
rect 573 1167 591 1183
rect 607 1167 625 1183
rect 641 1167 659 1183
rect 675 1167 693 1183
rect 709 1167 727 1183
rect 743 1167 761 1183
rect 777 1167 795 1183
rect 811 1167 829 1183
rect 845 1167 863 1183
rect 879 1167 897 1183
rect 913 1167 931 1183
rect 947 1167 965 1183
rect 981 1167 999 1183
rect 1015 1167 1033 1183
rect 1049 1167 1067 1183
rect 1083 1167 1101 1183
rect 1117 1167 1135 1183
rect 1151 1167 1169 1183
rect 1185 1167 1203 1183
rect 1219 1167 1237 1183
rect 1253 1167 1271 1183
rect 1287 1167 1305 1183
rect 1321 1167 1339 1183
rect 1355 1167 1373 1183
rect 1389 1167 1407 1183
rect 1423 1167 1441 1183
rect 1457 1167 1475 1183
rect 1491 1167 1509 1183
rect 1525 1167 1543 1183
rect 1559 1167 1577 1183
rect 1593 1167 1611 1183
rect 1627 1167 1645 1183
rect 1661 1167 1679 1183
rect 1695 1167 1713 1183
rect 1729 1167 1747 1183
rect 1763 1167 1781 1183
rect 1797 1167 1815 1183
rect 1831 1167 1849 1183
rect 1865 1167 1883 1183
rect 1899 1167 1917 1183
rect 1933 1167 1951 1183
rect 1967 1167 1985 1183
rect 2001 1167 2019 1183
rect 2035 1167 2053 1183
rect 2069 1167 2087 1183
rect 2103 1167 2121 1183
rect 2137 1167 2155 1183
rect 2171 1167 2189 1183
rect 2205 1167 2223 1183
rect 2239 1167 2257 1183
rect 2273 1167 2291 1183
rect 2307 1167 2325 1183
rect 2341 1167 2359 1183
rect 2375 1167 2393 1183
rect 2409 1167 2427 1183
rect 2443 1167 2461 1183
rect 2477 1167 2495 1183
rect 2511 1167 2529 1183
rect 2545 1167 2563 1183
rect 2579 1167 2597 1183
rect 2613 1167 2631 1183
rect 2647 1167 2665 1183
rect 2681 1167 2699 1183
rect 2715 1167 2733 1183
rect 2749 1167 2767 1183
rect 2783 1167 2801 1183
rect 2817 1167 2835 1183
rect 2851 1167 2869 1183
rect 2885 1167 2903 1183
rect 2919 1167 2937 1183
rect 2953 1167 2971 1183
rect 2987 1167 3005 1183
rect 3021 1167 3039 1183
rect 3055 1167 3073 1183
rect 3089 1167 3107 1183
rect 3123 1167 3141 1183
rect 3157 1167 3175 1183
rect 3191 1167 3209 1183
rect 3225 1167 3243 1183
rect 3259 1167 3277 1183
rect 3293 1167 3311 1183
rect 3327 1167 3345 1183
rect 3361 1167 3379 1183
rect 3395 1167 3413 1183
rect 3429 1167 3447 1183
rect 3463 1167 3472 1183
rect -166 1158 3472 1167
rect -166 1133 -132 1158
rect -166 1117 -157 1133
rect -141 1117 -132 1133
rect -166 1099 -132 1117
rect -166 1083 -157 1099
rect -141 1083 -132 1099
rect -166 1065 -132 1083
rect -166 1049 -157 1065
rect -141 1049 -132 1065
rect -166 1031 -132 1049
rect -166 1015 -157 1031
rect -141 1015 -132 1031
rect 3438 1133 3472 1158
rect 3438 1117 3447 1133
rect 3463 1117 3472 1133
rect 3438 1099 3472 1117
rect 3438 1083 3447 1099
rect 3463 1083 3472 1099
rect 3438 1065 3472 1083
rect 3438 1049 3447 1065
rect 3463 1049 3472 1065
rect 3438 1031 3472 1049
rect -166 997 -132 1015
rect -166 981 -157 997
rect -141 981 -132 997
rect -166 963 -132 981
rect -166 947 -157 963
rect -141 947 -132 963
rect -166 929 -132 947
rect -166 913 -157 929
rect -141 913 -132 929
rect -166 895 -132 913
rect -166 879 -157 895
rect -141 879 -132 895
rect -166 861 -132 879
rect -166 845 -157 861
rect -141 845 -132 861
rect -166 827 -132 845
rect -166 811 -157 827
rect -141 811 -132 827
rect -166 793 -132 811
rect -166 777 -157 793
rect -141 777 -132 793
rect -166 759 -132 777
rect -166 743 -157 759
rect -141 743 -132 759
rect -166 725 -132 743
rect -166 709 -157 725
rect -141 709 -132 725
rect -166 691 -132 709
rect -166 675 -157 691
rect -141 675 -132 691
rect -166 657 -132 675
rect -166 641 -157 657
rect -141 641 -132 657
rect -166 623 -132 641
rect -166 607 -157 623
rect -141 607 -132 623
rect -166 589 -132 607
rect -166 573 -157 589
rect -141 573 -132 589
rect -166 555 -132 573
rect -166 539 -157 555
rect -141 539 -132 555
rect -166 521 -132 539
rect -166 505 -157 521
rect -141 505 -132 521
rect -166 487 -132 505
rect -166 471 -157 487
rect -141 471 -132 487
rect -166 453 -132 471
rect -166 437 -157 453
rect -141 437 -132 453
rect -166 419 -132 437
rect -166 403 -157 419
rect -141 403 -132 419
rect -166 385 -132 403
rect -166 369 -157 385
rect -141 369 -132 385
rect -166 351 -132 369
rect -166 335 -157 351
rect -141 335 -132 351
rect -166 317 -132 335
rect -166 301 -157 317
rect -141 301 -132 317
rect -166 283 -132 301
rect -166 267 -157 283
rect -141 267 -132 283
rect -166 249 -132 267
rect -166 233 -157 249
rect -141 233 -132 249
rect -166 215 -132 233
rect -166 199 -157 215
rect -141 199 -132 215
rect -166 181 -132 199
rect -166 165 -157 181
rect -141 165 -132 181
rect -166 147 -132 165
rect -166 131 -157 147
rect -141 131 -132 147
rect -166 113 -132 131
rect -166 97 -157 113
rect -141 97 -132 113
rect -166 79 -132 97
rect -166 63 -157 79
rect -141 63 -132 79
rect -166 45 -132 63
rect -166 29 -157 45
rect -141 29 -132 45
rect -166 11 -132 29
rect -166 -5 -157 11
rect -141 -5 -132 11
rect 3438 1015 3447 1031
rect 3463 1015 3472 1031
rect 3438 997 3472 1015
rect 3438 981 3447 997
rect 3463 981 3472 997
rect 3438 963 3472 981
rect 3438 947 3447 963
rect 3463 947 3472 963
rect 3438 929 3472 947
rect 3438 913 3447 929
rect 3463 913 3472 929
rect 3438 895 3472 913
rect 3438 879 3447 895
rect 3463 879 3472 895
rect 3438 861 3472 879
rect 3438 845 3447 861
rect 3463 845 3472 861
rect 3438 827 3472 845
rect 3438 811 3447 827
rect 3463 811 3472 827
rect 3438 793 3472 811
rect 3438 777 3447 793
rect 3463 777 3472 793
rect 3438 759 3472 777
rect 3438 743 3447 759
rect 3463 743 3472 759
rect 3438 725 3472 743
rect 3438 709 3447 725
rect 3463 709 3472 725
rect 3438 691 3472 709
rect 3438 675 3447 691
rect 3463 675 3472 691
rect 3438 657 3472 675
rect 3438 641 3447 657
rect 3463 641 3472 657
rect 3438 623 3472 641
rect 3438 607 3447 623
rect 3463 607 3472 623
rect 3438 589 3472 607
rect 3438 573 3447 589
rect 3463 573 3472 589
rect 3438 555 3472 573
rect 3438 539 3447 555
rect 3463 539 3472 555
rect 3438 521 3472 539
rect 3438 505 3447 521
rect 3463 505 3472 521
rect 3438 487 3472 505
rect 3438 471 3447 487
rect 3463 471 3472 487
rect 3438 453 3472 471
rect 3438 437 3447 453
rect 3463 437 3472 453
rect 3438 419 3472 437
rect 3438 403 3447 419
rect 3463 403 3472 419
rect 3438 385 3472 403
rect 3438 369 3447 385
rect 3463 369 3472 385
rect 3438 351 3472 369
rect 3438 335 3447 351
rect 3463 335 3472 351
rect 3438 317 3472 335
rect 3438 301 3447 317
rect 3463 301 3472 317
rect 3438 283 3472 301
rect 3438 267 3447 283
rect 3463 267 3472 283
rect 3438 249 3472 267
rect 3438 233 3447 249
rect 3463 233 3472 249
rect 3438 215 3472 233
rect 3438 199 3447 215
rect 3463 199 3472 215
rect 3438 181 3472 199
rect 3438 165 3447 181
rect 3463 165 3472 181
rect 3438 147 3472 165
rect 3438 131 3447 147
rect 3463 131 3472 147
rect 3438 113 3472 131
rect 3438 97 3447 113
rect 3463 97 3472 113
rect 3438 79 3472 97
rect 3438 63 3447 79
rect 3463 63 3472 79
rect 3438 45 3472 63
rect 3438 29 3447 45
rect 3463 29 3472 45
rect 3438 11 3472 29
rect -166 -23 -132 -5
rect -166 -39 -157 -23
rect -141 -39 -132 -23
rect -166 -57 -132 -39
rect -166 -73 -157 -57
rect -141 -73 -132 -57
rect -166 -91 -132 -73
rect -166 -107 -157 -91
rect -141 -107 -132 -91
rect -166 -132 -132 -107
rect 3438 -5 3447 11
rect 3463 -5 3472 11
rect 3438 -23 3472 -5
rect 3438 -39 3447 -23
rect 3463 -39 3472 -23
rect 3438 -57 3472 -39
rect 3438 -73 3447 -57
rect 3463 -73 3472 -57
rect 3438 -91 3472 -73
rect 3438 -107 3447 -91
rect 3463 -107 3472 -91
rect 3438 -132 3472 -107
rect -166 -141 3472 -132
rect -166 -157 -157 -141
rect -141 -157 -123 -141
rect -107 -157 -89 -141
rect -73 -157 -55 -141
rect -39 -157 -21 -141
rect -5 -157 13 -141
rect 29 -157 47 -141
rect 63 -157 81 -141
rect 97 -157 115 -141
rect 131 -157 149 -141
rect 165 -157 183 -141
rect 199 -157 217 -141
rect 233 -157 251 -141
rect 267 -157 285 -141
rect 301 -157 319 -141
rect 335 -157 353 -141
rect 369 -157 387 -141
rect 403 -157 421 -141
rect 437 -157 455 -141
rect 471 -157 489 -141
rect 505 -157 523 -141
rect 539 -157 557 -141
rect 573 -157 591 -141
rect 607 -157 625 -141
rect 641 -157 659 -141
rect 675 -157 693 -141
rect 709 -157 727 -141
rect 743 -157 761 -141
rect 777 -157 795 -141
rect 811 -157 829 -141
rect 845 -157 863 -141
rect 879 -157 897 -141
rect 913 -157 931 -141
rect 947 -157 965 -141
rect 981 -157 999 -141
rect 1015 -157 1033 -141
rect 1049 -157 1067 -141
rect 1083 -157 1101 -141
rect 1117 -157 1135 -141
rect 1151 -157 1169 -141
rect 1185 -157 1203 -141
rect 1219 -157 1237 -141
rect 1253 -157 1271 -141
rect 1287 -157 1305 -141
rect 1321 -157 1339 -141
rect 1355 -157 1373 -141
rect 1389 -157 1407 -141
rect 1423 -157 1441 -141
rect 1457 -157 1475 -141
rect 1491 -157 1509 -141
rect 1525 -157 1543 -141
rect 1559 -157 1577 -141
rect 1593 -157 1611 -141
rect 1627 -157 1645 -141
rect 1661 -157 1679 -141
rect 1695 -157 1713 -141
rect 1729 -157 1747 -141
rect 1763 -157 1781 -141
rect 1797 -157 1815 -141
rect 1831 -157 1849 -141
rect 1865 -157 1883 -141
rect 1899 -157 1917 -141
rect 1933 -157 1951 -141
rect 1967 -157 1985 -141
rect 2001 -157 2019 -141
rect 2035 -157 2053 -141
rect 2069 -157 2087 -141
rect 2103 -157 2121 -141
rect 2137 -157 2155 -141
rect 2171 -157 2189 -141
rect 2205 -157 2223 -141
rect 2239 -157 2257 -141
rect 2273 -157 2291 -141
rect 2307 -157 2325 -141
rect 2341 -157 2359 -141
rect 2375 -157 2393 -141
rect 2409 -157 2427 -141
rect 2443 -157 2461 -141
rect 2477 -157 2495 -141
rect 2511 -157 2529 -141
rect 2545 -157 2563 -141
rect 2579 -157 2597 -141
rect 2613 -157 2631 -141
rect 2647 -157 2665 -141
rect 2681 -157 2699 -141
rect 2715 -157 2733 -141
rect 2749 -157 2767 -141
rect 2783 -157 2801 -141
rect 2817 -157 2835 -141
rect 2851 -157 2869 -141
rect 2885 -157 2903 -141
rect 2919 -157 2937 -141
rect 2953 -157 2971 -141
rect 2987 -157 3005 -141
rect 3021 -157 3039 -141
rect 3055 -157 3073 -141
rect 3089 -157 3107 -141
rect 3123 -157 3141 -141
rect 3157 -157 3175 -141
rect 3191 -157 3209 -141
rect 3225 -157 3243 -141
rect 3259 -157 3277 -141
rect 3293 -157 3311 -141
rect 3327 -157 3345 -141
rect 3361 -157 3379 -141
rect 3395 -157 3413 -141
rect 3429 -157 3447 -141
rect 3463 -157 3472 -141
rect -166 -166 3472 -157
<< nsubdiff >>
rect 0 1014 3306 1026
rect 0 998 21 1014
rect 37 998 55 1014
rect 71 998 89 1014
rect 105 1005 3201 1014
rect 105 998 149 1005
rect 0 989 149 998
rect 165 989 183 1005
rect 199 989 217 1005
rect 233 989 251 1005
rect 267 989 285 1005
rect 301 989 319 1005
rect 335 989 353 1005
rect 369 989 387 1005
rect 403 989 421 1005
rect 437 989 455 1005
rect 471 989 489 1005
rect 505 989 523 1005
rect 539 989 557 1005
rect 573 989 591 1005
rect 607 989 625 1005
rect 641 989 659 1005
rect 675 989 693 1005
rect 709 989 727 1005
rect 743 989 761 1005
rect 777 989 795 1005
rect 811 989 829 1005
rect 845 989 863 1005
rect 879 989 897 1005
rect 913 989 931 1005
rect 947 989 965 1005
rect 981 989 999 1005
rect 1015 989 1033 1005
rect 1049 989 1067 1005
rect 1083 989 1101 1005
rect 1117 989 1135 1005
rect 1151 989 1169 1005
rect 1185 989 1203 1005
rect 1219 989 1237 1005
rect 1253 989 1271 1005
rect 1287 989 1305 1005
rect 1321 989 1339 1005
rect 1355 989 1373 1005
rect 1389 989 1407 1005
rect 1423 989 1441 1005
rect 1457 989 1475 1005
rect 1491 989 1509 1005
rect 1525 989 1543 1005
rect 1559 989 1577 1005
rect 1593 989 1611 1005
rect 1627 989 1645 1005
rect 1661 989 1679 1005
rect 1695 989 1713 1005
rect 1729 989 1747 1005
rect 1763 989 1781 1005
rect 1797 989 1815 1005
rect 1831 989 1849 1005
rect 1865 989 1883 1005
rect 1899 989 1917 1005
rect 1933 989 1951 1005
rect 1967 989 1985 1005
rect 2001 989 2019 1005
rect 2035 989 2053 1005
rect 2069 989 2087 1005
rect 2103 989 2121 1005
rect 2137 989 2155 1005
rect 2171 989 2189 1005
rect 2205 989 2223 1005
rect 2239 989 2257 1005
rect 2273 989 2291 1005
rect 2307 989 2325 1005
rect 2341 989 2359 1005
rect 2375 989 2393 1005
rect 2409 989 2427 1005
rect 2443 989 2461 1005
rect 2477 989 2495 1005
rect 2511 989 2529 1005
rect 2545 989 2563 1005
rect 2579 989 2597 1005
rect 2613 989 2631 1005
rect 2647 989 2665 1005
rect 2681 989 2699 1005
rect 2715 989 2733 1005
rect 2749 989 2767 1005
rect 2783 989 2801 1005
rect 2817 989 2835 1005
rect 2851 989 2869 1005
rect 2885 989 2903 1005
rect 2919 989 2937 1005
rect 2953 989 2971 1005
rect 2987 989 3005 1005
rect 3021 989 3039 1005
rect 3055 989 3073 1005
rect 3089 989 3107 1005
rect 3123 989 3141 1005
rect 3157 998 3201 1005
rect 3217 998 3235 1014
rect 3251 998 3269 1014
rect 3285 998 3306 1014
rect 3157 989 3306 998
rect 0 980 3306 989
rect 0 964 21 980
rect 37 964 55 980
rect 71 964 89 980
rect 105 971 3201 980
rect 105 964 149 971
rect 0 955 149 964
rect 165 955 183 971
rect 199 955 217 971
rect 233 955 251 971
rect 267 955 285 971
rect 301 955 319 971
rect 335 955 353 971
rect 369 955 387 971
rect 403 955 421 971
rect 437 955 455 971
rect 471 955 489 971
rect 505 955 523 971
rect 539 955 557 971
rect 573 955 591 971
rect 607 955 625 971
rect 641 955 659 971
rect 675 955 693 971
rect 709 955 727 971
rect 743 955 761 971
rect 777 955 795 971
rect 811 955 829 971
rect 845 955 863 971
rect 879 955 897 971
rect 913 955 931 971
rect 947 955 965 971
rect 981 955 999 971
rect 1015 955 1033 971
rect 1049 955 1067 971
rect 1083 955 1101 971
rect 1117 955 1135 971
rect 1151 955 1169 971
rect 1185 955 1203 971
rect 1219 955 1237 971
rect 1253 955 1271 971
rect 1287 955 1305 971
rect 1321 955 1339 971
rect 1355 955 1373 971
rect 1389 955 1407 971
rect 1423 955 1441 971
rect 1457 955 1475 971
rect 1491 955 1509 971
rect 1525 955 1543 971
rect 1559 955 1577 971
rect 1593 955 1611 971
rect 1627 955 1645 971
rect 1661 955 1679 971
rect 1695 955 1713 971
rect 1729 955 1747 971
rect 1763 955 1781 971
rect 1797 955 1815 971
rect 1831 955 1849 971
rect 1865 955 1883 971
rect 1899 955 1917 971
rect 1933 955 1951 971
rect 1967 955 1985 971
rect 2001 955 2019 971
rect 2035 955 2053 971
rect 2069 955 2087 971
rect 2103 955 2121 971
rect 2137 955 2155 971
rect 2171 955 2189 971
rect 2205 955 2223 971
rect 2239 955 2257 971
rect 2273 955 2291 971
rect 2307 955 2325 971
rect 2341 955 2359 971
rect 2375 955 2393 971
rect 2409 955 2427 971
rect 2443 955 2461 971
rect 2477 955 2495 971
rect 2511 955 2529 971
rect 2545 955 2563 971
rect 2579 955 2597 971
rect 2613 955 2631 971
rect 2647 955 2665 971
rect 2681 955 2699 971
rect 2715 955 2733 971
rect 2749 955 2767 971
rect 2783 955 2801 971
rect 2817 955 2835 971
rect 2851 955 2869 971
rect 2885 955 2903 971
rect 2919 955 2937 971
rect 2953 955 2971 971
rect 2987 955 3005 971
rect 3021 955 3039 971
rect 3055 955 3073 971
rect 3089 955 3107 971
rect 3123 955 3141 971
rect 3157 964 3201 971
rect 3217 964 3235 980
rect 3251 964 3269 980
rect 3285 964 3306 980
rect 3157 955 3306 964
rect 0 946 3306 955
rect 0 930 21 946
rect 37 930 55 946
rect 71 930 89 946
rect 105 937 3201 946
rect 105 930 149 937
rect 0 921 149 930
rect 165 921 183 937
rect 199 921 217 937
rect 233 921 251 937
rect 267 921 285 937
rect 301 921 319 937
rect 335 921 353 937
rect 369 921 387 937
rect 403 921 421 937
rect 437 921 455 937
rect 471 921 489 937
rect 505 921 523 937
rect 539 921 557 937
rect 573 921 591 937
rect 607 921 625 937
rect 641 921 659 937
rect 675 921 693 937
rect 709 921 727 937
rect 743 921 761 937
rect 777 921 795 937
rect 811 921 829 937
rect 845 921 863 937
rect 879 921 897 937
rect 913 921 931 937
rect 947 921 965 937
rect 981 921 999 937
rect 1015 921 1033 937
rect 1049 921 1067 937
rect 1083 921 1101 937
rect 1117 921 1135 937
rect 1151 921 1169 937
rect 1185 921 1203 937
rect 1219 921 1237 937
rect 1253 921 1271 937
rect 1287 921 1305 937
rect 1321 921 1339 937
rect 1355 921 1373 937
rect 1389 921 1407 937
rect 1423 921 1441 937
rect 1457 921 1475 937
rect 1491 921 1509 937
rect 1525 921 1543 937
rect 1559 921 1577 937
rect 1593 921 1611 937
rect 1627 921 1645 937
rect 1661 921 1679 937
rect 1695 921 1713 937
rect 1729 921 1747 937
rect 1763 921 1781 937
rect 1797 921 1815 937
rect 1831 921 1849 937
rect 1865 921 1883 937
rect 1899 921 1917 937
rect 1933 921 1951 937
rect 1967 921 1985 937
rect 2001 921 2019 937
rect 2035 921 2053 937
rect 2069 921 2087 937
rect 2103 921 2121 937
rect 2137 921 2155 937
rect 2171 921 2189 937
rect 2205 921 2223 937
rect 2239 921 2257 937
rect 2273 921 2291 937
rect 2307 921 2325 937
rect 2341 921 2359 937
rect 2375 921 2393 937
rect 2409 921 2427 937
rect 2443 921 2461 937
rect 2477 921 2495 937
rect 2511 921 2529 937
rect 2545 921 2563 937
rect 2579 921 2597 937
rect 2613 921 2631 937
rect 2647 921 2665 937
rect 2681 921 2699 937
rect 2715 921 2733 937
rect 2749 921 2767 937
rect 2783 921 2801 937
rect 2817 921 2835 937
rect 2851 921 2869 937
rect 2885 921 2903 937
rect 2919 921 2937 937
rect 2953 921 2971 937
rect 2987 921 3005 937
rect 3021 921 3039 937
rect 3055 921 3073 937
rect 3089 921 3107 937
rect 3123 921 3141 937
rect 3157 930 3201 937
rect 3217 930 3235 946
rect 3251 930 3269 946
rect 3285 930 3306 946
rect 3157 921 3306 930
rect 0 912 3306 921
rect 0 896 21 912
rect 37 896 55 912
rect 71 896 89 912
rect 105 900 3201 912
rect 105 896 126 900
rect 0 878 126 896
rect 0 862 21 878
rect 37 862 55 878
rect 71 862 89 878
rect 105 862 126 878
rect 0 844 126 862
rect 0 828 21 844
rect 37 828 55 844
rect 71 828 89 844
rect 105 828 126 844
rect 0 810 126 828
rect 0 794 21 810
rect 37 794 55 810
rect 71 794 89 810
rect 105 794 126 810
rect 3180 896 3201 900
rect 3217 896 3235 912
rect 3251 896 3269 912
rect 3285 896 3306 912
rect 3180 878 3306 896
rect 3180 862 3201 878
rect 3217 862 3235 878
rect 3251 862 3269 878
rect 3285 862 3306 878
rect 3180 844 3306 862
rect 3180 828 3201 844
rect 3217 828 3235 844
rect 3251 828 3269 844
rect 3285 828 3306 844
rect 3180 810 3306 828
rect 0 776 126 794
rect 0 760 21 776
rect 37 760 55 776
rect 71 760 89 776
rect 105 760 126 776
rect 0 742 126 760
rect 0 726 21 742
rect 37 726 55 742
rect 71 726 89 742
rect 105 726 126 742
rect 0 708 126 726
rect 0 692 21 708
rect 37 692 55 708
rect 71 692 89 708
rect 105 692 126 708
rect 0 674 126 692
rect 3180 794 3201 810
rect 3217 794 3235 810
rect 3251 794 3269 810
rect 3285 794 3306 810
rect 3180 776 3306 794
rect 3180 760 3201 776
rect 3217 760 3235 776
rect 3251 760 3269 776
rect 3285 760 3306 776
rect 3180 742 3306 760
rect 3180 726 3201 742
rect 3217 726 3235 742
rect 3251 726 3269 742
rect 3285 726 3306 742
rect 3180 708 3306 726
rect 3180 692 3201 708
rect 3217 692 3235 708
rect 3251 692 3269 708
rect 3285 692 3306 708
rect 0 658 21 674
rect 37 658 55 674
rect 71 658 89 674
rect 105 658 126 674
rect 0 640 126 658
rect 0 624 21 640
rect 37 624 55 640
rect 71 624 89 640
rect 105 624 126 640
rect 0 606 126 624
rect 0 590 21 606
rect 37 590 55 606
rect 71 590 89 606
rect 105 590 126 606
rect 0 576 126 590
rect 3180 674 3306 692
rect 3180 658 3201 674
rect 3217 658 3235 674
rect 3251 658 3269 674
rect 3285 658 3306 674
rect 3180 640 3306 658
rect 3180 624 3201 640
rect 3217 624 3235 640
rect 3251 624 3269 640
rect 3285 624 3306 640
rect 3180 606 3306 624
rect 3180 590 3201 606
rect 3217 590 3235 606
rect 3251 590 3269 606
rect 3285 590 3306 606
rect 3180 576 3306 590
rect 0 572 3306 576
rect 0 556 21 572
rect 37 556 55 572
rect 71 556 89 572
rect 105 556 3201 572
rect 3217 556 3235 572
rect 3251 556 3269 572
rect 3285 556 3306 572
rect 0 555 3306 556
rect 0 539 149 555
rect 165 539 183 555
rect 199 539 217 555
rect 233 539 251 555
rect 267 539 285 555
rect 301 539 319 555
rect 335 539 353 555
rect 369 539 387 555
rect 403 539 421 555
rect 437 539 455 555
rect 471 539 489 555
rect 505 539 523 555
rect 539 539 557 555
rect 573 539 591 555
rect 607 539 625 555
rect 641 539 659 555
rect 675 539 693 555
rect 709 539 727 555
rect 743 539 761 555
rect 777 539 795 555
rect 811 539 829 555
rect 845 539 863 555
rect 879 539 897 555
rect 913 539 931 555
rect 947 539 965 555
rect 981 539 999 555
rect 1015 539 1033 555
rect 1049 539 1067 555
rect 1083 539 1101 555
rect 1117 539 1135 555
rect 1151 539 1169 555
rect 1185 539 1203 555
rect 1219 539 1237 555
rect 1253 539 1271 555
rect 1287 539 1305 555
rect 1321 539 1339 555
rect 1355 539 1373 555
rect 1389 539 1407 555
rect 1423 539 1441 555
rect 1457 539 1475 555
rect 1491 539 1509 555
rect 1525 539 1543 555
rect 1559 539 1577 555
rect 1593 539 1611 555
rect 1627 539 1645 555
rect 1661 539 1679 555
rect 1695 539 1713 555
rect 1729 539 1747 555
rect 1763 539 1781 555
rect 1797 539 1815 555
rect 1831 539 1849 555
rect 1865 539 1883 555
rect 1899 539 1917 555
rect 1933 539 1951 555
rect 1967 539 1985 555
rect 2001 539 2019 555
rect 2035 539 2053 555
rect 2069 539 2087 555
rect 2103 539 2121 555
rect 2137 539 2155 555
rect 2171 539 2189 555
rect 2205 539 2223 555
rect 2239 539 2257 555
rect 2273 539 2291 555
rect 2307 539 2325 555
rect 2341 539 2359 555
rect 2375 539 2393 555
rect 2409 539 2427 555
rect 2443 539 2461 555
rect 2477 539 2495 555
rect 2511 539 2529 555
rect 2545 539 2563 555
rect 2579 539 2597 555
rect 2613 539 2631 555
rect 2647 539 2665 555
rect 2681 539 2699 555
rect 2715 539 2733 555
rect 2749 539 2767 555
rect 2783 539 2801 555
rect 2817 539 2835 555
rect 2851 539 2869 555
rect 2885 539 2903 555
rect 2919 539 2937 555
rect 2953 539 2971 555
rect 2987 539 3005 555
rect 3021 539 3039 555
rect 3055 539 3073 555
rect 3089 539 3107 555
rect 3123 539 3141 555
rect 3157 539 3306 555
rect 0 538 3306 539
rect 0 522 21 538
rect 37 522 55 538
rect 71 522 89 538
rect 105 522 3201 538
rect 3217 522 3235 538
rect 3251 522 3269 538
rect 3285 522 3306 538
rect 0 521 3306 522
rect 0 505 149 521
rect 165 505 183 521
rect 199 505 217 521
rect 233 505 251 521
rect 267 505 285 521
rect 301 505 319 521
rect 335 505 353 521
rect 369 505 387 521
rect 403 505 421 521
rect 437 505 455 521
rect 471 505 489 521
rect 505 505 523 521
rect 539 505 557 521
rect 573 505 591 521
rect 607 505 625 521
rect 641 505 659 521
rect 675 505 693 521
rect 709 505 727 521
rect 743 505 761 521
rect 777 505 795 521
rect 811 505 829 521
rect 845 505 863 521
rect 879 505 897 521
rect 913 505 931 521
rect 947 505 965 521
rect 981 505 999 521
rect 1015 505 1033 521
rect 1049 505 1067 521
rect 1083 505 1101 521
rect 1117 505 1135 521
rect 1151 505 1169 521
rect 1185 505 1203 521
rect 1219 505 1237 521
rect 1253 505 1271 521
rect 1287 505 1305 521
rect 1321 505 1339 521
rect 1355 505 1373 521
rect 1389 505 1407 521
rect 1423 505 1441 521
rect 1457 505 1475 521
rect 1491 505 1509 521
rect 1525 505 1543 521
rect 1559 505 1577 521
rect 1593 505 1611 521
rect 1627 505 1645 521
rect 1661 505 1679 521
rect 1695 505 1713 521
rect 1729 505 1747 521
rect 1763 505 1781 521
rect 1797 505 1815 521
rect 1831 505 1849 521
rect 1865 505 1883 521
rect 1899 505 1917 521
rect 1933 505 1951 521
rect 1967 505 1985 521
rect 2001 505 2019 521
rect 2035 505 2053 521
rect 2069 505 2087 521
rect 2103 505 2121 521
rect 2137 505 2155 521
rect 2171 505 2189 521
rect 2205 505 2223 521
rect 2239 505 2257 521
rect 2273 505 2291 521
rect 2307 505 2325 521
rect 2341 505 2359 521
rect 2375 505 2393 521
rect 2409 505 2427 521
rect 2443 505 2461 521
rect 2477 505 2495 521
rect 2511 505 2529 521
rect 2545 505 2563 521
rect 2579 505 2597 521
rect 2613 505 2631 521
rect 2647 505 2665 521
rect 2681 505 2699 521
rect 2715 505 2733 521
rect 2749 505 2767 521
rect 2783 505 2801 521
rect 2817 505 2835 521
rect 2851 505 2869 521
rect 2885 505 2903 521
rect 2919 505 2937 521
rect 2953 505 2971 521
rect 2987 505 3005 521
rect 3021 505 3039 521
rect 3055 505 3073 521
rect 3089 505 3107 521
rect 3123 505 3141 521
rect 3157 505 3306 521
rect 0 504 3306 505
rect 0 488 21 504
rect 37 488 55 504
rect 71 488 89 504
rect 105 488 3201 504
rect 3217 488 3235 504
rect 3251 488 3269 504
rect 3285 488 3306 504
rect 0 487 3306 488
rect 0 471 149 487
rect 165 471 183 487
rect 199 471 217 487
rect 233 471 251 487
rect 267 471 285 487
rect 301 471 319 487
rect 335 471 353 487
rect 369 471 387 487
rect 403 471 421 487
rect 437 471 455 487
rect 471 471 489 487
rect 505 471 523 487
rect 539 471 557 487
rect 573 471 591 487
rect 607 471 625 487
rect 641 471 659 487
rect 675 471 693 487
rect 709 471 727 487
rect 743 471 761 487
rect 777 471 795 487
rect 811 471 829 487
rect 845 471 863 487
rect 879 471 897 487
rect 913 471 931 487
rect 947 471 965 487
rect 981 471 999 487
rect 1015 471 1033 487
rect 1049 471 1067 487
rect 1083 471 1101 487
rect 1117 471 1135 487
rect 1151 471 1169 487
rect 1185 471 1203 487
rect 1219 471 1237 487
rect 1253 471 1271 487
rect 1287 471 1305 487
rect 1321 471 1339 487
rect 1355 471 1373 487
rect 1389 471 1407 487
rect 1423 471 1441 487
rect 1457 471 1475 487
rect 1491 471 1509 487
rect 1525 471 1543 487
rect 1559 471 1577 487
rect 1593 471 1611 487
rect 1627 471 1645 487
rect 1661 471 1679 487
rect 1695 471 1713 487
rect 1729 471 1747 487
rect 1763 471 1781 487
rect 1797 471 1815 487
rect 1831 471 1849 487
rect 1865 471 1883 487
rect 1899 471 1917 487
rect 1933 471 1951 487
rect 1967 471 1985 487
rect 2001 471 2019 487
rect 2035 471 2053 487
rect 2069 471 2087 487
rect 2103 471 2121 487
rect 2137 471 2155 487
rect 2171 471 2189 487
rect 2205 471 2223 487
rect 2239 471 2257 487
rect 2273 471 2291 487
rect 2307 471 2325 487
rect 2341 471 2359 487
rect 2375 471 2393 487
rect 2409 471 2427 487
rect 2443 471 2461 487
rect 2477 471 2495 487
rect 2511 471 2529 487
rect 2545 471 2563 487
rect 2579 471 2597 487
rect 2613 471 2631 487
rect 2647 471 2665 487
rect 2681 471 2699 487
rect 2715 471 2733 487
rect 2749 471 2767 487
rect 2783 471 2801 487
rect 2817 471 2835 487
rect 2851 471 2869 487
rect 2885 471 2903 487
rect 2919 471 2937 487
rect 2953 471 2971 487
rect 2987 471 3005 487
rect 3021 471 3039 487
rect 3055 471 3073 487
rect 3089 471 3107 487
rect 3123 471 3141 487
rect 3157 471 3306 487
rect 0 470 3306 471
rect 0 454 21 470
rect 37 454 55 470
rect 71 454 89 470
rect 105 454 3201 470
rect 3217 454 3235 470
rect 3251 454 3269 470
rect 3285 454 3306 470
rect 0 450 3306 454
rect 0 436 126 450
rect 0 420 21 436
rect 37 420 55 436
rect 71 420 89 436
rect 105 420 126 436
rect 0 402 126 420
rect 0 386 21 402
rect 37 386 55 402
rect 71 386 89 402
rect 105 386 126 402
rect 0 368 126 386
rect 0 352 21 368
rect 37 352 55 368
rect 71 352 89 368
rect 105 352 126 368
rect 0 334 126 352
rect 3180 436 3306 450
rect 3180 420 3201 436
rect 3217 420 3235 436
rect 3251 420 3269 436
rect 3285 420 3306 436
rect 3180 402 3306 420
rect 3180 386 3201 402
rect 3217 386 3235 402
rect 3251 386 3269 402
rect 3285 386 3306 402
rect 3180 368 3306 386
rect 3180 352 3201 368
rect 3217 352 3235 368
rect 3251 352 3269 368
rect 3285 352 3306 368
rect 0 318 21 334
rect 37 318 55 334
rect 71 318 89 334
rect 105 318 126 334
rect 0 300 126 318
rect 0 284 21 300
rect 37 284 55 300
rect 71 284 89 300
rect 105 284 126 300
rect 0 266 126 284
rect 0 250 21 266
rect 37 250 55 266
rect 71 250 89 266
rect 105 250 126 266
rect 0 232 126 250
rect 0 216 21 232
rect 37 216 55 232
rect 71 216 89 232
rect 105 216 126 232
rect 3180 334 3306 352
rect 3180 318 3201 334
rect 3217 318 3235 334
rect 3251 318 3269 334
rect 3285 318 3306 334
rect 3180 300 3306 318
rect 3180 284 3201 300
rect 3217 284 3235 300
rect 3251 284 3269 300
rect 3285 284 3306 300
rect 3180 266 3306 284
rect 3180 250 3201 266
rect 3217 250 3235 266
rect 3251 250 3269 266
rect 3285 250 3306 266
rect 3180 232 3306 250
rect 0 198 126 216
rect 0 182 21 198
rect 37 182 55 198
rect 71 182 89 198
rect 105 182 126 198
rect 0 164 126 182
rect 0 148 21 164
rect 37 148 55 164
rect 71 148 89 164
rect 105 148 126 164
rect 0 130 126 148
rect 0 114 21 130
rect 37 114 55 130
rect 71 114 89 130
rect 105 126 126 130
rect 3180 216 3201 232
rect 3217 216 3235 232
rect 3251 216 3269 232
rect 3285 216 3306 232
rect 3180 198 3306 216
rect 3180 182 3201 198
rect 3217 182 3235 198
rect 3251 182 3269 198
rect 3285 182 3306 198
rect 3180 164 3306 182
rect 3180 148 3201 164
rect 3217 148 3235 164
rect 3251 148 3269 164
rect 3285 148 3306 164
rect 3180 130 3306 148
rect 3180 126 3201 130
rect 105 114 3201 126
rect 3217 114 3235 130
rect 3251 114 3269 130
rect 3285 114 3306 130
rect 0 105 3306 114
rect 0 96 149 105
rect 0 80 21 96
rect 37 80 55 96
rect 71 80 89 96
rect 105 89 149 96
rect 165 89 183 105
rect 199 89 217 105
rect 233 89 251 105
rect 267 89 285 105
rect 301 89 319 105
rect 335 89 353 105
rect 369 89 387 105
rect 403 89 421 105
rect 437 89 455 105
rect 471 89 489 105
rect 505 89 523 105
rect 539 89 557 105
rect 573 89 591 105
rect 607 89 625 105
rect 641 89 659 105
rect 675 89 693 105
rect 709 89 727 105
rect 743 89 761 105
rect 777 89 795 105
rect 811 89 829 105
rect 845 89 863 105
rect 879 89 897 105
rect 913 89 931 105
rect 947 89 965 105
rect 981 89 999 105
rect 1015 89 1033 105
rect 1049 89 1067 105
rect 1083 89 1101 105
rect 1117 89 1135 105
rect 1151 89 1169 105
rect 1185 89 1203 105
rect 1219 89 1237 105
rect 1253 89 1271 105
rect 1287 89 1305 105
rect 1321 89 1339 105
rect 1355 89 1373 105
rect 1389 89 1407 105
rect 1423 89 1441 105
rect 1457 89 1475 105
rect 1491 89 1509 105
rect 1525 89 1543 105
rect 1559 89 1577 105
rect 1593 89 1611 105
rect 1627 89 1645 105
rect 1661 89 1679 105
rect 1695 89 1713 105
rect 1729 89 1747 105
rect 1763 89 1781 105
rect 1797 89 1815 105
rect 1831 89 1849 105
rect 1865 89 1883 105
rect 1899 89 1917 105
rect 1933 89 1951 105
rect 1967 89 1985 105
rect 2001 89 2019 105
rect 2035 89 2053 105
rect 2069 89 2087 105
rect 2103 89 2121 105
rect 2137 89 2155 105
rect 2171 89 2189 105
rect 2205 89 2223 105
rect 2239 89 2257 105
rect 2273 89 2291 105
rect 2307 89 2325 105
rect 2341 89 2359 105
rect 2375 89 2393 105
rect 2409 89 2427 105
rect 2443 89 2461 105
rect 2477 89 2495 105
rect 2511 89 2529 105
rect 2545 89 2563 105
rect 2579 89 2597 105
rect 2613 89 2631 105
rect 2647 89 2665 105
rect 2681 89 2699 105
rect 2715 89 2733 105
rect 2749 89 2767 105
rect 2783 89 2801 105
rect 2817 89 2835 105
rect 2851 89 2869 105
rect 2885 89 2903 105
rect 2919 89 2937 105
rect 2953 89 2971 105
rect 2987 89 3005 105
rect 3021 89 3039 105
rect 3055 89 3073 105
rect 3089 89 3107 105
rect 3123 89 3141 105
rect 3157 96 3306 105
rect 3157 89 3201 96
rect 105 80 3201 89
rect 3217 80 3235 96
rect 3251 80 3269 96
rect 3285 80 3306 96
rect 0 71 3306 80
rect 0 62 149 71
rect 0 46 21 62
rect 37 46 55 62
rect 71 46 89 62
rect 105 55 149 62
rect 165 55 183 71
rect 199 55 217 71
rect 233 55 251 71
rect 267 55 285 71
rect 301 55 319 71
rect 335 55 353 71
rect 369 55 387 71
rect 403 55 421 71
rect 437 55 455 71
rect 471 55 489 71
rect 505 55 523 71
rect 539 55 557 71
rect 573 55 591 71
rect 607 55 625 71
rect 641 55 659 71
rect 675 55 693 71
rect 709 55 727 71
rect 743 55 761 71
rect 777 55 795 71
rect 811 55 829 71
rect 845 55 863 71
rect 879 55 897 71
rect 913 55 931 71
rect 947 55 965 71
rect 981 55 999 71
rect 1015 55 1033 71
rect 1049 55 1067 71
rect 1083 55 1101 71
rect 1117 55 1135 71
rect 1151 55 1169 71
rect 1185 55 1203 71
rect 1219 55 1237 71
rect 1253 55 1271 71
rect 1287 55 1305 71
rect 1321 55 1339 71
rect 1355 55 1373 71
rect 1389 55 1407 71
rect 1423 55 1441 71
rect 1457 55 1475 71
rect 1491 55 1509 71
rect 1525 55 1543 71
rect 1559 55 1577 71
rect 1593 55 1611 71
rect 1627 55 1645 71
rect 1661 55 1679 71
rect 1695 55 1713 71
rect 1729 55 1747 71
rect 1763 55 1781 71
rect 1797 55 1815 71
rect 1831 55 1849 71
rect 1865 55 1883 71
rect 1899 55 1917 71
rect 1933 55 1951 71
rect 1967 55 1985 71
rect 2001 55 2019 71
rect 2035 55 2053 71
rect 2069 55 2087 71
rect 2103 55 2121 71
rect 2137 55 2155 71
rect 2171 55 2189 71
rect 2205 55 2223 71
rect 2239 55 2257 71
rect 2273 55 2291 71
rect 2307 55 2325 71
rect 2341 55 2359 71
rect 2375 55 2393 71
rect 2409 55 2427 71
rect 2443 55 2461 71
rect 2477 55 2495 71
rect 2511 55 2529 71
rect 2545 55 2563 71
rect 2579 55 2597 71
rect 2613 55 2631 71
rect 2647 55 2665 71
rect 2681 55 2699 71
rect 2715 55 2733 71
rect 2749 55 2767 71
rect 2783 55 2801 71
rect 2817 55 2835 71
rect 2851 55 2869 71
rect 2885 55 2903 71
rect 2919 55 2937 71
rect 2953 55 2971 71
rect 2987 55 3005 71
rect 3021 55 3039 71
rect 3055 55 3073 71
rect 3089 55 3107 71
rect 3123 55 3141 71
rect 3157 62 3306 71
rect 3157 55 3201 62
rect 105 46 3201 55
rect 3217 46 3235 62
rect 3251 46 3269 62
rect 3285 46 3306 62
rect 0 37 3306 46
rect 0 28 149 37
rect 0 12 21 28
rect 37 12 55 28
rect 71 12 89 28
rect 105 21 149 28
rect 165 21 183 37
rect 199 21 217 37
rect 233 21 251 37
rect 267 21 285 37
rect 301 21 319 37
rect 335 21 353 37
rect 369 21 387 37
rect 403 21 421 37
rect 437 21 455 37
rect 471 21 489 37
rect 505 21 523 37
rect 539 21 557 37
rect 573 21 591 37
rect 607 21 625 37
rect 641 21 659 37
rect 675 21 693 37
rect 709 21 727 37
rect 743 21 761 37
rect 777 21 795 37
rect 811 21 829 37
rect 845 21 863 37
rect 879 21 897 37
rect 913 21 931 37
rect 947 21 965 37
rect 981 21 999 37
rect 1015 21 1033 37
rect 1049 21 1067 37
rect 1083 21 1101 37
rect 1117 21 1135 37
rect 1151 21 1169 37
rect 1185 21 1203 37
rect 1219 21 1237 37
rect 1253 21 1271 37
rect 1287 21 1305 37
rect 1321 21 1339 37
rect 1355 21 1373 37
rect 1389 21 1407 37
rect 1423 21 1441 37
rect 1457 21 1475 37
rect 1491 21 1509 37
rect 1525 21 1543 37
rect 1559 21 1577 37
rect 1593 21 1611 37
rect 1627 21 1645 37
rect 1661 21 1679 37
rect 1695 21 1713 37
rect 1729 21 1747 37
rect 1763 21 1781 37
rect 1797 21 1815 37
rect 1831 21 1849 37
rect 1865 21 1883 37
rect 1899 21 1917 37
rect 1933 21 1951 37
rect 1967 21 1985 37
rect 2001 21 2019 37
rect 2035 21 2053 37
rect 2069 21 2087 37
rect 2103 21 2121 37
rect 2137 21 2155 37
rect 2171 21 2189 37
rect 2205 21 2223 37
rect 2239 21 2257 37
rect 2273 21 2291 37
rect 2307 21 2325 37
rect 2341 21 2359 37
rect 2375 21 2393 37
rect 2409 21 2427 37
rect 2443 21 2461 37
rect 2477 21 2495 37
rect 2511 21 2529 37
rect 2545 21 2563 37
rect 2579 21 2597 37
rect 2613 21 2631 37
rect 2647 21 2665 37
rect 2681 21 2699 37
rect 2715 21 2733 37
rect 2749 21 2767 37
rect 2783 21 2801 37
rect 2817 21 2835 37
rect 2851 21 2869 37
rect 2885 21 2903 37
rect 2919 21 2937 37
rect 2953 21 2971 37
rect 2987 21 3005 37
rect 3021 21 3039 37
rect 3055 21 3073 37
rect 3089 21 3107 37
rect 3123 21 3141 37
rect 3157 28 3306 37
rect 3157 21 3201 28
rect 105 12 3201 21
rect 3217 12 3235 28
rect 3251 12 3269 28
rect 3285 12 3306 28
rect 0 0 3306 12
<< psubdiffcont >>
rect -157 1167 -141 1183
rect -123 1167 -107 1183
rect -89 1167 -73 1183
rect -55 1167 -39 1183
rect -21 1167 -5 1183
rect 13 1167 29 1183
rect 47 1167 63 1183
rect 81 1167 97 1183
rect 115 1167 131 1183
rect 149 1167 165 1183
rect 183 1167 199 1183
rect 217 1167 233 1183
rect 251 1167 267 1183
rect 285 1167 301 1183
rect 319 1167 335 1183
rect 353 1167 369 1183
rect 387 1167 403 1183
rect 421 1167 437 1183
rect 455 1167 471 1183
rect 489 1167 505 1183
rect 523 1167 539 1183
rect 557 1167 573 1183
rect 591 1167 607 1183
rect 625 1167 641 1183
rect 659 1167 675 1183
rect 693 1167 709 1183
rect 727 1167 743 1183
rect 761 1167 777 1183
rect 795 1167 811 1183
rect 829 1167 845 1183
rect 863 1167 879 1183
rect 897 1167 913 1183
rect 931 1167 947 1183
rect 965 1167 981 1183
rect 999 1167 1015 1183
rect 1033 1167 1049 1183
rect 1067 1167 1083 1183
rect 1101 1167 1117 1183
rect 1135 1167 1151 1183
rect 1169 1167 1185 1183
rect 1203 1167 1219 1183
rect 1237 1167 1253 1183
rect 1271 1167 1287 1183
rect 1305 1167 1321 1183
rect 1339 1167 1355 1183
rect 1373 1167 1389 1183
rect 1407 1167 1423 1183
rect 1441 1167 1457 1183
rect 1475 1167 1491 1183
rect 1509 1167 1525 1183
rect 1543 1167 1559 1183
rect 1577 1167 1593 1183
rect 1611 1167 1627 1183
rect 1645 1167 1661 1183
rect 1679 1167 1695 1183
rect 1713 1167 1729 1183
rect 1747 1167 1763 1183
rect 1781 1167 1797 1183
rect 1815 1167 1831 1183
rect 1849 1167 1865 1183
rect 1883 1167 1899 1183
rect 1917 1167 1933 1183
rect 1951 1167 1967 1183
rect 1985 1167 2001 1183
rect 2019 1167 2035 1183
rect 2053 1167 2069 1183
rect 2087 1167 2103 1183
rect 2121 1167 2137 1183
rect 2155 1167 2171 1183
rect 2189 1167 2205 1183
rect 2223 1167 2239 1183
rect 2257 1167 2273 1183
rect 2291 1167 2307 1183
rect 2325 1167 2341 1183
rect 2359 1167 2375 1183
rect 2393 1167 2409 1183
rect 2427 1167 2443 1183
rect 2461 1167 2477 1183
rect 2495 1167 2511 1183
rect 2529 1167 2545 1183
rect 2563 1167 2579 1183
rect 2597 1167 2613 1183
rect 2631 1167 2647 1183
rect 2665 1167 2681 1183
rect 2699 1167 2715 1183
rect 2733 1167 2749 1183
rect 2767 1167 2783 1183
rect 2801 1167 2817 1183
rect 2835 1167 2851 1183
rect 2869 1167 2885 1183
rect 2903 1167 2919 1183
rect 2937 1167 2953 1183
rect 2971 1167 2987 1183
rect 3005 1167 3021 1183
rect 3039 1167 3055 1183
rect 3073 1167 3089 1183
rect 3107 1167 3123 1183
rect 3141 1167 3157 1183
rect 3175 1167 3191 1183
rect 3209 1167 3225 1183
rect 3243 1167 3259 1183
rect 3277 1167 3293 1183
rect 3311 1167 3327 1183
rect 3345 1167 3361 1183
rect 3379 1167 3395 1183
rect 3413 1167 3429 1183
rect 3447 1167 3463 1183
rect -157 1117 -141 1133
rect -157 1083 -141 1099
rect -157 1049 -141 1065
rect -157 1015 -141 1031
rect 3447 1117 3463 1133
rect 3447 1083 3463 1099
rect 3447 1049 3463 1065
rect -157 981 -141 997
rect -157 947 -141 963
rect -157 913 -141 929
rect -157 879 -141 895
rect -157 845 -141 861
rect -157 811 -141 827
rect -157 777 -141 793
rect -157 743 -141 759
rect -157 709 -141 725
rect -157 675 -141 691
rect -157 641 -141 657
rect -157 607 -141 623
rect -157 573 -141 589
rect -157 539 -141 555
rect -157 505 -141 521
rect -157 471 -141 487
rect -157 437 -141 453
rect -157 403 -141 419
rect -157 369 -141 385
rect -157 335 -141 351
rect -157 301 -141 317
rect -157 267 -141 283
rect -157 233 -141 249
rect -157 199 -141 215
rect -157 165 -141 181
rect -157 131 -141 147
rect -157 97 -141 113
rect -157 63 -141 79
rect -157 29 -141 45
rect -157 -5 -141 11
rect 3447 1015 3463 1031
rect 3447 981 3463 997
rect 3447 947 3463 963
rect 3447 913 3463 929
rect 3447 879 3463 895
rect 3447 845 3463 861
rect 3447 811 3463 827
rect 3447 777 3463 793
rect 3447 743 3463 759
rect 3447 709 3463 725
rect 3447 675 3463 691
rect 3447 641 3463 657
rect 3447 607 3463 623
rect 3447 573 3463 589
rect 3447 539 3463 555
rect 3447 505 3463 521
rect 3447 471 3463 487
rect 3447 437 3463 453
rect 3447 403 3463 419
rect 3447 369 3463 385
rect 3447 335 3463 351
rect 3447 301 3463 317
rect 3447 267 3463 283
rect 3447 233 3463 249
rect 3447 199 3463 215
rect 3447 165 3463 181
rect 3447 131 3463 147
rect 3447 97 3463 113
rect 3447 63 3463 79
rect 3447 29 3463 45
rect -157 -39 -141 -23
rect -157 -73 -141 -57
rect -157 -107 -141 -91
rect 3447 -5 3463 11
rect 3447 -39 3463 -23
rect 3447 -73 3463 -57
rect 3447 -107 3463 -91
rect -157 -157 -141 -141
rect -123 -157 -107 -141
rect -89 -157 -73 -141
rect -55 -157 -39 -141
rect -21 -157 -5 -141
rect 13 -157 29 -141
rect 47 -157 63 -141
rect 81 -157 97 -141
rect 115 -157 131 -141
rect 149 -157 165 -141
rect 183 -157 199 -141
rect 217 -157 233 -141
rect 251 -157 267 -141
rect 285 -157 301 -141
rect 319 -157 335 -141
rect 353 -157 369 -141
rect 387 -157 403 -141
rect 421 -157 437 -141
rect 455 -157 471 -141
rect 489 -157 505 -141
rect 523 -157 539 -141
rect 557 -157 573 -141
rect 591 -157 607 -141
rect 625 -157 641 -141
rect 659 -157 675 -141
rect 693 -157 709 -141
rect 727 -157 743 -141
rect 761 -157 777 -141
rect 795 -157 811 -141
rect 829 -157 845 -141
rect 863 -157 879 -141
rect 897 -157 913 -141
rect 931 -157 947 -141
rect 965 -157 981 -141
rect 999 -157 1015 -141
rect 1033 -157 1049 -141
rect 1067 -157 1083 -141
rect 1101 -157 1117 -141
rect 1135 -157 1151 -141
rect 1169 -157 1185 -141
rect 1203 -157 1219 -141
rect 1237 -157 1253 -141
rect 1271 -157 1287 -141
rect 1305 -157 1321 -141
rect 1339 -157 1355 -141
rect 1373 -157 1389 -141
rect 1407 -157 1423 -141
rect 1441 -157 1457 -141
rect 1475 -157 1491 -141
rect 1509 -157 1525 -141
rect 1543 -157 1559 -141
rect 1577 -157 1593 -141
rect 1611 -157 1627 -141
rect 1645 -157 1661 -141
rect 1679 -157 1695 -141
rect 1713 -157 1729 -141
rect 1747 -157 1763 -141
rect 1781 -157 1797 -141
rect 1815 -157 1831 -141
rect 1849 -157 1865 -141
rect 1883 -157 1899 -141
rect 1917 -157 1933 -141
rect 1951 -157 1967 -141
rect 1985 -157 2001 -141
rect 2019 -157 2035 -141
rect 2053 -157 2069 -141
rect 2087 -157 2103 -141
rect 2121 -157 2137 -141
rect 2155 -157 2171 -141
rect 2189 -157 2205 -141
rect 2223 -157 2239 -141
rect 2257 -157 2273 -141
rect 2291 -157 2307 -141
rect 2325 -157 2341 -141
rect 2359 -157 2375 -141
rect 2393 -157 2409 -141
rect 2427 -157 2443 -141
rect 2461 -157 2477 -141
rect 2495 -157 2511 -141
rect 2529 -157 2545 -141
rect 2563 -157 2579 -141
rect 2597 -157 2613 -141
rect 2631 -157 2647 -141
rect 2665 -157 2681 -141
rect 2699 -157 2715 -141
rect 2733 -157 2749 -141
rect 2767 -157 2783 -141
rect 2801 -157 2817 -141
rect 2835 -157 2851 -141
rect 2869 -157 2885 -141
rect 2903 -157 2919 -141
rect 2937 -157 2953 -141
rect 2971 -157 2987 -141
rect 3005 -157 3021 -141
rect 3039 -157 3055 -141
rect 3073 -157 3089 -141
rect 3107 -157 3123 -141
rect 3141 -157 3157 -141
rect 3175 -157 3191 -141
rect 3209 -157 3225 -141
rect 3243 -157 3259 -141
rect 3277 -157 3293 -141
rect 3311 -157 3327 -141
rect 3345 -157 3361 -141
rect 3379 -157 3395 -141
rect 3413 -157 3429 -141
rect 3447 -157 3463 -141
<< nsubdiffcont >>
rect 21 998 37 1014
rect 55 998 71 1014
rect 89 998 105 1014
rect 149 989 165 1005
rect 183 989 199 1005
rect 217 989 233 1005
rect 251 989 267 1005
rect 285 989 301 1005
rect 319 989 335 1005
rect 353 989 369 1005
rect 387 989 403 1005
rect 421 989 437 1005
rect 455 989 471 1005
rect 489 989 505 1005
rect 523 989 539 1005
rect 557 989 573 1005
rect 591 989 607 1005
rect 625 989 641 1005
rect 659 989 675 1005
rect 693 989 709 1005
rect 727 989 743 1005
rect 761 989 777 1005
rect 795 989 811 1005
rect 829 989 845 1005
rect 863 989 879 1005
rect 897 989 913 1005
rect 931 989 947 1005
rect 965 989 981 1005
rect 999 989 1015 1005
rect 1033 989 1049 1005
rect 1067 989 1083 1005
rect 1101 989 1117 1005
rect 1135 989 1151 1005
rect 1169 989 1185 1005
rect 1203 989 1219 1005
rect 1237 989 1253 1005
rect 1271 989 1287 1005
rect 1305 989 1321 1005
rect 1339 989 1355 1005
rect 1373 989 1389 1005
rect 1407 989 1423 1005
rect 1441 989 1457 1005
rect 1475 989 1491 1005
rect 1509 989 1525 1005
rect 1543 989 1559 1005
rect 1577 989 1593 1005
rect 1611 989 1627 1005
rect 1645 989 1661 1005
rect 1679 989 1695 1005
rect 1713 989 1729 1005
rect 1747 989 1763 1005
rect 1781 989 1797 1005
rect 1815 989 1831 1005
rect 1849 989 1865 1005
rect 1883 989 1899 1005
rect 1917 989 1933 1005
rect 1951 989 1967 1005
rect 1985 989 2001 1005
rect 2019 989 2035 1005
rect 2053 989 2069 1005
rect 2087 989 2103 1005
rect 2121 989 2137 1005
rect 2155 989 2171 1005
rect 2189 989 2205 1005
rect 2223 989 2239 1005
rect 2257 989 2273 1005
rect 2291 989 2307 1005
rect 2325 989 2341 1005
rect 2359 989 2375 1005
rect 2393 989 2409 1005
rect 2427 989 2443 1005
rect 2461 989 2477 1005
rect 2495 989 2511 1005
rect 2529 989 2545 1005
rect 2563 989 2579 1005
rect 2597 989 2613 1005
rect 2631 989 2647 1005
rect 2665 989 2681 1005
rect 2699 989 2715 1005
rect 2733 989 2749 1005
rect 2767 989 2783 1005
rect 2801 989 2817 1005
rect 2835 989 2851 1005
rect 2869 989 2885 1005
rect 2903 989 2919 1005
rect 2937 989 2953 1005
rect 2971 989 2987 1005
rect 3005 989 3021 1005
rect 3039 989 3055 1005
rect 3073 989 3089 1005
rect 3107 989 3123 1005
rect 3141 989 3157 1005
rect 3201 998 3217 1014
rect 3235 998 3251 1014
rect 3269 998 3285 1014
rect 21 964 37 980
rect 55 964 71 980
rect 89 964 105 980
rect 149 955 165 971
rect 183 955 199 971
rect 217 955 233 971
rect 251 955 267 971
rect 285 955 301 971
rect 319 955 335 971
rect 353 955 369 971
rect 387 955 403 971
rect 421 955 437 971
rect 455 955 471 971
rect 489 955 505 971
rect 523 955 539 971
rect 557 955 573 971
rect 591 955 607 971
rect 625 955 641 971
rect 659 955 675 971
rect 693 955 709 971
rect 727 955 743 971
rect 761 955 777 971
rect 795 955 811 971
rect 829 955 845 971
rect 863 955 879 971
rect 897 955 913 971
rect 931 955 947 971
rect 965 955 981 971
rect 999 955 1015 971
rect 1033 955 1049 971
rect 1067 955 1083 971
rect 1101 955 1117 971
rect 1135 955 1151 971
rect 1169 955 1185 971
rect 1203 955 1219 971
rect 1237 955 1253 971
rect 1271 955 1287 971
rect 1305 955 1321 971
rect 1339 955 1355 971
rect 1373 955 1389 971
rect 1407 955 1423 971
rect 1441 955 1457 971
rect 1475 955 1491 971
rect 1509 955 1525 971
rect 1543 955 1559 971
rect 1577 955 1593 971
rect 1611 955 1627 971
rect 1645 955 1661 971
rect 1679 955 1695 971
rect 1713 955 1729 971
rect 1747 955 1763 971
rect 1781 955 1797 971
rect 1815 955 1831 971
rect 1849 955 1865 971
rect 1883 955 1899 971
rect 1917 955 1933 971
rect 1951 955 1967 971
rect 1985 955 2001 971
rect 2019 955 2035 971
rect 2053 955 2069 971
rect 2087 955 2103 971
rect 2121 955 2137 971
rect 2155 955 2171 971
rect 2189 955 2205 971
rect 2223 955 2239 971
rect 2257 955 2273 971
rect 2291 955 2307 971
rect 2325 955 2341 971
rect 2359 955 2375 971
rect 2393 955 2409 971
rect 2427 955 2443 971
rect 2461 955 2477 971
rect 2495 955 2511 971
rect 2529 955 2545 971
rect 2563 955 2579 971
rect 2597 955 2613 971
rect 2631 955 2647 971
rect 2665 955 2681 971
rect 2699 955 2715 971
rect 2733 955 2749 971
rect 2767 955 2783 971
rect 2801 955 2817 971
rect 2835 955 2851 971
rect 2869 955 2885 971
rect 2903 955 2919 971
rect 2937 955 2953 971
rect 2971 955 2987 971
rect 3005 955 3021 971
rect 3039 955 3055 971
rect 3073 955 3089 971
rect 3107 955 3123 971
rect 3141 955 3157 971
rect 3201 964 3217 980
rect 3235 964 3251 980
rect 3269 964 3285 980
rect 21 930 37 946
rect 55 930 71 946
rect 89 930 105 946
rect 149 921 165 937
rect 183 921 199 937
rect 217 921 233 937
rect 251 921 267 937
rect 285 921 301 937
rect 319 921 335 937
rect 353 921 369 937
rect 387 921 403 937
rect 421 921 437 937
rect 455 921 471 937
rect 489 921 505 937
rect 523 921 539 937
rect 557 921 573 937
rect 591 921 607 937
rect 625 921 641 937
rect 659 921 675 937
rect 693 921 709 937
rect 727 921 743 937
rect 761 921 777 937
rect 795 921 811 937
rect 829 921 845 937
rect 863 921 879 937
rect 897 921 913 937
rect 931 921 947 937
rect 965 921 981 937
rect 999 921 1015 937
rect 1033 921 1049 937
rect 1067 921 1083 937
rect 1101 921 1117 937
rect 1135 921 1151 937
rect 1169 921 1185 937
rect 1203 921 1219 937
rect 1237 921 1253 937
rect 1271 921 1287 937
rect 1305 921 1321 937
rect 1339 921 1355 937
rect 1373 921 1389 937
rect 1407 921 1423 937
rect 1441 921 1457 937
rect 1475 921 1491 937
rect 1509 921 1525 937
rect 1543 921 1559 937
rect 1577 921 1593 937
rect 1611 921 1627 937
rect 1645 921 1661 937
rect 1679 921 1695 937
rect 1713 921 1729 937
rect 1747 921 1763 937
rect 1781 921 1797 937
rect 1815 921 1831 937
rect 1849 921 1865 937
rect 1883 921 1899 937
rect 1917 921 1933 937
rect 1951 921 1967 937
rect 1985 921 2001 937
rect 2019 921 2035 937
rect 2053 921 2069 937
rect 2087 921 2103 937
rect 2121 921 2137 937
rect 2155 921 2171 937
rect 2189 921 2205 937
rect 2223 921 2239 937
rect 2257 921 2273 937
rect 2291 921 2307 937
rect 2325 921 2341 937
rect 2359 921 2375 937
rect 2393 921 2409 937
rect 2427 921 2443 937
rect 2461 921 2477 937
rect 2495 921 2511 937
rect 2529 921 2545 937
rect 2563 921 2579 937
rect 2597 921 2613 937
rect 2631 921 2647 937
rect 2665 921 2681 937
rect 2699 921 2715 937
rect 2733 921 2749 937
rect 2767 921 2783 937
rect 2801 921 2817 937
rect 2835 921 2851 937
rect 2869 921 2885 937
rect 2903 921 2919 937
rect 2937 921 2953 937
rect 2971 921 2987 937
rect 3005 921 3021 937
rect 3039 921 3055 937
rect 3073 921 3089 937
rect 3107 921 3123 937
rect 3141 921 3157 937
rect 3201 930 3217 946
rect 3235 930 3251 946
rect 3269 930 3285 946
rect 21 896 37 912
rect 55 896 71 912
rect 89 896 105 912
rect 21 862 37 878
rect 55 862 71 878
rect 89 862 105 878
rect 21 828 37 844
rect 55 828 71 844
rect 89 828 105 844
rect 21 794 37 810
rect 55 794 71 810
rect 89 794 105 810
rect 3201 896 3217 912
rect 3235 896 3251 912
rect 3269 896 3285 912
rect 3201 862 3217 878
rect 3235 862 3251 878
rect 3269 862 3285 878
rect 3201 828 3217 844
rect 3235 828 3251 844
rect 3269 828 3285 844
rect 21 760 37 776
rect 55 760 71 776
rect 89 760 105 776
rect 21 726 37 742
rect 55 726 71 742
rect 89 726 105 742
rect 21 692 37 708
rect 55 692 71 708
rect 89 692 105 708
rect 3201 794 3217 810
rect 3235 794 3251 810
rect 3269 794 3285 810
rect 3201 760 3217 776
rect 3235 760 3251 776
rect 3269 760 3285 776
rect 3201 726 3217 742
rect 3235 726 3251 742
rect 3269 726 3285 742
rect 3201 692 3217 708
rect 3235 692 3251 708
rect 3269 692 3285 708
rect 21 658 37 674
rect 55 658 71 674
rect 89 658 105 674
rect 21 624 37 640
rect 55 624 71 640
rect 89 624 105 640
rect 21 590 37 606
rect 55 590 71 606
rect 89 590 105 606
rect 3201 658 3217 674
rect 3235 658 3251 674
rect 3269 658 3285 674
rect 3201 624 3217 640
rect 3235 624 3251 640
rect 3269 624 3285 640
rect 3201 590 3217 606
rect 3235 590 3251 606
rect 3269 590 3285 606
rect 21 556 37 572
rect 55 556 71 572
rect 89 556 105 572
rect 3201 556 3217 572
rect 3235 556 3251 572
rect 3269 556 3285 572
rect 149 539 165 555
rect 183 539 199 555
rect 217 539 233 555
rect 251 539 267 555
rect 285 539 301 555
rect 319 539 335 555
rect 353 539 369 555
rect 387 539 403 555
rect 421 539 437 555
rect 455 539 471 555
rect 489 539 505 555
rect 523 539 539 555
rect 557 539 573 555
rect 591 539 607 555
rect 625 539 641 555
rect 659 539 675 555
rect 693 539 709 555
rect 727 539 743 555
rect 761 539 777 555
rect 795 539 811 555
rect 829 539 845 555
rect 863 539 879 555
rect 897 539 913 555
rect 931 539 947 555
rect 965 539 981 555
rect 999 539 1015 555
rect 1033 539 1049 555
rect 1067 539 1083 555
rect 1101 539 1117 555
rect 1135 539 1151 555
rect 1169 539 1185 555
rect 1203 539 1219 555
rect 1237 539 1253 555
rect 1271 539 1287 555
rect 1305 539 1321 555
rect 1339 539 1355 555
rect 1373 539 1389 555
rect 1407 539 1423 555
rect 1441 539 1457 555
rect 1475 539 1491 555
rect 1509 539 1525 555
rect 1543 539 1559 555
rect 1577 539 1593 555
rect 1611 539 1627 555
rect 1645 539 1661 555
rect 1679 539 1695 555
rect 1713 539 1729 555
rect 1747 539 1763 555
rect 1781 539 1797 555
rect 1815 539 1831 555
rect 1849 539 1865 555
rect 1883 539 1899 555
rect 1917 539 1933 555
rect 1951 539 1967 555
rect 1985 539 2001 555
rect 2019 539 2035 555
rect 2053 539 2069 555
rect 2087 539 2103 555
rect 2121 539 2137 555
rect 2155 539 2171 555
rect 2189 539 2205 555
rect 2223 539 2239 555
rect 2257 539 2273 555
rect 2291 539 2307 555
rect 2325 539 2341 555
rect 2359 539 2375 555
rect 2393 539 2409 555
rect 2427 539 2443 555
rect 2461 539 2477 555
rect 2495 539 2511 555
rect 2529 539 2545 555
rect 2563 539 2579 555
rect 2597 539 2613 555
rect 2631 539 2647 555
rect 2665 539 2681 555
rect 2699 539 2715 555
rect 2733 539 2749 555
rect 2767 539 2783 555
rect 2801 539 2817 555
rect 2835 539 2851 555
rect 2869 539 2885 555
rect 2903 539 2919 555
rect 2937 539 2953 555
rect 2971 539 2987 555
rect 3005 539 3021 555
rect 3039 539 3055 555
rect 3073 539 3089 555
rect 3107 539 3123 555
rect 3141 539 3157 555
rect 21 522 37 538
rect 55 522 71 538
rect 89 522 105 538
rect 3201 522 3217 538
rect 3235 522 3251 538
rect 3269 522 3285 538
rect 149 505 165 521
rect 183 505 199 521
rect 217 505 233 521
rect 251 505 267 521
rect 285 505 301 521
rect 319 505 335 521
rect 353 505 369 521
rect 387 505 403 521
rect 421 505 437 521
rect 455 505 471 521
rect 489 505 505 521
rect 523 505 539 521
rect 557 505 573 521
rect 591 505 607 521
rect 625 505 641 521
rect 659 505 675 521
rect 693 505 709 521
rect 727 505 743 521
rect 761 505 777 521
rect 795 505 811 521
rect 829 505 845 521
rect 863 505 879 521
rect 897 505 913 521
rect 931 505 947 521
rect 965 505 981 521
rect 999 505 1015 521
rect 1033 505 1049 521
rect 1067 505 1083 521
rect 1101 505 1117 521
rect 1135 505 1151 521
rect 1169 505 1185 521
rect 1203 505 1219 521
rect 1237 505 1253 521
rect 1271 505 1287 521
rect 1305 505 1321 521
rect 1339 505 1355 521
rect 1373 505 1389 521
rect 1407 505 1423 521
rect 1441 505 1457 521
rect 1475 505 1491 521
rect 1509 505 1525 521
rect 1543 505 1559 521
rect 1577 505 1593 521
rect 1611 505 1627 521
rect 1645 505 1661 521
rect 1679 505 1695 521
rect 1713 505 1729 521
rect 1747 505 1763 521
rect 1781 505 1797 521
rect 1815 505 1831 521
rect 1849 505 1865 521
rect 1883 505 1899 521
rect 1917 505 1933 521
rect 1951 505 1967 521
rect 1985 505 2001 521
rect 2019 505 2035 521
rect 2053 505 2069 521
rect 2087 505 2103 521
rect 2121 505 2137 521
rect 2155 505 2171 521
rect 2189 505 2205 521
rect 2223 505 2239 521
rect 2257 505 2273 521
rect 2291 505 2307 521
rect 2325 505 2341 521
rect 2359 505 2375 521
rect 2393 505 2409 521
rect 2427 505 2443 521
rect 2461 505 2477 521
rect 2495 505 2511 521
rect 2529 505 2545 521
rect 2563 505 2579 521
rect 2597 505 2613 521
rect 2631 505 2647 521
rect 2665 505 2681 521
rect 2699 505 2715 521
rect 2733 505 2749 521
rect 2767 505 2783 521
rect 2801 505 2817 521
rect 2835 505 2851 521
rect 2869 505 2885 521
rect 2903 505 2919 521
rect 2937 505 2953 521
rect 2971 505 2987 521
rect 3005 505 3021 521
rect 3039 505 3055 521
rect 3073 505 3089 521
rect 3107 505 3123 521
rect 3141 505 3157 521
rect 21 488 37 504
rect 55 488 71 504
rect 89 488 105 504
rect 3201 488 3217 504
rect 3235 488 3251 504
rect 3269 488 3285 504
rect 149 471 165 487
rect 183 471 199 487
rect 217 471 233 487
rect 251 471 267 487
rect 285 471 301 487
rect 319 471 335 487
rect 353 471 369 487
rect 387 471 403 487
rect 421 471 437 487
rect 455 471 471 487
rect 489 471 505 487
rect 523 471 539 487
rect 557 471 573 487
rect 591 471 607 487
rect 625 471 641 487
rect 659 471 675 487
rect 693 471 709 487
rect 727 471 743 487
rect 761 471 777 487
rect 795 471 811 487
rect 829 471 845 487
rect 863 471 879 487
rect 897 471 913 487
rect 931 471 947 487
rect 965 471 981 487
rect 999 471 1015 487
rect 1033 471 1049 487
rect 1067 471 1083 487
rect 1101 471 1117 487
rect 1135 471 1151 487
rect 1169 471 1185 487
rect 1203 471 1219 487
rect 1237 471 1253 487
rect 1271 471 1287 487
rect 1305 471 1321 487
rect 1339 471 1355 487
rect 1373 471 1389 487
rect 1407 471 1423 487
rect 1441 471 1457 487
rect 1475 471 1491 487
rect 1509 471 1525 487
rect 1543 471 1559 487
rect 1577 471 1593 487
rect 1611 471 1627 487
rect 1645 471 1661 487
rect 1679 471 1695 487
rect 1713 471 1729 487
rect 1747 471 1763 487
rect 1781 471 1797 487
rect 1815 471 1831 487
rect 1849 471 1865 487
rect 1883 471 1899 487
rect 1917 471 1933 487
rect 1951 471 1967 487
rect 1985 471 2001 487
rect 2019 471 2035 487
rect 2053 471 2069 487
rect 2087 471 2103 487
rect 2121 471 2137 487
rect 2155 471 2171 487
rect 2189 471 2205 487
rect 2223 471 2239 487
rect 2257 471 2273 487
rect 2291 471 2307 487
rect 2325 471 2341 487
rect 2359 471 2375 487
rect 2393 471 2409 487
rect 2427 471 2443 487
rect 2461 471 2477 487
rect 2495 471 2511 487
rect 2529 471 2545 487
rect 2563 471 2579 487
rect 2597 471 2613 487
rect 2631 471 2647 487
rect 2665 471 2681 487
rect 2699 471 2715 487
rect 2733 471 2749 487
rect 2767 471 2783 487
rect 2801 471 2817 487
rect 2835 471 2851 487
rect 2869 471 2885 487
rect 2903 471 2919 487
rect 2937 471 2953 487
rect 2971 471 2987 487
rect 3005 471 3021 487
rect 3039 471 3055 487
rect 3073 471 3089 487
rect 3107 471 3123 487
rect 3141 471 3157 487
rect 21 454 37 470
rect 55 454 71 470
rect 89 454 105 470
rect 3201 454 3217 470
rect 3235 454 3251 470
rect 3269 454 3285 470
rect 21 420 37 436
rect 55 420 71 436
rect 89 420 105 436
rect 21 386 37 402
rect 55 386 71 402
rect 89 386 105 402
rect 21 352 37 368
rect 55 352 71 368
rect 89 352 105 368
rect 3201 420 3217 436
rect 3235 420 3251 436
rect 3269 420 3285 436
rect 3201 386 3217 402
rect 3235 386 3251 402
rect 3269 386 3285 402
rect 3201 352 3217 368
rect 3235 352 3251 368
rect 3269 352 3285 368
rect 21 318 37 334
rect 55 318 71 334
rect 89 318 105 334
rect 21 284 37 300
rect 55 284 71 300
rect 89 284 105 300
rect 21 250 37 266
rect 55 250 71 266
rect 89 250 105 266
rect 21 216 37 232
rect 55 216 71 232
rect 89 216 105 232
rect 3201 318 3217 334
rect 3235 318 3251 334
rect 3269 318 3285 334
rect 3201 284 3217 300
rect 3235 284 3251 300
rect 3269 284 3285 300
rect 3201 250 3217 266
rect 3235 250 3251 266
rect 3269 250 3285 266
rect 21 182 37 198
rect 55 182 71 198
rect 89 182 105 198
rect 21 148 37 164
rect 55 148 71 164
rect 89 148 105 164
rect 21 114 37 130
rect 55 114 71 130
rect 89 114 105 130
rect 3201 216 3217 232
rect 3235 216 3251 232
rect 3269 216 3285 232
rect 3201 182 3217 198
rect 3235 182 3251 198
rect 3269 182 3285 198
rect 3201 148 3217 164
rect 3235 148 3251 164
rect 3269 148 3285 164
rect 3201 114 3217 130
rect 3235 114 3251 130
rect 3269 114 3285 130
rect 21 80 37 96
rect 55 80 71 96
rect 89 80 105 96
rect 149 89 165 105
rect 183 89 199 105
rect 217 89 233 105
rect 251 89 267 105
rect 285 89 301 105
rect 319 89 335 105
rect 353 89 369 105
rect 387 89 403 105
rect 421 89 437 105
rect 455 89 471 105
rect 489 89 505 105
rect 523 89 539 105
rect 557 89 573 105
rect 591 89 607 105
rect 625 89 641 105
rect 659 89 675 105
rect 693 89 709 105
rect 727 89 743 105
rect 761 89 777 105
rect 795 89 811 105
rect 829 89 845 105
rect 863 89 879 105
rect 897 89 913 105
rect 931 89 947 105
rect 965 89 981 105
rect 999 89 1015 105
rect 1033 89 1049 105
rect 1067 89 1083 105
rect 1101 89 1117 105
rect 1135 89 1151 105
rect 1169 89 1185 105
rect 1203 89 1219 105
rect 1237 89 1253 105
rect 1271 89 1287 105
rect 1305 89 1321 105
rect 1339 89 1355 105
rect 1373 89 1389 105
rect 1407 89 1423 105
rect 1441 89 1457 105
rect 1475 89 1491 105
rect 1509 89 1525 105
rect 1543 89 1559 105
rect 1577 89 1593 105
rect 1611 89 1627 105
rect 1645 89 1661 105
rect 1679 89 1695 105
rect 1713 89 1729 105
rect 1747 89 1763 105
rect 1781 89 1797 105
rect 1815 89 1831 105
rect 1849 89 1865 105
rect 1883 89 1899 105
rect 1917 89 1933 105
rect 1951 89 1967 105
rect 1985 89 2001 105
rect 2019 89 2035 105
rect 2053 89 2069 105
rect 2087 89 2103 105
rect 2121 89 2137 105
rect 2155 89 2171 105
rect 2189 89 2205 105
rect 2223 89 2239 105
rect 2257 89 2273 105
rect 2291 89 2307 105
rect 2325 89 2341 105
rect 2359 89 2375 105
rect 2393 89 2409 105
rect 2427 89 2443 105
rect 2461 89 2477 105
rect 2495 89 2511 105
rect 2529 89 2545 105
rect 2563 89 2579 105
rect 2597 89 2613 105
rect 2631 89 2647 105
rect 2665 89 2681 105
rect 2699 89 2715 105
rect 2733 89 2749 105
rect 2767 89 2783 105
rect 2801 89 2817 105
rect 2835 89 2851 105
rect 2869 89 2885 105
rect 2903 89 2919 105
rect 2937 89 2953 105
rect 2971 89 2987 105
rect 3005 89 3021 105
rect 3039 89 3055 105
rect 3073 89 3089 105
rect 3107 89 3123 105
rect 3141 89 3157 105
rect 3201 80 3217 96
rect 3235 80 3251 96
rect 3269 80 3285 96
rect 21 46 37 62
rect 55 46 71 62
rect 89 46 105 62
rect 149 55 165 71
rect 183 55 199 71
rect 217 55 233 71
rect 251 55 267 71
rect 285 55 301 71
rect 319 55 335 71
rect 353 55 369 71
rect 387 55 403 71
rect 421 55 437 71
rect 455 55 471 71
rect 489 55 505 71
rect 523 55 539 71
rect 557 55 573 71
rect 591 55 607 71
rect 625 55 641 71
rect 659 55 675 71
rect 693 55 709 71
rect 727 55 743 71
rect 761 55 777 71
rect 795 55 811 71
rect 829 55 845 71
rect 863 55 879 71
rect 897 55 913 71
rect 931 55 947 71
rect 965 55 981 71
rect 999 55 1015 71
rect 1033 55 1049 71
rect 1067 55 1083 71
rect 1101 55 1117 71
rect 1135 55 1151 71
rect 1169 55 1185 71
rect 1203 55 1219 71
rect 1237 55 1253 71
rect 1271 55 1287 71
rect 1305 55 1321 71
rect 1339 55 1355 71
rect 1373 55 1389 71
rect 1407 55 1423 71
rect 1441 55 1457 71
rect 1475 55 1491 71
rect 1509 55 1525 71
rect 1543 55 1559 71
rect 1577 55 1593 71
rect 1611 55 1627 71
rect 1645 55 1661 71
rect 1679 55 1695 71
rect 1713 55 1729 71
rect 1747 55 1763 71
rect 1781 55 1797 71
rect 1815 55 1831 71
rect 1849 55 1865 71
rect 1883 55 1899 71
rect 1917 55 1933 71
rect 1951 55 1967 71
rect 1985 55 2001 71
rect 2019 55 2035 71
rect 2053 55 2069 71
rect 2087 55 2103 71
rect 2121 55 2137 71
rect 2155 55 2171 71
rect 2189 55 2205 71
rect 2223 55 2239 71
rect 2257 55 2273 71
rect 2291 55 2307 71
rect 2325 55 2341 71
rect 2359 55 2375 71
rect 2393 55 2409 71
rect 2427 55 2443 71
rect 2461 55 2477 71
rect 2495 55 2511 71
rect 2529 55 2545 71
rect 2563 55 2579 71
rect 2597 55 2613 71
rect 2631 55 2647 71
rect 2665 55 2681 71
rect 2699 55 2715 71
rect 2733 55 2749 71
rect 2767 55 2783 71
rect 2801 55 2817 71
rect 2835 55 2851 71
rect 2869 55 2885 71
rect 2903 55 2919 71
rect 2937 55 2953 71
rect 2971 55 2987 71
rect 3005 55 3021 71
rect 3039 55 3055 71
rect 3073 55 3089 71
rect 3107 55 3123 71
rect 3141 55 3157 71
rect 3201 46 3217 62
rect 3235 46 3251 62
rect 3269 46 3285 62
rect 21 12 37 28
rect 55 12 71 28
rect 89 12 105 28
rect 149 21 165 37
rect 183 21 199 37
rect 217 21 233 37
rect 251 21 267 37
rect 285 21 301 37
rect 319 21 335 37
rect 353 21 369 37
rect 387 21 403 37
rect 421 21 437 37
rect 455 21 471 37
rect 489 21 505 37
rect 523 21 539 37
rect 557 21 573 37
rect 591 21 607 37
rect 625 21 641 37
rect 659 21 675 37
rect 693 21 709 37
rect 727 21 743 37
rect 761 21 777 37
rect 795 21 811 37
rect 829 21 845 37
rect 863 21 879 37
rect 897 21 913 37
rect 931 21 947 37
rect 965 21 981 37
rect 999 21 1015 37
rect 1033 21 1049 37
rect 1067 21 1083 37
rect 1101 21 1117 37
rect 1135 21 1151 37
rect 1169 21 1185 37
rect 1203 21 1219 37
rect 1237 21 1253 37
rect 1271 21 1287 37
rect 1305 21 1321 37
rect 1339 21 1355 37
rect 1373 21 1389 37
rect 1407 21 1423 37
rect 1441 21 1457 37
rect 1475 21 1491 37
rect 1509 21 1525 37
rect 1543 21 1559 37
rect 1577 21 1593 37
rect 1611 21 1627 37
rect 1645 21 1661 37
rect 1679 21 1695 37
rect 1713 21 1729 37
rect 1747 21 1763 37
rect 1781 21 1797 37
rect 1815 21 1831 37
rect 1849 21 1865 37
rect 1883 21 1899 37
rect 1917 21 1933 37
rect 1951 21 1967 37
rect 1985 21 2001 37
rect 2019 21 2035 37
rect 2053 21 2069 37
rect 2087 21 2103 37
rect 2121 21 2137 37
rect 2155 21 2171 37
rect 2189 21 2205 37
rect 2223 21 2239 37
rect 2257 21 2273 37
rect 2291 21 2307 37
rect 2325 21 2341 37
rect 2359 21 2375 37
rect 2393 21 2409 37
rect 2427 21 2443 37
rect 2461 21 2477 37
rect 2495 21 2511 37
rect 2529 21 2545 37
rect 2563 21 2579 37
rect 2597 21 2613 37
rect 2631 21 2647 37
rect 2665 21 2681 37
rect 2699 21 2715 37
rect 2733 21 2749 37
rect 2767 21 2783 37
rect 2801 21 2817 37
rect 2835 21 2851 37
rect 2869 21 2885 37
rect 2903 21 2919 37
rect 2937 21 2953 37
rect 2971 21 2987 37
rect 3005 21 3021 37
rect 3039 21 3055 37
rect 3073 21 3089 37
rect 3107 21 3123 37
rect 3141 21 3157 37
rect 3201 12 3217 28
rect 3235 12 3251 28
rect 3269 12 3285 28
<< pdiode >>
rect 264 780 3042 801
rect 264 764 285 780
rect 301 764 319 780
rect 335 764 353 780
rect 369 764 387 780
rect 403 764 421 780
rect 437 764 455 780
rect 471 764 489 780
rect 505 764 523 780
rect 539 764 557 780
rect 573 764 591 780
rect 607 764 625 780
rect 641 764 659 780
rect 675 764 693 780
rect 709 764 727 780
rect 743 764 761 780
rect 777 764 795 780
rect 811 764 829 780
rect 845 764 863 780
rect 879 764 897 780
rect 913 764 931 780
rect 947 764 965 780
rect 981 764 999 780
rect 1015 764 1033 780
rect 1049 764 1067 780
rect 1083 764 1101 780
rect 1117 764 1135 780
rect 1151 764 1169 780
rect 1185 764 1203 780
rect 1219 764 1237 780
rect 1253 764 1271 780
rect 1287 764 1305 780
rect 1321 764 1339 780
rect 1355 764 1373 780
rect 1389 764 1407 780
rect 1423 764 1441 780
rect 1457 764 1475 780
rect 1491 764 1509 780
rect 1525 764 1543 780
rect 1559 764 1577 780
rect 1593 764 1611 780
rect 1627 764 1645 780
rect 1661 764 1679 780
rect 1695 764 1713 780
rect 1729 764 1747 780
rect 1763 764 1781 780
rect 1797 764 1815 780
rect 1831 764 1849 780
rect 1865 764 1883 780
rect 1899 764 1917 780
rect 1933 764 1951 780
rect 1967 764 1985 780
rect 2001 764 2019 780
rect 2035 764 2053 780
rect 2069 764 2087 780
rect 2103 764 2121 780
rect 2137 764 2155 780
rect 2171 764 2189 780
rect 2205 764 2223 780
rect 2239 764 2257 780
rect 2273 764 2291 780
rect 2307 764 2325 780
rect 2341 764 2359 780
rect 2375 764 2393 780
rect 2409 764 2427 780
rect 2443 764 2461 780
rect 2477 764 2495 780
rect 2511 764 2529 780
rect 2545 764 2563 780
rect 2579 764 2597 780
rect 2613 764 2631 780
rect 2647 764 2665 780
rect 2681 764 2699 780
rect 2715 764 2733 780
rect 2749 764 2767 780
rect 2783 764 2801 780
rect 2817 764 2835 780
rect 2851 764 2869 780
rect 2885 764 2903 780
rect 2919 764 2937 780
rect 2953 764 2971 780
rect 2987 764 3005 780
rect 3021 764 3042 780
rect 264 746 3042 764
rect 264 730 285 746
rect 301 730 319 746
rect 335 730 353 746
rect 369 730 387 746
rect 403 730 421 746
rect 437 730 455 746
rect 471 730 489 746
rect 505 730 523 746
rect 539 730 557 746
rect 573 730 591 746
rect 607 730 625 746
rect 641 730 659 746
rect 675 730 693 746
rect 709 730 727 746
rect 743 730 761 746
rect 777 730 795 746
rect 811 730 829 746
rect 845 730 863 746
rect 879 730 897 746
rect 913 730 931 746
rect 947 730 965 746
rect 981 730 999 746
rect 1015 730 1033 746
rect 1049 730 1067 746
rect 1083 730 1101 746
rect 1117 730 1135 746
rect 1151 730 1169 746
rect 1185 730 1203 746
rect 1219 730 1237 746
rect 1253 730 1271 746
rect 1287 730 1305 746
rect 1321 730 1339 746
rect 1355 730 1373 746
rect 1389 730 1407 746
rect 1423 730 1441 746
rect 1457 730 1475 746
rect 1491 730 1509 746
rect 1525 730 1543 746
rect 1559 730 1577 746
rect 1593 730 1611 746
rect 1627 730 1645 746
rect 1661 730 1679 746
rect 1695 730 1713 746
rect 1729 730 1747 746
rect 1763 730 1781 746
rect 1797 730 1815 746
rect 1831 730 1849 746
rect 1865 730 1883 746
rect 1899 730 1917 746
rect 1933 730 1951 746
rect 1967 730 1985 746
rect 2001 730 2019 746
rect 2035 730 2053 746
rect 2069 730 2087 746
rect 2103 730 2121 746
rect 2137 730 2155 746
rect 2171 730 2189 746
rect 2205 730 2223 746
rect 2239 730 2257 746
rect 2273 730 2291 746
rect 2307 730 2325 746
rect 2341 730 2359 746
rect 2375 730 2393 746
rect 2409 730 2427 746
rect 2443 730 2461 746
rect 2477 730 2495 746
rect 2511 730 2529 746
rect 2545 730 2563 746
rect 2579 730 2597 746
rect 2613 730 2631 746
rect 2647 730 2665 746
rect 2681 730 2699 746
rect 2715 730 2733 746
rect 2749 730 2767 746
rect 2783 730 2801 746
rect 2817 730 2835 746
rect 2851 730 2869 746
rect 2885 730 2903 746
rect 2919 730 2937 746
rect 2953 730 2971 746
rect 2987 730 3005 746
rect 3021 730 3042 746
rect 264 712 3042 730
rect 264 696 285 712
rect 301 696 319 712
rect 335 696 353 712
rect 369 696 387 712
rect 403 696 421 712
rect 437 696 455 712
rect 471 696 489 712
rect 505 696 523 712
rect 539 696 557 712
rect 573 696 591 712
rect 607 696 625 712
rect 641 696 659 712
rect 675 696 693 712
rect 709 696 727 712
rect 743 696 761 712
rect 777 696 795 712
rect 811 696 829 712
rect 845 696 863 712
rect 879 696 897 712
rect 913 696 931 712
rect 947 696 965 712
rect 981 696 999 712
rect 1015 696 1033 712
rect 1049 696 1067 712
rect 1083 696 1101 712
rect 1117 696 1135 712
rect 1151 696 1169 712
rect 1185 696 1203 712
rect 1219 696 1237 712
rect 1253 696 1271 712
rect 1287 696 1305 712
rect 1321 696 1339 712
rect 1355 696 1373 712
rect 1389 696 1407 712
rect 1423 696 1441 712
rect 1457 696 1475 712
rect 1491 696 1509 712
rect 1525 696 1543 712
rect 1559 696 1577 712
rect 1593 696 1611 712
rect 1627 696 1645 712
rect 1661 696 1679 712
rect 1695 696 1713 712
rect 1729 696 1747 712
rect 1763 696 1781 712
rect 1797 696 1815 712
rect 1831 696 1849 712
rect 1865 696 1883 712
rect 1899 696 1917 712
rect 1933 696 1951 712
rect 1967 696 1985 712
rect 2001 696 2019 712
rect 2035 696 2053 712
rect 2069 696 2087 712
rect 2103 696 2121 712
rect 2137 696 2155 712
rect 2171 696 2189 712
rect 2205 696 2223 712
rect 2239 696 2257 712
rect 2273 696 2291 712
rect 2307 696 2325 712
rect 2341 696 2359 712
rect 2375 696 2393 712
rect 2409 696 2427 712
rect 2443 696 2461 712
rect 2477 696 2495 712
rect 2511 696 2529 712
rect 2545 696 2563 712
rect 2579 696 2597 712
rect 2613 696 2631 712
rect 2647 696 2665 712
rect 2681 696 2699 712
rect 2715 696 2733 712
rect 2749 696 2767 712
rect 2783 696 2801 712
rect 2817 696 2835 712
rect 2851 696 2869 712
rect 2885 696 2903 712
rect 2919 696 2937 712
rect 2953 696 2971 712
rect 2987 696 3005 712
rect 3021 696 3042 712
rect 264 675 3042 696
rect 264 330 3042 351
rect 264 314 285 330
rect 301 314 319 330
rect 335 314 353 330
rect 369 314 387 330
rect 403 314 421 330
rect 437 314 455 330
rect 471 314 489 330
rect 505 314 523 330
rect 539 314 557 330
rect 573 314 591 330
rect 607 314 625 330
rect 641 314 659 330
rect 675 314 693 330
rect 709 314 727 330
rect 743 314 761 330
rect 777 314 795 330
rect 811 314 829 330
rect 845 314 863 330
rect 879 314 897 330
rect 913 314 931 330
rect 947 314 965 330
rect 981 314 999 330
rect 1015 314 1033 330
rect 1049 314 1067 330
rect 1083 314 1101 330
rect 1117 314 1135 330
rect 1151 314 1169 330
rect 1185 314 1203 330
rect 1219 314 1237 330
rect 1253 314 1271 330
rect 1287 314 1305 330
rect 1321 314 1339 330
rect 1355 314 1373 330
rect 1389 314 1407 330
rect 1423 314 1441 330
rect 1457 314 1475 330
rect 1491 314 1509 330
rect 1525 314 1543 330
rect 1559 314 1577 330
rect 1593 314 1611 330
rect 1627 314 1645 330
rect 1661 314 1679 330
rect 1695 314 1713 330
rect 1729 314 1747 330
rect 1763 314 1781 330
rect 1797 314 1815 330
rect 1831 314 1849 330
rect 1865 314 1883 330
rect 1899 314 1917 330
rect 1933 314 1951 330
rect 1967 314 1985 330
rect 2001 314 2019 330
rect 2035 314 2053 330
rect 2069 314 2087 330
rect 2103 314 2121 330
rect 2137 314 2155 330
rect 2171 314 2189 330
rect 2205 314 2223 330
rect 2239 314 2257 330
rect 2273 314 2291 330
rect 2307 314 2325 330
rect 2341 314 2359 330
rect 2375 314 2393 330
rect 2409 314 2427 330
rect 2443 314 2461 330
rect 2477 314 2495 330
rect 2511 314 2529 330
rect 2545 314 2563 330
rect 2579 314 2597 330
rect 2613 314 2631 330
rect 2647 314 2665 330
rect 2681 314 2699 330
rect 2715 314 2733 330
rect 2749 314 2767 330
rect 2783 314 2801 330
rect 2817 314 2835 330
rect 2851 314 2869 330
rect 2885 314 2903 330
rect 2919 314 2937 330
rect 2953 314 2971 330
rect 2987 314 3005 330
rect 3021 314 3042 330
rect 264 296 3042 314
rect 264 280 285 296
rect 301 280 319 296
rect 335 280 353 296
rect 369 280 387 296
rect 403 280 421 296
rect 437 280 455 296
rect 471 280 489 296
rect 505 280 523 296
rect 539 280 557 296
rect 573 280 591 296
rect 607 280 625 296
rect 641 280 659 296
rect 675 280 693 296
rect 709 280 727 296
rect 743 280 761 296
rect 777 280 795 296
rect 811 280 829 296
rect 845 280 863 296
rect 879 280 897 296
rect 913 280 931 296
rect 947 280 965 296
rect 981 280 999 296
rect 1015 280 1033 296
rect 1049 280 1067 296
rect 1083 280 1101 296
rect 1117 280 1135 296
rect 1151 280 1169 296
rect 1185 280 1203 296
rect 1219 280 1237 296
rect 1253 280 1271 296
rect 1287 280 1305 296
rect 1321 280 1339 296
rect 1355 280 1373 296
rect 1389 280 1407 296
rect 1423 280 1441 296
rect 1457 280 1475 296
rect 1491 280 1509 296
rect 1525 280 1543 296
rect 1559 280 1577 296
rect 1593 280 1611 296
rect 1627 280 1645 296
rect 1661 280 1679 296
rect 1695 280 1713 296
rect 1729 280 1747 296
rect 1763 280 1781 296
rect 1797 280 1815 296
rect 1831 280 1849 296
rect 1865 280 1883 296
rect 1899 280 1917 296
rect 1933 280 1951 296
rect 1967 280 1985 296
rect 2001 280 2019 296
rect 2035 280 2053 296
rect 2069 280 2087 296
rect 2103 280 2121 296
rect 2137 280 2155 296
rect 2171 280 2189 296
rect 2205 280 2223 296
rect 2239 280 2257 296
rect 2273 280 2291 296
rect 2307 280 2325 296
rect 2341 280 2359 296
rect 2375 280 2393 296
rect 2409 280 2427 296
rect 2443 280 2461 296
rect 2477 280 2495 296
rect 2511 280 2529 296
rect 2545 280 2563 296
rect 2579 280 2597 296
rect 2613 280 2631 296
rect 2647 280 2665 296
rect 2681 280 2699 296
rect 2715 280 2733 296
rect 2749 280 2767 296
rect 2783 280 2801 296
rect 2817 280 2835 296
rect 2851 280 2869 296
rect 2885 280 2903 296
rect 2919 280 2937 296
rect 2953 280 2971 296
rect 2987 280 3005 296
rect 3021 280 3042 296
rect 264 262 3042 280
rect 264 246 285 262
rect 301 246 319 262
rect 335 246 353 262
rect 369 246 387 262
rect 403 246 421 262
rect 437 246 455 262
rect 471 246 489 262
rect 505 246 523 262
rect 539 246 557 262
rect 573 246 591 262
rect 607 246 625 262
rect 641 246 659 262
rect 675 246 693 262
rect 709 246 727 262
rect 743 246 761 262
rect 777 246 795 262
rect 811 246 829 262
rect 845 246 863 262
rect 879 246 897 262
rect 913 246 931 262
rect 947 246 965 262
rect 981 246 999 262
rect 1015 246 1033 262
rect 1049 246 1067 262
rect 1083 246 1101 262
rect 1117 246 1135 262
rect 1151 246 1169 262
rect 1185 246 1203 262
rect 1219 246 1237 262
rect 1253 246 1271 262
rect 1287 246 1305 262
rect 1321 246 1339 262
rect 1355 246 1373 262
rect 1389 246 1407 262
rect 1423 246 1441 262
rect 1457 246 1475 262
rect 1491 246 1509 262
rect 1525 246 1543 262
rect 1559 246 1577 262
rect 1593 246 1611 262
rect 1627 246 1645 262
rect 1661 246 1679 262
rect 1695 246 1713 262
rect 1729 246 1747 262
rect 1763 246 1781 262
rect 1797 246 1815 262
rect 1831 246 1849 262
rect 1865 246 1883 262
rect 1899 246 1917 262
rect 1933 246 1951 262
rect 1967 246 1985 262
rect 2001 246 2019 262
rect 2035 246 2053 262
rect 2069 246 2087 262
rect 2103 246 2121 262
rect 2137 246 2155 262
rect 2171 246 2189 262
rect 2205 246 2223 262
rect 2239 246 2257 262
rect 2273 246 2291 262
rect 2307 246 2325 262
rect 2341 246 2359 262
rect 2375 246 2393 262
rect 2409 246 2427 262
rect 2443 246 2461 262
rect 2477 246 2495 262
rect 2511 246 2529 262
rect 2545 246 2563 262
rect 2579 246 2597 262
rect 2613 246 2631 262
rect 2647 246 2665 262
rect 2681 246 2699 262
rect 2715 246 2733 262
rect 2749 246 2767 262
rect 2783 246 2801 262
rect 2817 246 2835 262
rect 2851 246 2869 262
rect 2885 246 2903 262
rect 2919 246 2937 262
rect 2953 246 2971 262
rect 2987 246 3005 262
rect 3021 246 3042 262
rect 264 225 3042 246
<< pdiodecont >>
rect 285 764 301 780
rect 319 764 335 780
rect 353 764 369 780
rect 387 764 403 780
rect 421 764 437 780
rect 455 764 471 780
rect 489 764 505 780
rect 523 764 539 780
rect 557 764 573 780
rect 591 764 607 780
rect 625 764 641 780
rect 659 764 675 780
rect 693 764 709 780
rect 727 764 743 780
rect 761 764 777 780
rect 795 764 811 780
rect 829 764 845 780
rect 863 764 879 780
rect 897 764 913 780
rect 931 764 947 780
rect 965 764 981 780
rect 999 764 1015 780
rect 1033 764 1049 780
rect 1067 764 1083 780
rect 1101 764 1117 780
rect 1135 764 1151 780
rect 1169 764 1185 780
rect 1203 764 1219 780
rect 1237 764 1253 780
rect 1271 764 1287 780
rect 1305 764 1321 780
rect 1339 764 1355 780
rect 1373 764 1389 780
rect 1407 764 1423 780
rect 1441 764 1457 780
rect 1475 764 1491 780
rect 1509 764 1525 780
rect 1543 764 1559 780
rect 1577 764 1593 780
rect 1611 764 1627 780
rect 1645 764 1661 780
rect 1679 764 1695 780
rect 1713 764 1729 780
rect 1747 764 1763 780
rect 1781 764 1797 780
rect 1815 764 1831 780
rect 1849 764 1865 780
rect 1883 764 1899 780
rect 1917 764 1933 780
rect 1951 764 1967 780
rect 1985 764 2001 780
rect 2019 764 2035 780
rect 2053 764 2069 780
rect 2087 764 2103 780
rect 2121 764 2137 780
rect 2155 764 2171 780
rect 2189 764 2205 780
rect 2223 764 2239 780
rect 2257 764 2273 780
rect 2291 764 2307 780
rect 2325 764 2341 780
rect 2359 764 2375 780
rect 2393 764 2409 780
rect 2427 764 2443 780
rect 2461 764 2477 780
rect 2495 764 2511 780
rect 2529 764 2545 780
rect 2563 764 2579 780
rect 2597 764 2613 780
rect 2631 764 2647 780
rect 2665 764 2681 780
rect 2699 764 2715 780
rect 2733 764 2749 780
rect 2767 764 2783 780
rect 2801 764 2817 780
rect 2835 764 2851 780
rect 2869 764 2885 780
rect 2903 764 2919 780
rect 2937 764 2953 780
rect 2971 764 2987 780
rect 3005 764 3021 780
rect 285 730 301 746
rect 319 730 335 746
rect 353 730 369 746
rect 387 730 403 746
rect 421 730 437 746
rect 455 730 471 746
rect 489 730 505 746
rect 523 730 539 746
rect 557 730 573 746
rect 591 730 607 746
rect 625 730 641 746
rect 659 730 675 746
rect 693 730 709 746
rect 727 730 743 746
rect 761 730 777 746
rect 795 730 811 746
rect 829 730 845 746
rect 863 730 879 746
rect 897 730 913 746
rect 931 730 947 746
rect 965 730 981 746
rect 999 730 1015 746
rect 1033 730 1049 746
rect 1067 730 1083 746
rect 1101 730 1117 746
rect 1135 730 1151 746
rect 1169 730 1185 746
rect 1203 730 1219 746
rect 1237 730 1253 746
rect 1271 730 1287 746
rect 1305 730 1321 746
rect 1339 730 1355 746
rect 1373 730 1389 746
rect 1407 730 1423 746
rect 1441 730 1457 746
rect 1475 730 1491 746
rect 1509 730 1525 746
rect 1543 730 1559 746
rect 1577 730 1593 746
rect 1611 730 1627 746
rect 1645 730 1661 746
rect 1679 730 1695 746
rect 1713 730 1729 746
rect 1747 730 1763 746
rect 1781 730 1797 746
rect 1815 730 1831 746
rect 1849 730 1865 746
rect 1883 730 1899 746
rect 1917 730 1933 746
rect 1951 730 1967 746
rect 1985 730 2001 746
rect 2019 730 2035 746
rect 2053 730 2069 746
rect 2087 730 2103 746
rect 2121 730 2137 746
rect 2155 730 2171 746
rect 2189 730 2205 746
rect 2223 730 2239 746
rect 2257 730 2273 746
rect 2291 730 2307 746
rect 2325 730 2341 746
rect 2359 730 2375 746
rect 2393 730 2409 746
rect 2427 730 2443 746
rect 2461 730 2477 746
rect 2495 730 2511 746
rect 2529 730 2545 746
rect 2563 730 2579 746
rect 2597 730 2613 746
rect 2631 730 2647 746
rect 2665 730 2681 746
rect 2699 730 2715 746
rect 2733 730 2749 746
rect 2767 730 2783 746
rect 2801 730 2817 746
rect 2835 730 2851 746
rect 2869 730 2885 746
rect 2903 730 2919 746
rect 2937 730 2953 746
rect 2971 730 2987 746
rect 3005 730 3021 746
rect 285 696 301 712
rect 319 696 335 712
rect 353 696 369 712
rect 387 696 403 712
rect 421 696 437 712
rect 455 696 471 712
rect 489 696 505 712
rect 523 696 539 712
rect 557 696 573 712
rect 591 696 607 712
rect 625 696 641 712
rect 659 696 675 712
rect 693 696 709 712
rect 727 696 743 712
rect 761 696 777 712
rect 795 696 811 712
rect 829 696 845 712
rect 863 696 879 712
rect 897 696 913 712
rect 931 696 947 712
rect 965 696 981 712
rect 999 696 1015 712
rect 1033 696 1049 712
rect 1067 696 1083 712
rect 1101 696 1117 712
rect 1135 696 1151 712
rect 1169 696 1185 712
rect 1203 696 1219 712
rect 1237 696 1253 712
rect 1271 696 1287 712
rect 1305 696 1321 712
rect 1339 696 1355 712
rect 1373 696 1389 712
rect 1407 696 1423 712
rect 1441 696 1457 712
rect 1475 696 1491 712
rect 1509 696 1525 712
rect 1543 696 1559 712
rect 1577 696 1593 712
rect 1611 696 1627 712
rect 1645 696 1661 712
rect 1679 696 1695 712
rect 1713 696 1729 712
rect 1747 696 1763 712
rect 1781 696 1797 712
rect 1815 696 1831 712
rect 1849 696 1865 712
rect 1883 696 1899 712
rect 1917 696 1933 712
rect 1951 696 1967 712
rect 1985 696 2001 712
rect 2019 696 2035 712
rect 2053 696 2069 712
rect 2087 696 2103 712
rect 2121 696 2137 712
rect 2155 696 2171 712
rect 2189 696 2205 712
rect 2223 696 2239 712
rect 2257 696 2273 712
rect 2291 696 2307 712
rect 2325 696 2341 712
rect 2359 696 2375 712
rect 2393 696 2409 712
rect 2427 696 2443 712
rect 2461 696 2477 712
rect 2495 696 2511 712
rect 2529 696 2545 712
rect 2563 696 2579 712
rect 2597 696 2613 712
rect 2631 696 2647 712
rect 2665 696 2681 712
rect 2699 696 2715 712
rect 2733 696 2749 712
rect 2767 696 2783 712
rect 2801 696 2817 712
rect 2835 696 2851 712
rect 2869 696 2885 712
rect 2903 696 2919 712
rect 2937 696 2953 712
rect 2971 696 2987 712
rect 3005 696 3021 712
rect 285 314 301 330
rect 319 314 335 330
rect 353 314 369 330
rect 387 314 403 330
rect 421 314 437 330
rect 455 314 471 330
rect 489 314 505 330
rect 523 314 539 330
rect 557 314 573 330
rect 591 314 607 330
rect 625 314 641 330
rect 659 314 675 330
rect 693 314 709 330
rect 727 314 743 330
rect 761 314 777 330
rect 795 314 811 330
rect 829 314 845 330
rect 863 314 879 330
rect 897 314 913 330
rect 931 314 947 330
rect 965 314 981 330
rect 999 314 1015 330
rect 1033 314 1049 330
rect 1067 314 1083 330
rect 1101 314 1117 330
rect 1135 314 1151 330
rect 1169 314 1185 330
rect 1203 314 1219 330
rect 1237 314 1253 330
rect 1271 314 1287 330
rect 1305 314 1321 330
rect 1339 314 1355 330
rect 1373 314 1389 330
rect 1407 314 1423 330
rect 1441 314 1457 330
rect 1475 314 1491 330
rect 1509 314 1525 330
rect 1543 314 1559 330
rect 1577 314 1593 330
rect 1611 314 1627 330
rect 1645 314 1661 330
rect 1679 314 1695 330
rect 1713 314 1729 330
rect 1747 314 1763 330
rect 1781 314 1797 330
rect 1815 314 1831 330
rect 1849 314 1865 330
rect 1883 314 1899 330
rect 1917 314 1933 330
rect 1951 314 1967 330
rect 1985 314 2001 330
rect 2019 314 2035 330
rect 2053 314 2069 330
rect 2087 314 2103 330
rect 2121 314 2137 330
rect 2155 314 2171 330
rect 2189 314 2205 330
rect 2223 314 2239 330
rect 2257 314 2273 330
rect 2291 314 2307 330
rect 2325 314 2341 330
rect 2359 314 2375 330
rect 2393 314 2409 330
rect 2427 314 2443 330
rect 2461 314 2477 330
rect 2495 314 2511 330
rect 2529 314 2545 330
rect 2563 314 2579 330
rect 2597 314 2613 330
rect 2631 314 2647 330
rect 2665 314 2681 330
rect 2699 314 2715 330
rect 2733 314 2749 330
rect 2767 314 2783 330
rect 2801 314 2817 330
rect 2835 314 2851 330
rect 2869 314 2885 330
rect 2903 314 2919 330
rect 2937 314 2953 330
rect 2971 314 2987 330
rect 3005 314 3021 330
rect 285 280 301 296
rect 319 280 335 296
rect 353 280 369 296
rect 387 280 403 296
rect 421 280 437 296
rect 455 280 471 296
rect 489 280 505 296
rect 523 280 539 296
rect 557 280 573 296
rect 591 280 607 296
rect 625 280 641 296
rect 659 280 675 296
rect 693 280 709 296
rect 727 280 743 296
rect 761 280 777 296
rect 795 280 811 296
rect 829 280 845 296
rect 863 280 879 296
rect 897 280 913 296
rect 931 280 947 296
rect 965 280 981 296
rect 999 280 1015 296
rect 1033 280 1049 296
rect 1067 280 1083 296
rect 1101 280 1117 296
rect 1135 280 1151 296
rect 1169 280 1185 296
rect 1203 280 1219 296
rect 1237 280 1253 296
rect 1271 280 1287 296
rect 1305 280 1321 296
rect 1339 280 1355 296
rect 1373 280 1389 296
rect 1407 280 1423 296
rect 1441 280 1457 296
rect 1475 280 1491 296
rect 1509 280 1525 296
rect 1543 280 1559 296
rect 1577 280 1593 296
rect 1611 280 1627 296
rect 1645 280 1661 296
rect 1679 280 1695 296
rect 1713 280 1729 296
rect 1747 280 1763 296
rect 1781 280 1797 296
rect 1815 280 1831 296
rect 1849 280 1865 296
rect 1883 280 1899 296
rect 1917 280 1933 296
rect 1951 280 1967 296
rect 1985 280 2001 296
rect 2019 280 2035 296
rect 2053 280 2069 296
rect 2087 280 2103 296
rect 2121 280 2137 296
rect 2155 280 2171 296
rect 2189 280 2205 296
rect 2223 280 2239 296
rect 2257 280 2273 296
rect 2291 280 2307 296
rect 2325 280 2341 296
rect 2359 280 2375 296
rect 2393 280 2409 296
rect 2427 280 2443 296
rect 2461 280 2477 296
rect 2495 280 2511 296
rect 2529 280 2545 296
rect 2563 280 2579 296
rect 2597 280 2613 296
rect 2631 280 2647 296
rect 2665 280 2681 296
rect 2699 280 2715 296
rect 2733 280 2749 296
rect 2767 280 2783 296
rect 2801 280 2817 296
rect 2835 280 2851 296
rect 2869 280 2885 296
rect 2903 280 2919 296
rect 2937 280 2953 296
rect 2971 280 2987 296
rect 3005 280 3021 296
rect 285 246 301 262
rect 319 246 335 262
rect 353 246 369 262
rect 387 246 403 262
rect 421 246 437 262
rect 455 246 471 262
rect 489 246 505 262
rect 523 246 539 262
rect 557 246 573 262
rect 591 246 607 262
rect 625 246 641 262
rect 659 246 675 262
rect 693 246 709 262
rect 727 246 743 262
rect 761 246 777 262
rect 795 246 811 262
rect 829 246 845 262
rect 863 246 879 262
rect 897 246 913 262
rect 931 246 947 262
rect 965 246 981 262
rect 999 246 1015 262
rect 1033 246 1049 262
rect 1067 246 1083 262
rect 1101 246 1117 262
rect 1135 246 1151 262
rect 1169 246 1185 262
rect 1203 246 1219 262
rect 1237 246 1253 262
rect 1271 246 1287 262
rect 1305 246 1321 262
rect 1339 246 1355 262
rect 1373 246 1389 262
rect 1407 246 1423 262
rect 1441 246 1457 262
rect 1475 246 1491 262
rect 1509 246 1525 262
rect 1543 246 1559 262
rect 1577 246 1593 262
rect 1611 246 1627 262
rect 1645 246 1661 262
rect 1679 246 1695 262
rect 1713 246 1729 262
rect 1747 246 1763 262
rect 1781 246 1797 262
rect 1815 246 1831 262
rect 1849 246 1865 262
rect 1883 246 1899 262
rect 1917 246 1933 262
rect 1951 246 1967 262
rect 1985 246 2001 262
rect 2019 246 2035 262
rect 2053 246 2069 262
rect 2087 246 2103 262
rect 2121 246 2137 262
rect 2155 246 2171 262
rect 2189 246 2205 262
rect 2223 246 2239 262
rect 2257 246 2273 262
rect 2291 246 2307 262
rect 2325 246 2341 262
rect 2359 246 2375 262
rect 2393 246 2409 262
rect 2427 246 2443 262
rect 2461 246 2477 262
rect 2495 246 2511 262
rect 2529 246 2545 262
rect 2563 246 2579 262
rect 2597 246 2613 262
rect 2631 246 2647 262
rect 2665 246 2681 262
rect 2699 246 2715 262
rect 2733 246 2749 262
rect 2767 246 2783 262
rect 2801 246 2817 262
rect 2835 246 2851 262
rect 2869 246 2885 262
rect 2903 246 2919 262
rect 2937 246 2953 262
rect 2971 246 2987 262
rect 3005 246 3021 262
<< metal1 >>
rect -166 1183 3472 1192
rect -166 1167 -157 1183
rect -141 1167 -123 1183
rect -107 1167 -89 1183
rect -73 1167 -55 1183
rect -39 1167 -21 1183
rect -5 1167 13 1183
rect 29 1167 47 1183
rect 63 1167 81 1183
rect 97 1167 115 1183
rect 131 1167 149 1183
rect 165 1167 183 1183
rect 199 1167 217 1183
rect 233 1167 251 1183
rect 267 1167 285 1183
rect 301 1167 319 1183
rect 335 1167 353 1183
rect 369 1167 387 1183
rect 403 1167 421 1183
rect 437 1167 455 1183
rect 471 1167 489 1183
rect 505 1167 523 1183
rect 539 1167 557 1183
rect 573 1167 591 1183
rect 607 1167 625 1183
rect 641 1167 659 1183
rect 675 1167 693 1183
rect 709 1167 727 1183
rect 743 1167 761 1183
rect 777 1167 795 1183
rect 811 1167 829 1183
rect 845 1167 863 1183
rect 879 1167 897 1183
rect 913 1167 931 1183
rect 947 1167 965 1183
rect 981 1167 999 1183
rect 1015 1167 1033 1183
rect 1049 1167 1067 1183
rect 1083 1167 1101 1183
rect 1117 1167 1135 1183
rect 1151 1167 1169 1183
rect 1185 1167 1203 1183
rect 1219 1167 1237 1183
rect 1253 1167 1271 1183
rect 1287 1167 1305 1183
rect 1321 1167 1339 1183
rect 1355 1167 1373 1183
rect 1389 1167 1407 1183
rect 1423 1167 1441 1183
rect 1457 1167 1475 1183
rect 1491 1167 1509 1183
rect 1525 1167 1543 1183
rect 1559 1167 1577 1183
rect 1593 1167 1611 1183
rect 1627 1167 1645 1183
rect 1661 1167 1679 1183
rect 1695 1167 1713 1183
rect 1729 1167 1747 1183
rect 1763 1167 1781 1183
rect 1797 1167 1815 1183
rect 1831 1167 1849 1183
rect 1865 1167 1883 1183
rect 1899 1167 1917 1183
rect 1933 1167 1951 1183
rect 1967 1167 1985 1183
rect 2001 1167 2019 1183
rect 2035 1167 2053 1183
rect 2069 1167 2087 1183
rect 2103 1167 2121 1183
rect 2137 1167 2155 1183
rect 2171 1167 2189 1183
rect 2205 1167 2223 1183
rect 2239 1167 2257 1183
rect 2273 1167 2291 1183
rect 2307 1167 2325 1183
rect 2341 1167 2359 1183
rect 2375 1167 2393 1183
rect 2409 1167 2427 1183
rect 2443 1167 2461 1183
rect 2477 1167 2495 1183
rect 2511 1167 2529 1183
rect 2545 1167 2563 1183
rect 2579 1167 2597 1183
rect 2613 1167 2631 1183
rect 2647 1167 2665 1183
rect 2681 1167 2699 1183
rect 2715 1167 2733 1183
rect 2749 1167 2767 1183
rect 2783 1167 2801 1183
rect 2817 1167 2835 1183
rect 2851 1167 2869 1183
rect 2885 1167 2903 1183
rect 2919 1167 2937 1183
rect 2953 1167 2971 1183
rect 2987 1167 3005 1183
rect 3021 1167 3039 1183
rect 3055 1167 3073 1183
rect 3089 1167 3107 1183
rect 3123 1167 3141 1183
rect 3157 1167 3175 1183
rect 3191 1167 3209 1183
rect 3225 1167 3243 1183
rect 3259 1167 3277 1183
rect 3293 1167 3311 1183
rect 3327 1167 3345 1183
rect 3361 1167 3379 1183
rect 3395 1167 3413 1183
rect 3429 1167 3447 1183
rect 3463 1167 3472 1183
rect -166 1158 3472 1167
rect -166 1133 -132 1158
rect -166 1117 -157 1133
rect -141 1117 -132 1133
rect -166 1099 -132 1117
rect -166 1083 -157 1099
rect -141 1083 -132 1099
rect -166 1065 -132 1083
rect -166 1049 -157 1065
rect -141 1049 -132 1065
rect -166 1031 -132 1049
rect -166 1015 -157 1031
rect -141 1015 -132 1031
rect 3438 1133 3472 1158
rect 3438 1117 3447 1133
rect 3463 1117 3472 1133
rect 3438 1099 3472 1117
rect 3438 1083 3447 1099
rect 3463 1083 3472 1099
rect 3438 1065 3472 1083
rect 3438 1049 3447 1065
rect 3463 1049 3472 1065
rect 3438 1031 3472 1049
rect -166 997 -132 1015
rect -166 981 -157 997
rect -141 981 -132 997
rect -166 963 -132 981
rect -166 947 -157 963
rect -141 947 -132 963
rect -166 929 -132 947
rect -166 913 -157 929
rect -141 913 -132 929
rect -166 895 -132 913
rect -166 879 -157 895
rect -141 879 -132 895
rect -166 861 -132 879
rect -166 845 -157 861
rect -141 845 -132 861
rect -166 827 -132 845
rect -166 811 -157 827
rect -141 811 -132 827
rect -166 793 -132 811
rect -166 777 -157 793
rect -141 777 -132 793
rect -166 759 -132 777
rect -166 743 -157 759
rect -141 743 -132 759
rect -166 725 -132 743
rect -166 709 -157 725
rect -141 709 -132 725
rect -166 691 -132 709
rect -166 675 -157 691
rect -141 675 -132 691
rect -166 657 -132 675
rect -166 641 -157 657
rect -141 641 -132 657
rect -166 623 -132 641
rect -166 607 -157 623
rect -141 607 -132 623
rect -166 589 -132 607
rect -166 573 -157 589
rect -141 573 -132 589
rect -166 555 -132 573
rect -166 539 -157 555
rect -141 539 -132 555
rect -166 521 -132 539
rect -166 505 -157 521
rect -141 505 -132 521
rect -166 487 -132 505
rect -166 471 -157 487
rect -141 471 -132 487
rect -166 453 -132 471
rect -166 437 -157 453
rect -141 437 -132 453
rect -166 419 -132 437
rect -166 403 -157 419
rect -141 403 -132 419
rect -166 385 -132 403
rect -166 369 -157 385
rect -141 369 -132 385
rect -166 351 -132 369
rect -166 335 -157 351
rect -141 335 -132 351
rect -166 317 -132 335
rect -166 301 -157 317
rect -141 301 -132 317
rect -166 283 -132 301
rect -166 267 -157 283
rect -141 267 -132 283
rect -166 249 -132 267
rect -166 233 -157 249
rect -141 233 -132 249
rect -166 215 -132 233
rect -166 199 -157 215
rect -141 199 -132 215
rect -166 181 -132 199
rect -166 165 -157 181
rect -141 165 -132 181
rect -166 147 -132 165
rect -166 131 -157 147
rect -141 131 -132 147
rect -166 113 -132 131
rect -166 97 -157 113
rect -141 97 -132 113
rect -166 79 -132 97
rect -166 63 -157 79
rect -141 63 -132 79
rect -166 45 -132 63
rect -166 29 -157 45
rect -141 29 -132 45
rect -166 11 -132 29
rect -166 -5 -157 11
rect -141 -5 -132 11
rect 0 1014 3306 1026
rect 0 998 21 1014
rect 37 998 55 1014
rect 71 998 89 1014
rect 105 1005 3201 1014
rect 105 998 149 1005
rect 0 989 149 998
rect 165 989 183 1005
rect 199 989 217 1005
rect 233 989 251 1005
rect 267 989 285 1005
rect 301 989 319 1005
rect 335 989 353 1005
rect 369 989 387 1005
rect 403 989 421 1005
rect 437 989 455 1005
rect 471 989 489 1005
rect 505 989 523 1005
rect 539 989 557 1005
rect 573 989 591 1005
rect 607 989 625 1005
rect 641 989 659 1005
rect 675 989 693 1005
rect 709 989 727 1005
rect 743 989 761 1005
rect 777 989 795 1005
rect 811 989 829 1005
rect 845 989 863 1005
rect 879 989 897 1005
rect 913 989 931 1005
rect 947 989 965 1005
rect 981 989 999 1005
rect 1015 989 1033 1005
rect 1049 989 1067 1005
rect 1083 989 1101 1005
rect 1117 989 1135 1005
rect 1151 989 1169 1005
rect 1185 989 1203 1005
rect 1219 989 1237 1005
rect 1253 989 1271 1005
rect 1287 989 1305 1005
rect 1321 989 1339 1005
rect 1355 989 1373 1005
rect 1389 989 1407 1005
rect 1423 989 1441 1005
rect 1457 989 1475 1005
rect 1491 989 1509 1005
rect 1525 989 1543 1005
rect 1559 989 1577 1005
rect 1593 989 1611 1005
rect 1627 989 1645 1005
rect 1661 989 1679 1005
rect 1695 989 1713 1005
rect 1729 989 1747 1005
rect 1763 989 1781 1005
rect 1797 989 1815 1005
rect 1831 989 1849 1005
rect 1865 989 1883 1005
rect 1899 989 1917 1005
rect 1933 989 1951 1005
rect 1967 989 1985 1005
rect 2001 989 2019 1005
rect 2035 989 2053 1005
rect 2069 989 2087 1005
rect 2103 989 2121 1005
rect 2137 989 2155 1005
rect 2171 989 2189 1005
rect 2205 989 2223 1005
rect 2239 989 2257 1005
rect 2273 989 2291 1005
rect 2307 989 2325 1005
rect 2341 989 2359 1005
rect 2375 989 2393 1005
rect 2409 989 2427 1005
rect 2443 989 2461 1005
rect 2477 989 2495 1005
rect 2511 989 2529 1005
rect 2545 989 2563 1005
rect 2579 989 2597 1005
rect 2613 989 2631 1005
rect 2647 989 2665 1005
rect 2681 989 2699 1005
rect 2715 989 2733 1005
rect 2749 989 2767 1005
rect 2783 989 2801 1005
rect 2817 989 2835 1005
rect 2851 989 2869 1005
rect 2885 989 2903 1005
rect 2919 989 2937 1005
rect 2953 989 2971 1005
rect 2987 989 3005 1005
rect 3021 989 3039 1005
rect 3055 989 3073 1005
rect 3089 989 3107 1005
rect 3123 989 3141 1005
rect 3157 998 3201 1005
rect 3217 998 3235 1014
rect 3251 998 3269 1014
rect 3285 998 3306 1014
rect 3157 989 3306 998
rect 0 980 3306 989
rect 0 964 21 980
rect 37 964 55 980
rect 71 964 89 980
rect 105 971 3201 980
rect 105 964 149 971
rect 0 955 149 964
rect 165 955 183 971
rect 199 955 217 971
rect 233 955 251 971
rect 267 955 285 971
rect 301 955 319 971
rect 335 955 353 971
rect 369 955 387 971
rect 403 955 421 971
rect 437 955 455 971
rect 471 955 489 971
rect 505 955 523 971
rect 539 955 557 971
rect 573 955 591 971
rect 607 955 625 971
rect 641 955 659 971
rect 675 955 693 971
rect 709 955 727 971
rect 743 955 761 971
rect 777 955 795 971
rect 811 955 829 971
rect 845 955 863 971
rect 879 955 897 971
rect 913 955 931 971
rect 947 955 965 971
rect 981 955 999 971
rect 1015 955 1033 971
rect 1049 955 1067 971
rect 1083 955 1101 971
rect 1117 955 1135 971
rect 1151 955 1169 971
rect 1185 955 1203 971
rect 1219 955 1237 971
rect 1253 955 1271 971
rect 1287 955 1305 971
rect 1321 955 1339 971
rect 1355 955 1373 971
rect 1389 955 1407 971
rect 1423 955 1441 971
rect 1457 955 1475 971
rect 1491 955 1509 971
rect 1525 955 1543 971
rect 1559 955 1577 971
rect 1593 955 1611 971
rect 1627 955 1645 971
rect 1661 955 1679 971
rect 1695 955 1713 971
rect 1729 955 1747 971
rect 1763 955 1781 971
rect 1797 955 1815 971
rect 1831 955 1849 971
rect 1865 955 1883 971
rect 1899 955 1917 971
rect 1933 955 1951 971
rect 1967 955 1985 971
rect 2001 955 2019 971
rect 2035 955 2053 971
rect 2069 955 2087 971
rect 2103 955 2121 971
rect 2137 955 2155 971
rect 2171 955 2189 971
rect 2205 955 2223 971
rect 2239 955 2257 971
rect 2273 955 2291 971
rect 2307 955 2325 971
rect 2341 955 2359 971
rect 2375 955 2393 971
rect 2409 955 2427 971
rect 2443 955 2461 971
rect 2477 955 2495 971
rect 2511 955 2529 971
rect 2545 955 2563 971
rect 2579 955 2597 971
rect 2613 955 2631 971
rect 2647 955 2665 971
rect 2681 955 2699 971
rect 2715 955 2733 971
rect 2749 955 2767 971
rect 2783 955 2801 971
rect 2817 955 2835 971
rect 2851 955 2869 971
rect 2885 955 2903 971
rect 2919 955 2937 971
rect 2953 955 2971 971
rect 2987 955 3005 971
rect 3021 955 3039 971
rect 3055 955 3073 971
rect 3089 955 3107 971
rect 3123 955 3141 971
rect 3157 964 3201 971
rect 3217 964 3235 980
rect 3251 964 3269 980
rect 3285 964 3306 980
rect 3157 955 3306 964
rect 0 946 3306 955
rect 0 930 21 946
rect 37 930 55 946
rect 71 930 89 946
rect 105 937 3201 946
rect 105 930 149 937
rect 0 921 149 930
rect 165 921 183 937
rect 199 921 217 937
rect 233 921 251 937
rect 267 921 285 937
rect 301 921 319 937
rect 335 921 353 937
rect 369 921 387 937
rect 403 921 421 937
rect 437 921 455 937
rect 471 921 489 937
rect 505 921 523 937
rect 539 921 557 937
rect 573 921 591 937
rect 607 921 625 937
rect 641 921 659 937
rect 675 921 693 937
rect 709 921 727 937
rect 743 921 761 937
rect 777 921 795 937
rect 811 921 829 937
rect 845 921 863 937
rect 879 921 897 937
rect 913 921 931 937
rect 947 921 965 937
rect 981 921 999 937
rect 1015 921 1033 937
rect 1049 921 1067 937
rect 1083 921 1101 937
rect 1117 921 1135 937
rect 1151 921 1169 937
rect 1185 921 1203 937
rect 1219 921 1237 937
rect 1253 921 1271 937
rect 1287 921 1305 937
rect 1321 921 1339 937
rect 1355 921 1373 937
rect 1389 921 1407 937
rect 1423 921 1441 937
rect 1457 921 1475 937
rect 1491 921 1509 937
rect 1525 921 1543 937
rect 1559 921 1577 937
rect 1593 921 1611 937
rect 1627 921 1645 937
rect 1661 921 1679 937
rect 1695 921 1713 937
rect 1729 921 1747 937
rect 1763 921 1781 937
rect 1797 921 1815 937
rect 1831 921 1849 937
rect 1865 921 1883 937
rect 1899 921 1917 937
rect 1933 921 1951 937
rect 1967 921 1985 937
rect 2001 921 2019 937
rect 2035 921 2053 937
rect 2069 921 2087 937
rect 2103 921 2121 937
rect 2137 921 2155 937
rect 2171 921 2189 937
rect 2205 921 2223 937
rect 2239 921 2257 937
rect 2273 921 2291 937
rect 2307 921 2325 937
rect 2341 921 2359 937
rect 2375 921 2393 937
rect 2409 921 2427 937
rect 2443 921 2461 937
rect 2477 921 2495 937
rect 2511 921 2529 937
rect 2545 921 2563 937
rect 2579 921 2597 937
rect 2613 921 2631 937
rect 2647 921 2665 937
rect 2681 921 2699 937
rect 2715 921 2733 937
rect 2749 921 2767 937
rect 2783 921 2801 937
rect 2817 921 2835 937
rect 2851 921 2869 937
rect 2885 921 2903 937
rect 2919 921 2937 937
rect 2953 921 2971 937
rect 2987 921 3005 937
rect 3021 921 3039 937
rect 3055 921 3073 937
rect 3089 921 3107 937
rect 3123 921 3141 937
rect 3157 930 3201 937
rect 3217 930 3235 946
rect 3251 930 3269 946
rect 3285 930 3306 946
rect 3157 921 3306 930
rect 0 912 3306 921
rect 0 896 21 912
rect 37 896 55 912
rect 71 896 89 912
rect 105 900 3201 912
rect 105 896 126 900
rect 0 878 126 896
rect 0 862 21 878
rect 37 862 55 878
rect 71 862 89 878
rect 105 862 126 878
rect 0 844 126 862
rect 0 828 21 844
rect 37 828 55 844
rect 71 828 89 844
rect 105 828 126 844
rect 0 810 126 828
rect 0 794 21 810
rect 37 794 55 810
rect 71 794 89 810
rect 105 794 126 810
rect 3180 896 3201 900
rect 3217 896 3235 912
rect 3251 896 3269 912
rect 3285 896 3306 912
rect 3180 878 3306 896
rect 3180 862 3201 878
rect 3217 862 3235 878
rect 3251 862 3269 878
rect 3285 862 3306 878
rect 3180 844 3306 862
rect 3180 828 3201 844
rect 3217 828 3235 844
rect 3251 828 3269 844
rect 3285 828 3306 844
rect 3180 810 3306 828
rect 0 776 126 794
rect 0 760 21 776
rect 37 760 55 776
rect 71 760 89 776
rect 105 760 126 776
rect 0 742 126 760
rect 0 726 21 742
rect 37 726 55 742
rect 71 726 89 742
rect 105 726 126 742
rect 0 708 126 726
rect 0 692 21 708
rect 37 692 55 708
rect 71 692 89 708
rect 105 692 126 708
rect 0 674 126 692
rect 264 780 3042 801
rect 264 764 285 780
rect 301 764 319 780
rect 335 764 353 780
rect 369 764 387 780
rect 403 764 421 780
rect 437 764 455 780
rect 471 764 489 780
rect 505 764 523 780
rect 539 764 557 780
rect 573 764 591 780
rect 607 764 625 780
rect 641 764 659 780
rect 675 764 693 780
rect 709 764 727 780
rect 743 764 761 780
rect 777 764 795 780
rect 811 764 829 780
rect 845 764 863 780
rect 879 764 897 780
rect 913 764 931 780
rect 947 764 965 780
rect 981 764 999 780
rect 1015 764 1033 780
rect 1049 764 1067 780
rect 1083 764 1101 780
rect 1117 764 1135 780
rect 1151 764 1169 780
rect 1185 764 1203 780
rect 1219 764 1237 780
rect 1253 764 1271 780
rect 1287 764 1305 780
rect 1321 764 1339 780
rect 1355 764 1373 780
rect 1389 764 1407 780
rect 1423 764 1441 780
rect 1457 764 1475 780
rect 1491 764 1509 780
rect 1525 764 1543 780
rect 1559 764 1577 780
rect 1593 764 1611 780
rect 1627 764 1645 780
rect 1661 764 1679 780
rect 1695 764 1713 780
rect 1729 764 1747 780
rect 1763 764 1781 780
rect 1797 764 1815 780
rect 1831 764 1849 780
rect 1865 764 1883 780
rect 1899 764 1917 780
rect 1933 764 1951 780
rect 1967 764 1985 780
rect 2001 764 2019 780
rect 2035 764 2053 780
rect 2069 764 2087 780
rect 2103 764 2121 780
rect 2137 764 2155 780
rect 2171 764 2189 780
rect 2205 764 2223 780
rect 2239 764 2257 780
rect 2273 764 2291 780
rect 2307 764 2325 780
rect 2341 764 2359 780
rect 2375 764 2393 780
rect 2409 764 2427 780
rect 2443 764 2461 780
rect 2477 764 2495 780
rect 2511 764 2529 780
rect 2545 764 2563 780
rect 2579 764 2597 780
rect 2613 764 2631 780
rect 2647 764 2665 780
rect 2681 764 2699 780
rect 2715 764 2733 780
rect 2749 764 2767 780
rect 2783 764 2801 780
rect 2817 764 2835 780
rect 2851 764 2869 780
rect 2885 764 2903 780
rect 2919 764 2937 780
rect 2953 764 2971 780
rect 2987 764 3005 780
rect 3021 764 3042 780
rect 264 746 3042 764
rect 264 730 285 746
rect 301 730 319 746
rect 335 730 353 746
rect 369 730 387 746
rect 403 730 421 746
rect 437 730 455 746
rect 471 730 489 746
rect 505 730 523 746
rect 539 730 557 746
rect 573 730 591 746
rect 607 730 625 746
rect 641 730 659 746
rect 675 730 693 746
rect 709 730 727 746
rect 743 730 761 746
rect 777 730 795 746
rect 811 730 829 746
rect 845 730 863 746
rect 879 730 897 746
rect 913 730 931 746
rect 947 730 965 746
rect 981 730 999 746
rect 1015 730 1033 746
rect 1049 730 1067 746
rect 1083 730 1101 746
rect 1117 730 1135 746
rect 1151 730 1169 746
rect 1185 730 1203 746
rect 1219 730 1237 746
rect 1253 730 1271 746
rect 1287 730 1305 746
rect 1321 730 1339 746
rect 1355 730 1373 746
rect 1389 730 1407 746
rect 1423 730 1441 746
rect 1457 730 1475 746
rect 1491 730 1509 746
rect 1525 730 1543 746
rect 1559 730 1577 746
rect 1593 730 1611 746
rect 1627 730 1645 746
rect 1661 730 1679 746
rect 1695 730 1713 746
rect 1729 730 1747 746
rect 1763 730 1781 746
rect 1797 730 1815 746
rect 1831 730 1849 746
rect 1865 730 1883 746
rect 1899 730 1917 746
rect 1933 730 1951 746
rect 1967 730 1985 746
rect 2001 730 2019 746
rect 2035 730 2053 746
rect 2069 730 2087 746
rect 2103 730 2121 746
rect 2137 730 2155 746
rect 2171 730 2189 746
rect 2205 730 2223 746
rect 2239 730 2257 746
rect 2273 730 2291 746
rect 2307 730 2325 746
rect 2341 730 2359 746
rect 2375 730 2393 746
rect 2409 730 2427 746
rect 2443 730 2461 746
rect 2477 730 2495 746
rect 2511 730 2529 746
rect 2545 730 2563 746
rect 2579 730 2597 746
rect 2613 730 2631 746
rect 2647 730 2665 746
rect 2681 730 2699 746
rect 2715 730 2733 746
rect 2749 730 2767 746
rect 2783 730 2801 746
rect 2817 730 2835 746
rect 2851 730 2869 746
rect 2885 730 2903 746
rect 2919 730 2937 746
rect 2953 730 2971 746
rect 2987 730 3005 746
rect 3021 730 3042 746
rect 264 712 3042 730
rect 264 696 285 712
rect 301 696 319 712
rect 335 696 353 712
rect 369 696 387 712
rect 403 696 421 712
rect 437 696 455 712
rect 471 696 489 712
rect 505 696 523 712
rect 539 696 557 712
rect 573 696 591 712
rect 607 696 625 712
rect 641 696 659 712
rect 675 696 693 712
rect 709 696 727 712
rect 743 696 761 712
rect 777 696 795 712
rect 811 696 829 712
rect 845 696 863 712
rect 879 696 897 712
rect 913 696 931 712
rect 947 696 965 712
rect 981 696 999 712
rect 1015 696 1033 712
rect 1049 696 1067 712
rect 1083 696 1101 712
rect 1117 696 1135 712
rect 1151 696 1169 712
rect 1185 696 1203 712
rect 1219 696 1237 712
rect 1253 696 1271 712
rect 1287 696 1305 712
rect 1321 696 1339 712
rect 1355 696 1373 712
rect 1389 696 1407 712
rect 1423 696 1441 712
rect 1457 696 1475 712
rect 1491 696 1509 712
rect 1525 696 1543 712
rect 1559 696 1577 712
rect 1593 696 1611 712
rect 1627 696 1645 712
rect 1661 696 1679 712
rect 1695 696 1713 712
rect 1729 696 1747 712
rect 1763 696 1781 712
rect 1797 696 1815 712
rect 1831 696 1849 712
rect 1865 696 1883 712
rect 1899 696 1917 712
rect 1933 696 1951 712
rect 1967 696 1985 712
rect 2001 696 2019 712
rect 2035 696 2053 712
rect 2069 696 2087 712
rect 2103 696 2121 712
rect 2137 696 2155 712
rect 2171 696 2189 712
rect 2205 696 2223 712
rect 2239 696 2257 712
rect 2273 696 2291 712
rect 2307 696 2325 712
rect 2341 696 2359 712
rect 2375 696 2393 712
rect 2409 696 2427 712
rect 2443 696 2461 712
rect 2477 696 2495 712
rect 2511 696 2529 712
rect 2545 696 2563 712
rect 2579 696 2597 712
rect 2613 696 2631 712
rect 2647 696 2665 712
rect 2681 696 2699 712
rect 2715 696 2733 712
rect 2749 696 2767 712
rect 2783 696 2801 712
rect 2817 696 2835 712
rect 2851 696 2869 712
rect 2885 696 2903 712
rect 2919 696 2937 712
rect 2953 696 2971 712
rect 2987 696 3005 712
rect 3021 696 3042 712
rect 264 675 3042 696
rect 3180 794 3201 810
rect 3217 794 3235 810
rect 3251 794 3269 810
rect 3285 794 3306 810
rect 3180 776 3306 794
rect 3180 760 3201 776
rect 3217 760 3235 776
rect 3251 760 3269 776
rect 3285 760 3306 776
rect 3180 742 3306 760
rect 3180 726 3201 742
rect 3217 726 3235 742
rect 3251 726 3269 742
rect 3285 726 3306 742
rect 3180 708 3306 726
rect 3180 692 3201 708
rect 3217 692 3235 708
rect 3251 692 3269 708
rect 3285 692 3306 708
rect 0 658 21 674
rect 37 658 55 674
rect 71 658 89 674
rect 105 658 126 674
rect 0 640 126 658
rect 0 624 21 640
rect 37 624 55 640
rect 71 624 89 640
rect 105 624 126 640
rect 0 606 126 624
rect 0 590 21 606
rect 37 590 55 606
rect 71 590 89 606
rect 105 590 126 606
rect 0 576 126 590
rect 3180 674 3306 692
rect 3180 658 3201 674
rect 3217 658 3235 674
rect 3251 658 3269 674
rect 3285 658 3306 674
rect 3180 640 3306 658
rect 3180 624 3201 640
rect 3217 624 3235 640
rect 3251 624 3269 640
rect 3285 624 3306 640
rect 3180 606 3306 624
rect 3180 590 3201 606
rect 3217 590 3235 606
rect 3251 590 3269 606
rect 3285 590 3306 606
rect 3180 576 3306 590
rect 0 572 3306 576
rect 0 556 21 572
rect 37 556 55 572
rect 71 556 89 572
rect 105 556 3201 572
rect 3217 556 3235 572
rect 3251 556 3269 572
rect 3285 556 3306 572
rect 0 555 3306 556
rect 0 539 149 555
rect 165 539 183 555
rect 199 539 217 555
rect 233 539 251 555
rect 267 539 285 555
rect 301 539 319 555
rect 335 539 353 555
rect 369 539 387 555
rect 403 539 421 555
rect 437 539 455 555
rect 471 539 489 555
rect 505 539 523 555
rect 539 539 557 555
rect 573 539 591 555
rect 607 539 625 555
rect 641 539 659 555
rect 675 539 693 555
rect 709 539 727 555
rect 743 539 761 555
rect 777 539 795 555
rect 811 539 829 555
rect 845 539 863 555
rect 879 539 897 555
rect 913 539 931 555
rect 947 539 965 555
rect 981 539 999 555
rect 1015 539 1033 555
rect 1049 539 1067 555
rect 1083 539 1101 555
rect 1117 539 1135 555
rect 1151 539 1169 555
rect 1185 539 1203 555
rect 1219 539 1237 555
rect 1253 539 1271 555
rect 1287 539 1305 555
rect 1321 539 1339 555
rect 1355 539 1373 555
rect 1389 539 1407 555
rect 1423 539 1441 555
rect 1457 539 1475 555
rect 1491 539 1509 555
rect 1525 539 1543 555
rect 1559 539 1577 555
rect 1593 539 1611 555
rect 1627 539 1645 555
rect 1661 539 1679 555
rect 1695 539 1713 555
rect 1729 539 1747 555
rect 1763 539 1781 555
rect 1797 539 1815 555
rect 1831 539 1849 555
rect 1865 539 1883 555
rect 1899 539 1917 555
rect 1933 539 1951 555
rect 1967 539 1985 555
rect 2001 539 2019 555
rect 2035 539 2053 555
rect 2069 539 2087 555
rect 2103 539 2121 555
rect 2137 539 2155 555
rect 2171 539 2189 555
rect 2205 539 2223 555
rect 2239 539 2257 555
rect 2273 539 2291 555
rect 2307 539 2325 555
rect 2341 539 2359 555
rect 2375 539 2393 555
rect 2409 539 2427 555
rect 2443 539 2461 555
rect 2477 539 2495 555
rect 2511 539 2529 555
rect 2545 539 2563 555
rect 2579 539 2597 555
rect 2613 539 2631 555
rect 2647 539 2665 555
rect 2681 539 2699 555
rect 2715 539 2733 555
rect 2749 539 2767 555
rect 2783 539 2801 555
rect 2817 539 2835 555
rect 2851 539 2869 555
rect 2885 539 2903 555
rect 2919 539 2937 555
rect 2953 539 2971 555
rect 2987 539 3005 555
rect 3021 539 3039 555
rect 3055 539 3073 555
rect 3089 539 3107 555
rect 3123 539 3141 555
rect 3157 539 3306 555
rect 0 538 3306 539
rect 0 522 21 538
rect 37 522 55 538
rect 71 522 89 538
rect 105 522 3201 538
rect 3217 522 3235 538
rect 3251 522 3269 538
rect 3285 522 3306 538
rect 0 521 3306 522
rect 0 505 149 521
rect 165 505 183 521
rect 199 505 217 521
rect 233 505 251 521
rect 267 505 285 521
rect 301 505 319 521
rect 335 505 353 521
rect 369 505 387 521
rect 403 505 421 521
rect 437 505 455 521
rect 471 505 489 521
rect 505 505 523 521
rect 539 505 557 521
rect 573 505 591 521
rect 607 505 625 521
rect 641 505 659 521
rect 675 505 693 521
rect 709 505 727 521
rect 743 505 761 521
rect 777 505 795 521
rect 811 505 829 521
rect 845 505 863 521
rect 879 505 897 521
rect 913 505 931 521
rect 947 505 965 521
rect 981 505 999 521
rect 1015 505 1033 521
rect 1049 505 1067 521
rect 1083 505 1101 521
rect 1117 505 1135 521
rect 1151 505 1169 521
rect 1185 505 1203 521
rect 1219 505 1237 521
rect 1253 505 1271 521
rect 1287 505 1305 521
rect 1321 505 1339 521
rect 1355 505 1373 521
rect 1389 505 1407 521
rect 1423 505 1441 521
rect 1457 505 1475 521
rect 1491 505 1509 521
rect 1525 505 1543 521
rect 1559 505 1577 521
rect 1593 505 1611 521
rect 1627 505 1645 521
rect 1661 505 1679 521
rect 1695 505 1713 521
rect 1729 505 1747 521
rect 1763 505 1781 521
rect 1797 505 1815 521
rect 1831 505 1849 521
rect 1865 505 1883 521
rect 1899 505 1917 521
rect 1933 505 1951 521
rect 1967 505 1985 521
rect 2001 505 2019 521
rect 2035 505 2053 521
rect 2069 505 2087 521
rect 2103 505 2121 521
rect 2137 505 2155 521
rect 2171 505 2189 521
rect 2205 505 2223 521
rect 2239 505 2257 521
rect 2273 505 2291 521
rect 2307 505 2325 521
rect 2341 505 2359 521
rect 2375 505 2393 521
rect 2409 505 2427 521
rect 2443 505 2461 521
rect 2477 505 2495 521
rect 2511 505 2529 521
rect 2545 505 2563 521
rect 2579 505 2597 521
rect 2613 505 2631 521
rect 2647 505 2665 521
rect 2681 505 2699 521
rect 2715 505 2733 521
rect 2749 505 2767 521
rect 2783 505 2801 521
rect 2817 505 2835 521
rect 2851 505 2869 521
rect 2885 505 2903 521
rect 2919 505 2937 521
rect 2953 505 2971 521
rect 2987 505 3005 521
rect 3021 505 3039 521
rect 3055 505 3073 521
rect 3089 505 3107 521
rect 3123 505 3141 521
rect 3157 505 3306 521
rect 0 504 3306 505
rect 0 488 21 504
rect 37 488 55 504
rect 71 488 89 504
rect 105 488 3201 504
rect 3217 488 3235 504
rect 3251 488 3269 504
rect 3285 488 3306 504
rect 0 487 3306 488
rect 0 471 149 487
rect 165 471 183 487
rect 199 471 217 487
rect 233 471 251 487
rect 267 471 285 487
rect 301 471 319 487
rect 335 471 353 487
rect 369 471 387 487
rect 403 471 421 487
rect 437 471 455 487
rect 471 471 489 487
rect 505 471 523 487
rect 539 471 557 487
rect 573 471 591 487
rect 607 471 625 487
rect 641 471 659 487
rect 675 471 693 487
rect 709 471 727 487
rect 743 471 761 487
rect 777 471 795 487
rect 811 471 829 487
rect 845 471 863 487
rect 879 471 897 487
rect 913 471 931 487
rect 947 471 965 487
rect 981 471 999 487
rect 1015 471 1033 487
rect 1049 471 1067 487
rect 1083 471 1101 487
rect 1117 471 1135 487
rect 1151 471 1169 487
rect 1185 471 1203 487
rect 1219 471 1237 487
rect 1253 471 1271 487
rect 1287 471 1305 487
rect 1321 471 1339 487
rect 1355 471 1373 487
rect 1389 471 1407 487
rect 1423 471 1441 487
rect 1457 471 1475 487
rect 1491 471 1509 487
rect 1525 471 1543 487
rect 1559 471 1577 487
rect 1593 471 1611 487
rect 1627 471 1645 487
rect 1661 471 1679 487
rect 1695 471 1713 487
rect 1729 471 1747 487
rect 1763 471 1781 487
rect 1797 471 1815 487
rect 1831 471 1849 487
rect 1865 471 1883 487
rect 1899 471 1917 487
rect 1933 471 1951 487
rect 1967 471 1985 487
rect 2001 471 2019 487
rect 2035 471 2053 487
rect 2069 471 2087 487
rect 2103 471 2121 487
rect 2137 471 2155 487
rect 2171 471 2189 487
rect 2205 471 2223 487
rect 2239 471 2257 487
rect 2273 471 2291 487
rect 2307 471 2325 487
rect 2341 471 2359 487
rect 2375 471 2393 487
rect 2409 471 2427 487
rect 2443 471 2461 487
rect 2477 471 2495 487
rect 2511 471 2529 487
rect 2545 471 2563 487
rect 2579 471 2597 487
rect 2613 471 2631 487
rect 2647 471 2665 487
rect 2681 471 2699 487
rect 2715 471 2733 487
rect 2749 471 2767 487
rect 2783 471 2801 487
rect 2817 471 2835 487
rect 2851 471 2869 487
rect 2885 471 2903 487
rect 2919 471 2937 487
rect 2953 471 2971 487
rect 2987 471 3005 487
rect 3021 471 3039 487
rect 3055 471 3073 487
rect 3089 471 3107 487
rect 3123 471 3141 487
rect 3157 471 3306 487
rect 0 470 3306 471
rect 0 454 21 470
rect 37 454 55 470
rect 71 454 89 470
rect 105 454 3201 470
rect 3217 454 3235 470
rect 3251 454 3269 470
rect 3285 454 3306 470
rect 0 450 3306 454
rect 0 436 126 450
rect 0 420 21 436
rect 37 420 55 436
rect 71 420 89 436
rect 105 420 126 436
rect 0 402 126 420
rect 0 386 21 402
rect 37 386 55 402
rect 71 386 89 402
rect 105 386 126 402
rect 0 368 126 386
rect 0 352 21 368
rect 37 352 55 368
rect 71 352 89 368
rect 105 352 126 368
rect 0 334 126 352
rect 3180 436 3306 450
rect 3180 420 3201 436
rect 3217 420 3235 436
rect 3251 420 3269 436
rect 3285 420 3306 436
rect 3180 402 3306 420
rect 3180 386 3201 402
rect 3217 386 3235 402
rect 3251 386 3269 402
rect 3285 386 3306 402
rect 3180 368 3306 386
rect 3180 352 3201 368
rect 3217 352 3235 368
rect 3251 352 3269 368
rect 3285 352 3306 368
rect 0 318 21 334
rect 37 318 55 334
rect 71 318 89 334
rect 105 318 126 334
rect 0 300 126 318
rect 0 284 21 300
rect 37 284 55 300
rect 71 284 89 300
rect 105 284 126 300
rect 0 266 126 284
rect 0 250 21 266
rect 37 250 55 266
rect 71 250 89 266
rect 105 250 126 266
rect 0 232 126 250
rect 0 216 21 232
rect 37 216 55 232
rect 71 216 89 232
rect 105 216 126 232
rect 264 330 3042 351
rect 264 314 285 330
rect 301 314 319 330
rect 335 314 353 330
rect 369 314 387 330
rect 403 314 421 330
rect 437 314 455 330
rect 471 314 489 330
rect 505 314 523 330
rect 539 314 557 330
rect 573 314 591 330
rect 607 314 625 330
rect 641 314 659 330
rect 675 314 693 330
rect 709 314 727 330
rect 743 314 761 330
rect 777 314 795 330
rect 811 314 829 330
rect 845 314 863 330
rect 879 314 897 330
rect 913 314 931 330
rect 947 314 965 330
rect 981 314 999 330
rect 1015 314 1033 330
rect 1049 314 1067 330
rect 1083 314 1101 330
rect 1117 314 1135 330
rect 1151 314 1169 330
rect 1185 314 1203 330
rect 1219 314 1237 330
rect 1253 314 1271 330
rect 1287 314 1305 330
rect 1321 314 1339 330
rect 1355 314 1373 330
rect 1389 314 1407 330
rect 1423 314 1441 330
rect 1457 314 1475 330
rect 1491 314 1509 330
rect 1525 314 1543 330
rect 1559 314 1577 330
rect 1593 314 1611 330
rect 1627 314 1645 330
rect 1661 314 1679 330
rect 1695 314 1713 330
rect 1729 314 1747 330
rect 1763 314 1781 330
rect 1797 314 1815 330
rect 1831 314 1849 330
rect 1865 314 1883 330
rect 1899 314 1917 330
rect 1933 314 1951 330
rect 1967 314 1985 330
rect 2001 314 2019 330
rect 2035 314 2053 330
rect 2069 314 2087 330
rect 2103 314 2121 330
rect 2137 314 2155 330
rect 2171 314 2189 330
rect 2205 314 2223 330
rect 2239 314 2257 330
rect 2273 314 2291 330
rect 2307 314 2325 330
rect 2341 314 2359 330
rect 2375 314 2393 330
rect 2409 314 2427 330
rect 2443 314 2461 330
rect 2477 314 2495 330
rect 2511 314 2529 330
rect 2545 314 2563 330
rect 2579 314 2597 330
rect 2613 314 2631 330
rect 2647 314 2665 330
rect 2681 314 2699 330
rect 2715 314 2733 330
rect 2749 314 2767 330
rect 2783 314 2801 330
rect 2817 314 2835 330
rect 2851 314 2869 330
rect 2885 314 2903 330
rect 2919 314 2937 330
rect 2953 314 2971 330
rect 2987 314 3005 330
rect 3021 314 3042 330
rect 264 296 3042 314
rect 264 280 285 296
rect 301 280 319 296
rect 335 280 353 296
rect 369 280 387 296
rect 403 280 421 296
rect 437 280 455 296
rect 471 280 489 296
rect 505 280 523 296
rect 539 280 557 296
rect 573 280 591 296
rect 607 280 625 296
rect 641 280 659 296
rect 675 280 693 296
rect 709 280 727 296
rect 743 280 761 296
rect 777 280 795 296
rect 811 280 829 296
rect 845 280 863 296
rect 879 280 897 296
rect 913 280 931 296
rect 947 280 965 296
rect 981 280 999 296
rect 1015 280 1033 296
rect 1049 280 1067 296
rect 1083 280 1101 296
rect 1117 280 1135 296
rect 1151 280 1169 296
rect 1185 280 1203 296
rect 1219 280 1237 296
rect 1253 280 1271 296
rect 1287 280 1305 296
rect 1321 280 1339 296
rect 1355 280 1373 296
rect 1389 280 1407 296
rect 1423 280 1441 296
rect 1457 280 1475 296
rect 1491 280 1509 296
rect 1525 280 1543 296
rect 1559 280 1577 296
rect 1593 280 1611 296
rect 1627 280 1645 296
rect 1661 280 1679 296
rect 1695 280 1713 296
rect 1729 280 1747 296
rect 1763 280 1781 296
rect 1797 280 1815 296
rect 1831 280 1849 296
rect 1865 280 1883 296
rect 1899 280 1917 296
rect 1933 280 1951 296
rect 1967 280 1985 296
rect 2001 280 2019 296
rect 2035 280 2053 296
rect 2069 280 2087 296
rect 2103 280 2121 296
rect 2137 280 2155 296
rect 2171 280 2189 296
rect 2205 280 2223 296
rect 2239 280 2257 296
rect 2273 280 2291 296
rect 2307 280 2325 296
rect 2341 280 2359 296
rect 2375 280 2393 296
rect 2409 280 2427 296
rect 2443 280 2461 296
rect 2477 280 2495 296
rect 2511 280 2529 296
rect 2545 280 2563 296
rect 2579 280 2597 296
rect 2613 280 2631 296
rect 2647 280 2665 296
rect 2681 280 2699 296
rect 2715 280 2733 296
rect 2749 280 2767 296
rect 2783 280 2801 296
rect 2817 280 2835 296
rect 2851 280 2869 296
rect 2885 280 2903 296
rect 2919 280 2937 296
rect 2953 280 2971 296
rect 2987 280 3005 296
rect 3021 280 3042 296
rect 264 262 3042 280
rect 264 246 285 262
rect 301 246 319 262
rect 335 246 353 262
rect 369 246 387 262
rect 403 246 421 262
rect 437 246 455 262
rect 471 246 489 262
rect 505 246 523 262
rect 539 246 557 262
rect 573 246 591 262
rect 607 246 625 262
rect 641 246 659 262
rect 675 246 693 262
rect 709 246 727 262
rect 743 246 761 262
rect 777 246 795 262
rect 811 246 829 262
rect 845 246 863 262
rect 879 246 897 262
rect 913 246 931 262
rect 947 246 965 262
rect 981 246 999 262
rect 1015 246 1033 262
rect 1049 246 1067 262
rect 1083 246 1101 262
rect 1117 246 1135 262
rect 1151 246 1169 262
rect 1185 246 1203 262
rect 1219 246 1237 262
rect 1253 246 1271 262
rect 1287 246 1305 262
rect 1321 246 1339 262
rect 1355 246 1373 262
rect 1389 246 1407 262
rect 1423 246 1441 262
rect 1457 246 1475 262
rect 1491 246 1509 262
rect 1525 246 1543 262
rect 1559 246 1577 262
rect 1593 246 1611 262
rect 1627 246 1645 262
rect 1661 246 1679 262
rect 1695 246 1713 262
rect 1729 246 1747 262
rect 1763 246 1781 262
rect 1797 246 1815 262
rect 1831 246 1849 262
rect 1865 246 1883 262
rect 1899 246 1917 262
rect 1933 246 1951 262
rect 1967 246 1985 262
rect 2001 246 2019 262
rect 2035 246 2053 262
rect 2069 246 2087 262
rect 2103 246 2121 262
rect 2137 246 2155 262
rect 2171 246 2189 262
rect 2205 246 2223 262
rect 2239 246 2257 262
rect 2273 246 2291 262
rect 2307 246 2325 262
rect 2341 246 2359 262
rect 2375 246 2393 262
rect 2409 246 2427 262
rect 2443 246 2461 262
rect 2477 246 2495 262
rect 2511 246 2529 262
rect 2545 246 2563 262
rect 2579 246 2597 262
rect 2613 246 2631 262
rect 2647 246 2665 262
rect 2681 246 2699 262
rect 2715 246 2733 262
rect 2749 246 2767 262
rect 2783 246 2801 262
rect 2817 246 2835 262
rect 2851 246 2869 262
rect 2885 246 2903 262
rect 2919 246 2937 262
rect 2953 246 2971 262
rect 2987 246 3005 262
rect 3021 246 3042 262
rect 264 225 3042 246
rect 3180 334 3306 352
rect 3180 318 3201 334
rect 3217 318 3235 334
rect 3251 318 3269 334
rect 3285 318 3306 334
rect 3180 300 3306 318
rect 3180 284 3201 300
rect 3217 284 3235 300
rect 3251 284 3269 300
rect 3285 284 3306 300
rect 3180 266 3306 284
rect 3180 250 3201 266
rect 3217 250 3235 266
rect 3251 250 3269 266
rect 3285 250 3306 266
rect 3180 232 3306 250
rect 0 198 126 216
rect 0 182 21 198
rect 37 182 55 198
rect 71 182 89 198
rect 105 182 126 198
rect 0 164 126 182
rect 0 148 21 164
rect 37 148 55 164
rect 71 148 89 164
rect 105 148 126 164
rect 0 130 126 148
rect 0 114 21 130
rect 37 114 55 130
rect 71 114 89 130
rect 105 126 126 130
rect 3180 216 3201 232
rect 3217 216 3235 232
rect 3251 216 3269 232
rect 3285 216 3306 232
rect 3180 198 3306 216
rect 3180 182 3201 198
rect 3217 182 3235 198
rect 3251 182 3269 198
rect 3285 182 3306 198
rect 3180 164 3306 182
rect 3180 148 3201 164
rect 3217 148 3235 164
rect 3251 148 3269 164
rect 3285 148 3306 164
rect 3180 130 3306 148
rect 3180 126 3201 130
rect 105 114 3201 126
rect 3217 114 3235 130
rect 3251 114 3269 130
rect 3285 114 3306 130
rect 0 105 3306 114
rect 0 96 149 105
rect 0 80 21 96
rect 37 80 55 96
rect 71 80 89 96
rect 105 89 149 96
rect 165 89 183 105
rect 199 89 217 105
rect 233 89 251 105
rect 267 89 285 105
rect 301 89 319 105
rect 335 89 353 105
rect 369 89 387 105
rect 403 89 421 105
rect 437 89 455 105
rect 471 89 489 105
rect 505 89 523 105
rect 539 89 557 105
rect 573 89 591 105
rect 607 89 625 105
rect 641 89 659 105
rect 675 89 693 105
rect 709 89 727 105
rect 743 89 761 105
rect 777 89 795 105
rect 811 89 829 105
rect 845 89 863 105
rect 879 89 897 105
rect 913 89 931 105
rect 947 89 965 105
rect 981 89 999 105
rect 1015 89 1033 105
rect 1049 89 1067 105
rect 1083 89 1101 105
rect 1117 89 1135 105
rect 1151 89 1169 105
rect 1185 89 1203 105
rect 1219 89 1237 105
rect 1253 89 1271 105
rect 1287 89 1305 105
rect 1321 89 1339 105
rect 1355 89 1373 105
rect 1389 89 1407 105
rect 1423 89 1441 105
rect 1457 89 1475 105
rect 1491 89 1509 105
rect 1525 89 1543 105
rect 1559 89 1577 105
rect 1593 89 1611 105
rect 1627 89 1645 105
rect 1661 89 1679 105
rect 1695 89 1713 105
rect 1729 89 1747 105
rect 1763 89 1781 105
rect 1797 89 1815 105
rect 1831 89 1849 105
rect 1865 89 1883 105
rect 1899 89 1917 105
rect 1933 89 1951 105
rect 1967 89 1985 105
rect 2001 89 2019 105
rect 2035 89 2053 105
rect 2069 89 2087 105
rect 2103 89 2121 105
rect 2137 89 2155 105
rect 2171 89 2189 105
rect 2205 89 2223 105
rect 2239 89 2257 105
rect 2273 89 2291 105
rect 2307 89 2325 105
rect 2341 89 2359 105
rect 2375 89 2393 105
rect 2409 89 2427 105
rect 2443 89 2461 105
rect 2477 89 2495 105
rect 2511 89 2529 105
rect 2545 89 2563 105
rect 2579 89 2597 105
rect 2613 89 2631 105
rect 2647 89 2665 105
rect 2681 89 2699 105
rect 2715 89 2733 105
rect 2749 89 2767 105
rect 2783 89 2801 105
rect 2817 89 2835 105
rect 2851 89 2869 105
rect 2885 89 2903 105
rect 2919 89 2937 105
rect 2953 89 2971 105
rect 2987 89 3005 105
rect 3021 89 3039 105
rect 3055 89 3073 105
rect 3089 89 3107 105
rect 3123 89 3141 105
rect 3157 96 3306 105
rect 3157 89 3201 96
rect 105 80 3201 89
rect 3217 80 3235 96
rect 3251 80 3269 96
rect 3285 80 3306 96
rect 0 71 3306 80
rect 0 62 149 71
rect 0 46 21 62
rect 37 46 55 62
rect 71 46 89 62
rect 105 55 149 62
rect 165 55 183 71
rect 199 55 217 71
rect 233 55 251 71
rect 267 55 285 71
rect 301 55 319 71
rect 335 55 353 71
rect 369 55 387 71
rect 403 55 421 71
rect 437 55 455 71
rect 471 55 489 71
rect 505 55 523 71
rect 539 55 557 71
rect 573 55 591 71
rect 607 55 625 71
rect 641 55 659 71
rect 675 55 693 71
rect 709 55 727 71
rect 743 55 761 71
rect 777 55 795 71
rect 811 55 829 71
rect 845 55 863 71
rect 879 55 897 71
rect 913 55 931 71
rect 947 55 965 71
rect 981 55 999 71
rect 1015 55 1033 71
rect 1049 55 1067 71
rect 1083 55 1101 71
rect 1117 55 1135 71
rect 1151 55 1169 71
rect 1185 55 1203 71
rect 1219 55 1237 71
rect 1253 55 1271 71
rect 1287 55 1305 71
rect 1321 55 1339 71
rect 1355 55 1373 71
rect 1389 55 1407 71
rect 1423 55 1441 71
rect 1457 55 1475 71
rect 1491 55 1509 71
rect 1525 55 1543 71
rect 1559 55 1577 71
rect 1593 55 1611 71
rect 1627 55 1645 71
rect 1661 55 1679 71
rect 1695 55 1713 71
rect 1729 55 1747 71
rect 1763 55 1781 71
rect 1797 55 1815 71
rect 1831 55 1849 71
rect 1865 55 1883 71
rect 1899 55 1917 71
rect 1933 55 1951 71
rect 1967 55 1985 71
rect 2001 55 2019 71
rect 2035 55 2053 71
rect 2069 55 2087 71
rect 2103 55 2121 71
rect 2137 55 2155 71
rect 2171 55 2189 71
rect 2205 55 2223 71
rect 2239 55 2257 71
rect 2273 55 2291 71
rect 2307 55 2325 71
rect 2341 55 2359 71
rect 2375 55 2393 71
rect 2409 55 2427 71
rect 2443 55 2461 71
rect 2477 55 2495 71
rect 2511 55 2529 71
rect 2545 55 2563 71
rect 2579 55 2597 71
rect 2613 55 2631 71
rect 2647 55 2665 71
rect 2681 55 2699 71
rect 2715 55 2733 71
rect 2749 55 2767 71
rect 2783 55 2801 71
rect 2817 55 2835 71
rect 2851 55 2869 71
rect 2885 55 2903 71
rect 2919 55 2937 71
rect 2953 55 2971 71
rect 2987 55 3005 71
rect 3021 55 3039 71
rect 3055 55 3073 71
rect 3089 55 3107 71
rect 3123 55 3141 71
rect 3157 62 3306 71
rect 3157 55 3201 62
rect 105 46 3201 55
rect 3217 46 3235 62
rect 3251 46 3269 62
rect 3285 46 3306 62
rect 0 37 3306 46
rect 0 28 149 37
rect 0 12 21 28
rect 37 12 55 28
rect 71 12 89 28
rect 105 21 149 28
rect 165 21 183 37
rect 199 21 217 37
rect 233 21 251 37
rect 267 21 285 37
rect 301 21 319 37
rect 335 21 353 37
rect 369 21 387 37
rect 403 21 421 37
rect 437 21 455 37
rect 471 21 489 37
rect 505 21 523 37
rect 539 21 557 37
rect 573 21 591 37
rect 607 21 625 37
rect 641 21 659 37
rect 675 21 693 37
rect 709 21 727 37
rect 743 21 761 37
rect 777 21 795 37
rect 811 21 829 37
rect 845 21 863 37
rect 879 21 897 37
rect 913 21 931 37
rect 947 21 965 37
rect 981 21 999 37
rect 1015 21 1033 37
rect 1049 21 1067 37
rect 1083 21 1101 37
rect 1117 21 1135 37
rect 1151 21 1169 37
rect 1185 21 1203 37
rect 1219 21 1237 37
rect 1253 21 1271 37
rect 1287 21 1305 37
rect 1321 21 1339 37
rect 1355 21 1373 37
rect 1389 21 1407 37
rect 1423 21 1441 37
rect 1457 21 1475 37
rect 1491 21 1509 37
rect 1525 21 1543 37
rect 1559 21 1577 37
rect 1593 21 1611 37
rect 1627 21 1645 37
rect 1661 21 1679 37
rect 1695 21 1713 37
rect 1729 21 1747 37
rect 1763 21 1781 37
rect 1797 21 1815 37
rect 1831 21 1849 37
rect 1865 21 1883 37
rect 1899 21 1917 37
rect 1933 21 1951 37
rect 1967 21 1985 37
rect 2001 21 2019 37
rect 2035 21 2053 37
rect 2069 21 2087 37
rect 2103 21 2121 37
rect 2137 21 2155 37
rect 2171 21 2189 37
rect 2205 21 2223 37
rect 2239 21 2257 37
rect 2273 21 2291 37
rect 2307 21 2325 37
rect 2341 21 2359 37
rect 2375 21 2393 37
rect 2409 21 2427 37
rect 2443 21 2461 37
rect 2477 21 2495 37
rect 2511 21 2529 37
rect 2545 21 2563 37
rect 2579 21 2597 37
rect 2613 21 2631 37
rect 2647 21 2665 37
rect 2681 21 2699 37
rect 2715 21 2733 37
rect 2749 21 2767 37
rect 2783 21 2801 37
rect 2817 21 2835 37
rect 2851 21 2869 37
rect 2885 21 2903 37
rect 2919 21 2937 37
rect 2953 21 2971 37
rect 2987 21 3005 37
rect 3021 21 3039 37
rect 3055 21 3073 37
rect 3089 21 3107 37
rect 3123 21 3141 37
rect 3157 28 3306 37
rect 3157 21 3201 28
rect 105 12 3201 21
rect 3217 12 3235 28
rect 3251 12 3269 28
rect 3285 12 3306 28
rect 0 0 3306 12
rect 3438 1015 3447 1031
rect 3463 1015 3472 1031
rect 3438 997 3472 1015
rect 3438 981 3447 997
rect 3463 981 3472 997
rect 3438 963 3472 981
rect 3438 947 3447 963
rect 3463 947 3472 963
rect 3438 929 3472 947
rect 3438 913 3447 929
rect 3463 913 3472 929
rect 3438 895 3472 913
rect 3438 879 3447 895
rect 3463 879 3472 895
rect 3438 861 3472 879
rect 3438 845 3447 861
rect 3463 845 3472 861
rect 3438 827 3472 845
rect 3438 811 3447 827
rect 3463 811 3472 827
rect 3438 793 3472 811
rect 3438 777 3447 793
rect 3463 777 3472 793
rect 3438 759 3472 777
rect 3438 743 3447 759
rect 3463 743 3472 759
rect 3438 725 3472 743
rect 3438 709 3447 725
rect 3463 709 3472 725
rect 3438 691 3472 709
rect 3438 675 3447 691
rect 3463 675 3472 691
rect 3438 657 3472 675
rect 3438 641 3447 657
rect 3463 641 3472 657
rect 3438 623 3472 641
rect 3438 607 3447 623
rect 3463 607 3472 623
rect 3438 589 3472 607
rect 3438 573 3447 589
rect 3463 573 3472 589
rect 3438 555 3472 573
rect 3438 539 3447 555
rect 3463 539 3472 555
rect 3438 521 3472 539
rect 3438 505 3447 521
rect 3463 505 3472 521
rect 3438 487 3472 505
rect 3438 471 3447 487
rect 3463 471 3472 487
rect 3438 453 3472 471
rect 3438 437 3447 453
rect 3463 437 3472 453
rect 3438 419 3472 437
rect 3438 403 3447 419
rect 3463 403 3472 419
rect 3438 385 3472 403
rect 3438 369 3447 385
rect 3463 369 3472 385
rect 3438 351 3472 369
rect 3438 335 3447 351
rect 3463 335 3472 351
rect 3438 317 3472 335
rect 3438 301 3447 317
rect 3463 301 3472 317
rect 3438 283 3472 301
rect 3438 267 3447 283
rect 3463 267 3472 283
rect 3438 249 3472 267
rect 3438 233 3447 249
rect 3463 233 3472 249
rect 3438 215 3472 233
rect 3438 199 3447 215
rect 3463 199 3472 215
rect 3438 181 3472 199
rect 3438 165 3447 181
rect 3463 165 3472 181
rect 3438 147 3472 165
rect 3438 131 3447 147
rect 3463 131 3472 147
rect 3438 113 3472 131
rect 3438 97 3447 113
rect 3463 97 3472 113
rect 3438 79 3472 97
rect 3438 63 3447 79
rect 3463 63 3472 79
rect 3438 45 3472 63
rect 3438 29 3447 45
rect 3463 29 3472 45
rect 3438 11 3472 29
rect -166 -23 -132 -5
rect -166 -39 -157 -23
rect -141 -39 -132 -23
rect -166 -57 -132 -39
rect -166 -73 -157 -57
rect -141 -73 -132 -57
rect -166 -91 -132 -73
rect -166 -107 -157 -91
rect -141 -107 -132 -91
rect -166 -132 -132 -107
rect 3438 -5 3447 11
rect 3463 -5 3472 11
rect 3438 -23 3472 -5
rect 3438 -39 3447 -23
rect 3463 -39 3472 -23
rect 3438 -57 3472 -39
rect 3438 -73 3447 -57
rect 3463 -73 3472 -57
rect 3438 -91 3472 -73
rect 3438 -107 3447 -91
rect 3463 -107 3472 -91
rect 3438 -132 3472 -107
rect -166 -141 3472 -132
rect -166 -157 -157 -141
rect -141 -157 -123 -141
rect -107 -157 -89 -141
rect -73 -157 -55 -141
rect -39 -157 -21 -141
rect -5 -157 13 -141
rect 29 -157 47 -141
rect 63 -157 81 -141
rect 97 -157 115 -141
rect 131 -157 149 -141
rect 165 -157 183 -141
rect 199 -157 217 -141
rect 233 -157 251 -141
rect 267 -157 285 -141
rect 301 -157 319 -141
rect 335 -157 353 -141
rect 369 -157 387 -141
rect 403 -157 421 -141
rect 437 -157 455 -141
rect 471 -157 489 -141
rect 505 -157 523 -141
rect 539 -157 557 -141
rect 573 -157 591 -141
rect 607 -157 625 -141
rect 641 -157 659 -141
rect 675 -157 693 -141
rect 709 -157 727 -141
rect 743 -157 761 -141
rect 777 -157 795 -141
rect 811 -157 829 -141
rect 845 -157 863 -141
rect 879 -157 897 -141
rect 913 -157 931 -141
rect 947 -157 965 -141
rect 981 -157 999 -141
rect 1015 -157 1033 -141
rect 1049 -157 1067 -141
rect 1083 -157 1101 -141
rect 1117 -157 1135 -141
rect 1151 -157 1169 -141
rect 1185 -157 1203 -141
rect 1219 -157 1237 -141
rect 1253 -157 1271 -141
rect 1287 -157 1305 -141
rect 1321 -157 1339 -141
rect 1355 -157 1373 -141
rect 1389 -157 1407 -141
rect 1423 -157 1441 -141
rect 1457 -157 1475 -141
rect 1491 -157 1509 -141
rect 1525 -157 1543 -141
rect 1559 -157 1577 -141
rect 1593 -157 1611 -141
rect 1627 -157 1645 -141
rect 1661 -157 1679 -141
rect 1695 -157 1713 -141
rect 1729 -157 1747 -141
rect 1763 -157 1781 -141
rect 1797 -157 1815 -141
rect 1831 -157 1849 -141
rect 1865 -157 1883 -141
rect 1899 -157 1917 -141
rect 1933 -157 1951 -141
rect 1967 -157 1985 -141
rect 2001 -157 2019 -141
rect 2035 -157 2053 -141
rect 2069 -157 2087 -141
rect 2103 -157 2121 -141
rect 2137 -157 2155 -141
rect 2171 -157 2189 -141
rect 2205 -157 2223 -141
rect 2239 -157 2257 -141
rect 2273 -157 2291 -141
rect 2307 -157 2325 -141
rect 2341 -157 2359 -141
rect 2375 -157 2393 -141
rect 2409 -157 2427 -141
rect 2443 -157 2461 -141
rect 2477 -157 2495 -141
rect 2511 -157 2529 -141
rect 2545 -157 2563 -141
rect 2579 -157 2597 -141
rect 2613 -157 2631 -141
rect 2647 -157 2665 -141
rect 2681 -157 2699 -141
rect 2715 -157 2733 -141
rect 2749 -157 2767 -141
rect 2783 -157 2801 -141
rect 2817 -157 2835 -141
rect 2851 -157 2869 -141
rect 2885 -157 2903 -141
rect 2919 -157 2937 -141
rect 2953 -157 2971 -141
rect 2987 -157 3005 -141
rect 3021 -157 3039 -141
rect 3055 -157 3073 -141
rect 3089 -157 3107 -141
rect 3123 -157 3141 -141
rect 3157 -157 3175 -141
rect 3191 -157 3209 -141
rect 3225 -157 3243 -141
rect 3259 -157 3277 -141
rect 3293 -157 3311 -141
rect 3327 -157 3345 -141
rect 3361 -157 3379 -141
rect 3395 -157 3413 -141
rect 3429 -157 3447 -141
rect 3463 -157 3472 -141
rect -166 -166 3472 -157
<< labels >>
flabel comment s 716 732 716 732 0 FreeSans 200 0 0 0 dpant
flabel comment s 704 284 704 284 0 FreeSans 200 0 0 0 dpant
rlabel comment s -149 -30 -149 -30 4 sub!
rlabel metal1 s -166 1158 3472 1192 4 guard
port 2 nsew
rlabel metal1 s -166 -166 3472 -132 4 guard
port 2 nsew
rlabel metal1 s 0 450 3306 576 4 cathode
port 3 nsew
rlabel metal1 s 0 0 3306 126 4 cathode
port 3 nsew
rlabel metal1 s 0 900 3306 1026 4 cathode
port 3 nsew
rlabel metal1 s 264 675 3042 801 4 anode
port 4 nsew
rlabel metal1 s 264 225 3042 351 4 anode
port 4 nsew
<< end >>
