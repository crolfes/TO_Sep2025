** Created by: circuit_gen.AN2D1_1
** Cell name: AN2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_AN2D1_1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AN2D1_2
** Cell name: AN2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_AN2D1_2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AN2D1_3
** Cell name: AN2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_AN2D1_3 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AN2D1
** Cell name: AN2D1
** Lib name: sg13g2
.SUBCKT sg13g2_AN2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AO21D1_1
** Cell name: AO21D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_AO21D1_1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AO21D1_2
** Cell name: AO21D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_AO21D1_2 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AO21D1_3
** Cell name: AO21D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_AO21D1_3 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AO21D1
** Cell name: AO21D1
** Lib name: sg13g2
.SUBCKT sg13g2_AO21D1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AOI21D1_1
** Cell name: AOI21D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_AOI21D1_1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 zn b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net13 a2 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u3 net13 a1 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AOI21D1_2
** Cell name: AOI21D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_AOI21D1_2 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 zn b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net13 a2 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u3 net13 a1 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AOI21D1_3
** Cell name: AOI21D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_AOI21D1_3 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 zn b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net13 a2 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u3 net13 a1 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AOI21D1
** Cell name: AOI21D1
** Lib name: sg13g2
.SUBCKT sg13g2_AOI21D1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 zn b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net13 a2 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u3 net13 a1 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ANTENNA
** Cell name: ANTENNA
** Lib name: sg13g2f
.SUBCKT sg13g2_ANTENNA i vdd vss
*.PININFO i:I vdd:B vss:B
Ddn_1 vss i dantenna m=1 w=1.485u l=970n a=1440.45f
DD0 i vdd dpantenna m=1 w=1.485u l=970n a=1440.45f
.ENDS


******* EOF

** Created by: circuit_gen.BUFFD1_1
** Cell name: BUFFD1_1
** Lib name: sg13g2
.SUBCKT sg13g2_BUFFD1_1 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.BUFFD1_2
** Cell name: BUFFD1_2
** Lib name: sg13g2
.SUBCKT sg13g2_BUFFD1_2 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.BUFFD1_3
** Cell name: BUFFD1_3
** Lib name: sg13g2
.SUBCKT sg13g2_BUFFD1_3 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.BUFFD1
** Cell name: BUFFD1
** Lib name: sg13g2
.SUBCKT sg13g2_BUFFD1 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.DFCNQD1
** Cell name: DFCNQD1
** Lib name: sg13g2
.SUBCKT sg13g2_DFCNQD1 cdn cp d q vdd vss
*.PININFO cdn:I cp:I d:I q:O vdd:B vss:B 
Mcpbn incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=0 $flip=0
Mcpbp incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07 $pos=0 $flip=0
Mcpn incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=1 $flip=1
Mcpp incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07 $pos=1 $flip=1
MI4 net52 incpb vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=3 $flip=1
MI7 net85 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07 $pos=3 $flip=1
Mdd0n d0 d net52 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=4 $flip=1
Mdd0p d0 d net85 vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07 $pos=4 $flip=1
MI47 d0 incp net59 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=5 $flip=0
MI45 d0 incpb net98 vdd sg13_lv_pmos l=1.300e-07 w=3.300e-07 $pos=5 $flip=0
MI48 net59 d1 net62 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=6 $flip=0
MI43 net98 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=3.050e-07 $pos=6 $flip=0
Mcdn0n net62 cdn vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=7 $flip=0
Md0d1n d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=8 $flip=1
Mcdn0p net98 cdn vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=8 $flip=0
Mswd1d2n d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=4.900e-07 $pos=9 $flip=0
Mdod1p d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.150e-07 $pos=9 $flip=1
MI23 d2 incpb net57 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=10 $flip=0
Mswd1d2p d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=1.030e-06 $pos=10 $flip=0
MI26 d2 incp net88 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=11 $flip=0
MI24 net57 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=12 $flip=0
MI28 net88 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=12 $flip=0
Mcdn1n net37 cdn vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=13 $flip=1
Mcdn1p d3 cdn vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07 $pos=13 $flip=1
Md2d3n d3 d2 net37 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=14 $flip=1
Md2d3p d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07 $pos=14 $flip=0
Mobp q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06 $pos=15 $flip=1
Mobn q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=16 $flip=1
.ENDS


******* EOF

** Created by: circuit_gen.DFQD1_1
** Cell name: DFQD1_1
** Lib name: sg13g2
.SUBCKT sg13g2_DFQD1_1 cp d q vdd vss
*.PININFO cp:I d:I q:O vdd:B vss:B 
MI4 net43 incpb vss vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI23 d2 incpb net42 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI5 d0 d net43 vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI47 d0 incp net50 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI48 net50 d1 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI24 net42 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI50 d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=3.750e-07
MI32_M_u2 incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI31_M_u2 incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI27_M_u2 q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI53_M_u2 d3 d2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI13_M_u2 d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.550e-07
MI6 d0 d net66 vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI32_M_u3 incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI31_M_u3 incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI27_M_u3 q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI53_M_u3 d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI13_M_u3 d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI7 net66 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07
MI52 d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI28 net74 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI26 d2 incp net74 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI45 d0 incpb net84 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI43 net84 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
.ENDS


******* EOF

** Created by: circuit_gen.DFQD1_2
** Cell name: DFQD1_2
** Lib name: sg13g2
.SUBCKT sg13g2_DFQD1_2 cp d q vdd vss
*.PININFO cp:I d:I q:O vdd:B vss:B 
MI4 net43 incpb vss vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI23 d2 incpb net42 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI5 d0 d net43 vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI47 d0 incp net50 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI48 net50 d1 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI24 net42 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI50 d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=3.750e-07
MI32_M_u2 incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI31_M_u2 incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI27_M_u2 q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI53_M_u2 d3 d2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI13_M_u2 d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.550e-07
MI6 d0 d net66 vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI32_M_u3 incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI31_M_u3 incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI27_M_u3 q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI53_M_u3 d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI13_M_u3 d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI7 net66 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07
MI52 d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI28 net74 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI26 d2 incp net74 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI45 d0 incpb net84 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI43 net84 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
.ENDS


******* EOF

** Created by: circuit_gen.DFQD1_3
** Cell name: DFQD1_3
** Lib name: sg13g2
.SUBCKT sg13g2_DFQD1_3 cp d q vdd vss
*.PININFO cp:I d:I q:O vdd:B vss:B 
MI4 net43 incpb vss vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI23 d2 incpb net42 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI5 d0 d net43 vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI47 d0 incp net50 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI48 net50 d1 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI24 net42 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI50 d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=3.750e-07
MI32_M_u2 incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI31_M_u2 incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI27_M_u2 q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI53_M_u2 d3 d2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI13_M_u2 d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.550e-07
MI6 d0 d net66 vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI32_M_u3 incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI31_M_u3 incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI27_M_u3 q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI53_M_u3 d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI13_M_u3 d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI7 net66 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07
MI52 d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI28 net74 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI26 d2 incp net74 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI45 d0 incpb net84 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI43 net84 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
.ENDS


******* EOF

** Created by: circuit_gen.DFQD1
** Cell name: DFQD1
** Lib name: sg13g2
.SUBCKT sg13g2_DFQD1 cp d q vdd vss
*.PININFO cp:I d:I q:O vdd:B vss:B 
MI4 net43 incpb vss vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI23 d2 incpb net42 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI5 d0 d net43 vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI47 d0 incp net50 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI48 net50 d1 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI24 net42 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI50 d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=3.750e-07
MI32_M_u2 incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI31_M_u2 incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI27_M_u2 q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI53_M_u2 d3 d2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI13_M_u2 d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.550e-07
MI6 d0 d net66 vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI32_M_u3 incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI31_M_u3 incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI27_M_u3 q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI53_M_u3 d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI13_M_u3 d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI7 net66 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07
MI52 d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI28 net74 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI26 d2 incp net74 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI45 d0 incpb net84 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI43 net84 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
.ENDS


******* EOF

** Created by: circuit_gen.FILL1
** Cell name: FILL1
** Lib name: sg13g2
.SUBCKT sg13g2_FILL1 vdd vss
*.PININFO vdd:B vss:B 
.ENDS


******* EOF

** Created by: circuit_gen.FILL2
** Cell name: FILL2
** Lib name: sg13g2
.SUBCKT sg13g2_FILL2 vdd vss
*.PININFO vdd:B vss:B 
.ENDS


******* EOF

** Created by: circuit_gen.FILL4
** Cell name: FILL4
** Lib name: sg13g2
.SUBCKT sg13g2_FILL4 vdd vss
*.PININFO vdd:B vss:B 
.ENDS


******* EOF

** Created by: circuit_gen.FILL8
** Cell name: FILL8
** Lib name: sg13g2
.SUBCKT sg13g2_FILL8 vdd vss
*.PININFO vdd:B vss:B 
.ENDS


******* EOF

** Created by: circuit_gen.INVD1_1
** Cell name: INVD1_1
** Lib name: sg13g2
.SUBCKT sg13g2_INVD1_1 i z vss vdd
*.PININFO i:I z:O vss:B vdd:B
M0 z i vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M1 z i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.INVD1_2
** Cell name: INVD1_2
** Lib name: sg13g2
.SUBCKT sg13g2_INVD1_2 i z vss vdd
*.PININFO i:I z:O vss:B vdd:B
M0 z i vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M1 z i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.INVD1_3
** Cell name: INVD1_3
** Lib name: sg13g2
.SUBCKT sg13g2_INVD1_3 i z vss vdd
*.PININFO i:I z:O vss:B vdd:B
M0 z i vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M1 z i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.INVD1
** Cell name: INVD1
** Lib name: sg13g2
.SUBCKT sg13g2_INVD1 i z vss vdd
*.PININFO i:I z:O vss:B vdd:B
M0 z i vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M1 z i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.MUX2D1_1
** Cell name: MUX2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_MUX2D1_1 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.050e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.100e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.700e-07
.ENDS


******* EOF

** Created by: circuit_gen.MUX2D1_2
** Cell name: MUX2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_MUX2D1_2 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.050e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.100e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.700e-07
.ENDS


******* EOF

** Created by: circuit_gen.MUX2D1_3
** Cell name: MUX2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_MUX2D1_3 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.050e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.100e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.700e-07
.ENDS


******* EOF

** Created by: circuit_gen.MUX2D1
** Cell name: MUX2D1
** Lib name: sg13g2
.SUBCKT sg13g2_MUX2D1 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.050e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.100e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.700e-07
.ENDS


******* EOF

** Created by: circuit_gen.ND2D1_1
** Cell name: ND2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_ND2D1_1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u3 zn a1 xi1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u4 xi1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND2D1_2
** Cell name: ND2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_ND2D1_2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u3 zn a1 xi1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u4 xi1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND2D1_3
** Cell name: ND2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_ND2D1_3 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u3 zn a1 xi1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u4 xi1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND2D1
** Cell name: ND2D1
** Lib name: sg13g2
.SUBCKT sg13g2_ND2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u3 zn a1 xi1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u4 xi1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND3D1_1
** Cell name: ND3D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_ND3D1_1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 xi1_net10 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u5 xi1_net10 a2 xi1_net13 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u6 xi1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND3D1_2
** Cell name: ND3D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_ND3D1_2 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 xi1_net10 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u5 xi1_net10 a2 xi1_net13 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u6 xi1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND3D1_3
** Cell name: ND3D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_ND3D1_3 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 xi1_net10 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u5 xi1_net10 a2 xi1_net13 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u6 xi1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND3D1
** Cell name: ND3D1
** Lib name: sg13g2
.SUBCKT sg13g2_ND3D1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 xi1_net10 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u5 xi1_net10 a2 xi1_net13 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u6 xi1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND4D1_1
** Cell name: ND4D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_ND4D1_1 a1 a2 a3 a4 vdd vss zn
*.PININFO a1:I a2:I a3:I a4:I zn:O vdd:B vss:B 
MI3 p0 a2 p1 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5 p2 a4 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4 p1 a3 p2 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MU53 zn a1 p0 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI7 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI2 zn a4 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI0 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND4D1_2
** Cell name: ND4D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_ND4D1_2 a1 a2 a3 a4 vdd vss zn
*.PININFO a1:I a2:I a3:I a4:I zn:O vdd:B vss:B 
MI3 p0 a2 p1 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5 p2 a4 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4 p1 a3 p2 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MU53 zn a1 p0 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI7 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI2 zn a4 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI0 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND4D1_3
** Cell name: ND4D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_ND4D1_3 a1 a2 a3 a4 vdd vss zn
*.PININFO a1:I a2:I a3:I a4:I zn:O vdd:B vss:B 
MI3 p0 a2 p1 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5 p2 a4 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4 p1 a3 p2 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MU53 zn a1 p0 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI7 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI2 zn a4 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI0 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND4D1
** Cell name: ND4D1
** Lib name: sg13g2
.SUBCKT sg13g2_ND4D1 a1 a2 a3 a4 vdd vss zn
*.PININFO a1:I a2:I a3:I a4:I zn:O vdd:B vss:B 
MI3 p0 a2 p1 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5 p2 a4 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4 p1 a3 p2 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MU53 zn a1 p0 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI7 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI2 zn a4 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI0 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR2D1_1
** Cell name: NR2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_NR2D1_1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR2D1_2
** Cell name: NR2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_NR2D1_2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR2D1_3
** Cell name: NR2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_NR2D1_3 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR2D1
** Cell name: NR2D1
** Lib name: sg13g2
.SUBCKT sg13g2_NR2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR3D1_1
** Cell name: NR3D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_NR3D1_1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_0 net37_0_ a2 net34_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_0 net34_0_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_1 net34_1_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_1 net37_1_ a2 net34_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_0 zn a1 net37_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_1 zn a1 net37_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR3D1_2
** Cell name: NR3D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_NR3D1_2 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_0 net37_0_ a2 net34_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_0 net34_0_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_1 net34_1_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_1 net37_1_ a2 net34_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_0 zn a1 net37_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_1 zn a1 net37_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR3D1_3
** Cell name: NR3D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_NR3D1_3 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_0 net37_0_ a2 net34_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_0 net34_0_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_1 net34_1_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_1 net37_1_ a2 net34_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_0 zn a1 net37_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_1 zn a1 net37_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR3D1
** Cell name: NR3D1
** Lib name: sg13g2
.SUBCKT sg13g2_NR3D1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_0 net37_0_ a2 net34_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_0 net34_0_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_1 net34_1_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_1 net37_1_ a2 net34_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_0 zn a1 net37_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_1 zn a1 net37_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OA21D1_1
** Cell name: OA21D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_OA21D1_1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OA21D1_2
** Cell name: OA21D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_OA21D1_2 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OA21D1_3
** Cell name: OA21D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_OA21D1_3 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OA21D1
** Cell name: OA21D1
** Lib name: sg13g2
.SUBCKT sg13g2_OA21D1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OAI21D1_1
** Cell name: OAI21D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_OAI21D1_1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OAI21D1_2
** Cell name: OAI21D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_OAI21D1_2 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OAI21D1_3
** Cell name: OAI21D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_OAI21D1_3 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OAI21D1
** Cell name: OAI21D1
** Lib name: sg13g2
.SUBCKT sg13g2_OAI21D1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OR2D1_1
** Cell name: OR2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_OR2D1_1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OR2D1_2
** Cell name: OR2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_OR2D1_2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OR2D1_3
** Cell name: OR2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_OR2D1_3 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OR2D1
** Cell name: OR2D1
** Lib name: sg13g2
.SUBCKT sg13g2_OR2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TAPCELL
** Cell name: TAPCELL
** Lib name: sg13g2
.SUBCKT sg13g2_TAPCELL vdd vss
*.PININFO vdd:B vss:B 
.ENDS


******* EOF

** Created by: circuit_gen.TIEH_1
** Cell name: TIEH_1
** Lib name: sg13g2
.SUBCKT sg13g2_TIEH_1 vdd vss z
*.PININFO z:O vdd:B vss:B 
M_u2 net6 net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEH_2
** Cell name: TIEH_2
** Lib name: sg13g2
.SUBCKT sg13g2_TIEH_2 vdd vss z
*.PININFO z:O vdd:B vss:B 
M_u2 net6 net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEH_3
** Cell name: TIEH_3
** Lib name: sg13g2
.SUBCKT sg13g2_TIEH_3 vdd vss z
*.PININFO z:O vdd:B vss:B 
M_u2 net6 net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEH
** Cell name: TIEH
** Lib name: sg13g2
.SUBCKT sg13g2_TIEH vdd vss z
*.PININFO z:O vdd:B vss:B 
M_u2 net6 net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEL_1
** Cell name: TIEL_1
** Lib name: sg13g2
.SUBCKT sg13g2_TIEL_1 vdd vss zn
*.PININFO zn:O vdd:B vss:B 
M_u2 zn net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 net6 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEL_2
** Cell name: TIEL_2
** Lib name: sg13g2
.SUBCKT sg13g2_TIEL_2 vdd vss zn
*.PININFO zn:O vdd:B vss:B 
M_u2 zn net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 net6 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEL_3
** Cell name: TIEL_3
** Lib name: sg13g2
.SUBCKT sg13g2_TIEL_3 vdd vss zn
*.PININFO zn:O vdd:B vss:B 
M_u2 zn net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 net6 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEL
** Cell name: TIEL
** Lib name: sg13g2
.SUBCKT sg13g2_TIEL vdd vss zn
*.PININFO zn:O vdd:B vss:B 
M_u2 zn net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 net6 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.XNR2D1_1
** Cell name: XNR2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_XNR2D1_1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XNR2D1_2
** Cell name: XNR2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_XNR2D1_2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XNR2D1_3
** Cell name: XNR2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_XNR2D1_3 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XNR2D1
** Cell name: XNR2D1
** Lib name: sg13g2
.SUBCKT sg13g2_XNR2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XOR2D1_1
** Cell name: XOR2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_XOR2D1_1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XOR2D1_2
** Cell name: XOR2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_XOR2D1_2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XOR2D1_3
** Cell name: XOR2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_XOR2D1_3 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XOR2D1
** Cell name: XOR2D1
** Lib name: sg13g2
.SUBCKT sg13g2_XOR2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

************************************************************************
* Customized version of the sg13g2_io because the LVS is trash
* Put the sub pin in order to be connected to VSS later, as god intended
* It would be helpful if there is a way to check LVS with IO and pads 
* without so much trouble
************************************************************************

************************************************************************
*
* Copyright 2024 IHP PDK Authors
* 
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
*    https://www.apache.org/licenses/LICENSE-2.0
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

**ptap1 (TIE SUB)
.subckt ptap1 1 2 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
* TODO: The LVS (up to aug/28) doesnt extract correctly
*       or extracts correctly, but cannot merge/compare
*R1 1 2 R=r A=A P=Perim w=w l=l
*D1 2 1 ptap1 A=A P=Perim
.ends ptap1

**ntap1 (TIE WELL)
.subckt ntap1 1 2 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
* TODO: The LVS (up to aug/28) doesnt extract correctly
*       or extracts correctly, but cannot merge/compare
*R1 1 2 R=r A=A P=Perim w=w l=l
*D1 1 2 ntap1 A=A P=Perim
.ends ntap1

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadIOVss
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadIOVss iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
DD4 sub iovss dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD2 sub iovss dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD3 iovss iovdd dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD1 iovss iovdd dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR2 vss sub / ptap1 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
XR0 iovss sub / ptap1 r=169.45m A=5.487n Perim=296.3u w=74.075u l=74.075u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_N43N43D4R
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N43N43D4R gate pad tie sub
*.PININFO gate:I pad:B tie:B
MN0<1> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<2> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<3> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<4> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<5> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<6> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<7> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<8> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<9> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<10> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<11> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<12> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<13> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<14> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<15> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<16> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<17> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<18> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<19> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<20> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<21> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<22> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<23> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<24> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<25> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<26> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<27> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<28> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<29> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<30> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<31> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<32> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<33> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<34> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<35> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<36> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<37> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<38> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<39> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<40> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<41> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<42> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<43> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<44> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<45> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<46> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<47> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<48> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<49> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<50> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<51> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<52> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<53> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<54> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<55> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<56> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<57> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<58> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<59> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<60> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<61> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<62> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<63> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<64> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<65> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<66> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<67> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<68> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<69> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<70> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<71> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<72> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<73> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<74> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<75> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<76> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<77> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<78> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<79> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<80> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<81> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<82> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<83> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<84> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<85> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<86> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<87> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<88> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<89> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<90> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<91> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<92> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<93> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<94> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<95> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<96> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<97> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<98> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<99> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<100> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<101> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<102> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<103> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<104> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<105> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<106> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<107> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<108> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<109> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<110> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<111> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<112> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<113> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<114> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<115> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<116> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<117> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<118> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<119> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<120> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<121> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<122> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<123> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<124> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<125> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<126> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<127> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<128> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<129> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<130> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<131> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<132> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<133> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<134> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<135> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<136> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<137> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<138> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<139> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<140> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<141> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<142> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<143> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<144> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<145> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<146> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<147> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<148> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<149> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<150> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<151> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<152> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<153> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<154> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<155> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<156> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<157> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<158> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<159> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<160> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<161> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<162> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<163> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<164> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<165> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<166> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<167> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<168> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<169> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<170> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<171> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<172> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
XR0 tie sub / ptap1 r=9.999 A=65.61p Perim=32.4u w=8.1u l=8.1u
DD0 sub gate dantenna m=1 w=480n l=480n a=230.4f p=1.92u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_RCClampResistor
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_RCClampResistor pin1 pin2 sub
*.PININFO pin1:B pin2:B
R$274 pin2 pin1 rppd w=1u l=520u ps=0 b=0 m=1
*RR29 net15 net16 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR28 net20 net21 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR27 net23 net24 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR24 net17 net18 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR23 net16 net17 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR21 net25 pin2 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR20 net22 net23 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR19 net19 net20 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR17 net24 net25 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR16 net21 net22 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR15 net18 net19 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR14 net5 net6 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR13 net8 net9 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR12 net11 net12 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR11 net14 net15 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR10 net2 net3 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR9 net1 net2 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
*RR8 net13 net14 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR7 net10 net11 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR6 net7 net8 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
*RR5 net4 net5 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
*RR4 net12 net13 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR3 net9 net10 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR2 net6 net7 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
*RR1 net3 net4 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
*RR0 pin1 net1 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_RCClampInverter
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_RCClampInverter in iovss out supply sub
*.PININFO in:B iovss:B out:B supply:B
MN1 iovss in iovss sub sg13_hv_nmos m=1 w=126.000u l=9.5u ng=14
MN0 out in iovss sub sg13_hv_nmos m=1 w=108.000u l=500.0n ng=12
XR0 iovss sub / ptap1 r=9.59 A=68.973p Perim=33.22u w=8.305u l=8.305u
MP0 out in supply supply sg13_hv_pmos m=1 w=350.000u l=500.0n ng=50
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadVdd
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadVdd iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XI0 net2 vdd iovss sub / sg13g2_Clamp_N43N43D4R
XI2 vdd net1 sub / sg13g2_RCClampResistor
XR1 iovss sub / ptap1 r=456.33m A=1.97n Perim=177.54u w=44.385u l=44.385u
XR0 vss sub / ptap1 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
XI1 net1 iovss net2 vdd sub / sg13g2_RCClampInverter
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadIOVdd
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadIOVdd iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XI0 net2 iovdd iovss sub / sg13g2_Clamp_N43N43D4R
XI2 iovdd net1 sub / sg13g2_RCClampResistor
XI1 net1 iovss net2 iovdd sub / sg13g2_RCClampInverter
XR1 iovss sub / ptap1 r=449.797m A=2n Perim=178.88u w=44.72u l=44.72u
XR0 vss sub / ptap1 r=22.832 A=23.523p Perim=19.4u w=4.85u l=4.85u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_DCNDiode
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_DCNDiode anode cathode guard sub
*.PININFO anode:B cathode:B guard:B
DD1 sub cathode dantenna m=1 w=1.26u l=27.78u a=35.0028p p=58.08u
DD0 sub cathode dantenna m=1 w=1.26u l=27.78u a=35.0028p p=58.08u
*XR0 anode sub / ptap1 r=5.191 A=141.253p Perim=47.54u w=11.885u l=11.885u
XR0 anode sub / ptap1 r=5.191 A=141.2964p Perim=221.76u w=11.885u l=11.885u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_DCPDiode
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_DCPDiode anode cathode guard sub
*.PININFO anode:B cathode:B guard:B
DD1 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.0028p p=58.08u
DD0 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.0028p p=58.08u
*XR0 guard sub / ptap1 r=17.289 A=33.524p Perim=23.16u w=5.79u l=5.79u
XR0 guard sub / ptap1 r=17.289 A=33.5104p Perim=197.12u w=5.79u l=5.79u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadVss
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadVss iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XI1 iovss vss iovss sub / sg13g2_DCNDiode
XI2 vss iovdd iovss sub / sg13g2_DCPDiode
XR1 iovss sub / ptap1 r=174.346m A=5.329n Perim=292u w=73u l=73u
XR0 vss sub / ptap1 r=22.832 A=23.523p Perim=19.4u w=4.85u l=4.85u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler4000
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler4000 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=63.078 A=5.856p Perim=9.68u w=2.42u l=2.42u
XR0 iovss sub / ptap1 r=625.742m A=1.416n Perim=150.5u w=37.625u l=37.625u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_io_inv_x1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_inv_x1 i nq vdd vss sub
*.PININFO i:I nq:O vdd:B vss:B
MN0 nq i vss sub sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MP0 nq i vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
XR0 vss sub / ptap1 r=258.978 A=624.1f Perim=3.16u w=790n l=790n
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_LevelUp
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_LevelUp i iovdd o vdd vss sub
*.PININFO i:I o:O iovdd:B vdd:B vss:B
MN0 net2 i vss sub sg13_lv_nmos m=1 w=2.75u l=130.00n ng=1
MP0 net2 i vdd vdd sg13_lv_pmos m=1 w=4.75u l=130.00n ng=1
MN3 o net4 vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN2 net4 i vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN1 net3 net2 vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MP3 o net4 iovdd iovdd sg13_hv_pmos m=1 w=3.9u l=450.00n ng=1
MP2 net3 net4 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
MP1 net4 net3 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
XR0 vss sub / ptap1 r=207.099 A=912.025f Perim=3.82u w=955n l=955n
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_io_nor2_x1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_nor2_x1 i0 i1 nq vdd vss sub
*.PININFO i0:I i1:I nq:O vdd:B vss:B
MN0 nq i0 vss sub sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MN1 nq i1 vss sub sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MP1 net1 i0 vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
MP0 nq i1 net1 vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
XR0 vss sub / ptap1 r=251.534 A=656.1f Perim=3.24u w=810n l=810n
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_io_tie
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_tie vdd vss sub
*.PININFO vdd:B vss:B
XR0 vss sub / ptap1 r=258.978 A=624.1f Perim=3.16u w=790n l=790n
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_io_nand2_x1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_nand2_x1 i0 i1 nq vdd vss sub
*.PININFO i0:I i1:I nq:O vdd:B vss:B
MP1 nq i1 vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
MP0 nq i0 vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
MN1 net1 i0 vss sub sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MN0 nq i1 net1 sub sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
XR0 vss sub / ptap1 r=251.534 A=656.1f Perim=3.24u w=810n l=810n
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_GateDecode
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_GateDecode core en iovdd ngate pgate vdd vss sub
*.PININFO core:I en:I ngate:O pgate:O iovdd:B vdd:B vss:B
XI2 en net3 vdd vss sub / sg13g2_io_inv_x1
XI4 net4 iovdd ngate vdd vss sub / sg13g2_LevelUp
XI3 net2 iovdd pgate vdd vss sub / sg13g2_LevelUp
XI0 core net3 net4 vdd vss sub / sg13g2_io_nor2_x1
XI5 vdd vss sub / sg13g2_io_tie
XI1 core en net2 vdd vss sub / sg13g2_io_nand2_x1
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_N2N2D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N2N2D gate iovss pad sub
*.PININFO gate:B iovss:B pad:B
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
MN1 iovss gate pad sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0 pad gate iovss sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
DD0 sub gate dantenna m=1 w=780.00n l=780.00n a=608.400f p=3.12u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_P2N2D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_P2N2D gate iovdd iovss pad sub
*.PININFO gate:B iovdd:B iovss:B pad:B
DD0 gate iovdd dpantenna m=1 w=480n l=480n a=230.4f p=1.92u
MP1 iovdd gate pad iovdd sg13_hv_pmos m=1 w=13.32u l=600.0n ng=2
MP0 pad gate iovdd iovdd sg13_hv_pmos m=1 w=13.32u l=600.0n ng=2
XR0 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_SecondaryProtection
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_SecondaryProtection core minus pad plus sub
*.PININFO core:B minus:B pad:B plus:B
*RR0 pad core 586.899 $SUB=sub $[res_rppd] m=1 l=2u w=1u ps=180n trise=0.0 b=0
RR0 pad core rppd m=1 l=2u w=1u
DD0 sub core dantenna m=1 w=640n l=3.1u a=1.984p p=7.48u
*XR1 minus sub / ptap1 r=46.556 A=9.03p Perim=12.02u w=3.005u l=3.005u
XR1 minus sub / ptap1 r=46.556 A=9.0304p Perim=53.12u w=3.005u l=3.005u
DD1 core plus dpantenna m=1 w=640n l=4.98u a=3.187p p=11.24u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_LevelDown
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_LevelDown core iovdd iovss pad vdd vss sub
*.PININFO core:O iovdd:B iovss:B pad:B vdd:B vss:B
MP0 net2 net4 vdd vdd sg13_hv_pmos m=1 w=4.65u l=450.00n ng=1
MN0 net2 net4 vss sub sg13_hv_nmos m=1 w=2.65u l=450.00n ng=1
MN1 core net2 vss sub sg13_lv_nmos m=1 w=2.75u l=130.00n ng=1
MP1 core net2 vdd vdd sg13_lv_pmos m=1 w=4.75u l=130.00n ng=1
*XR0 vss sub / ptap1 r=127.332 A=2.016p Perim=5.68u w=1.42u l=1.42u
XR0 vss sub / ptap1 r=127.332 A=2.019p Perim=14.06u w=1.42u l=1.42u
XI0 net4 iovss pad iovdd sub / sg13g2_SecondaryProtection
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadInOut4mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadInOut4mA c2p c2p_en iovdd iovss p2c pad vdd vss sub
*.PININFO c2p:I c2p_en:I p2c:O iovdd:B iovss:B pad:B vdd:B vss:B
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XI0 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
XI7 net2 iovss pad sub / sg13g2_Clamp_N2N2D
XI6 net1 iovdd iovss pad sub / sg13g2_Clamp_P2N2D
XI1 p2c iovdd iovss pad vdd vss sub / sg13g2_LevelDown
XR1 vss sub / ptap1 r=26.933 A=18.966p Perim=17.42u w=4.355u l=4.355u
XR0 iovss sub / ptap1 r=214.134m A=4.314n Perim=262.72u w=65.68u l=65.68u
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_P15N15D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_P15N15D gate iovdd iovss pad sub
*.PININFO gate:B iovdd:B iovss:B pad:B
DD0 gate iovdd dpantenna m=1 w=780.00n l=780.00n a=608.400f p=3.12u
XR0 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
MP1 pad gate iovdd iovdd sg13_hv_pmos m=1 w=199.8u l=600.0n ng=30
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_N15N15D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N15N15D gate iovss pad sub
*.PININFO gate:B iovss:B pad:B
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
MN0 pad gate iovss sub sg13_hv_nmos m=1 w=66.000u l=600.0n ng=15
DD0 sub gate dantenna m=1 w=780.00n l=780.00n a=608.400f p=3.12u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadInOut30mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadInOut30mA c2p c2p_en iovdd iovss p2c pad vdd vss sub
*.PININFO c2p:I c2p_en:I p2c:O iovdd:B iovss:B pad:B vdd:B vss:B
XI1 p2c iovdd iovss pad vdd vss sub / sg13g2_LevelDown
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XI7 net1 iovdd iovss pad sub / sg13g2_Clamp_P15N15D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI6 net2 iovss pad sub / sg13g2_Clamp_N15N15D
XR4 vss sub / ptap1 r=26.746 A=19.141p Perim=17.5u w=4.375u l=4.375u
XR3 iovss sub / ptap1 r=214.165m A=4.313n Perim=262.7u w=65.675u l=65.675u
XI0 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_LevelUpInv
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_LevelUpInv i iovdd o vdd vss sub
*.PININFO i:I o:O iovdd:B vdd:B vss:B
MN0 net2 i vss sub sg13_lv_nmos m=1 w=2.75u l=130.00n ng=1
MP0 net2 i vdd vdd sg13_lv_pmos m=1 w=4.75u l=130.00n ng=1
MN3 o net4 vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN2 net4 net2 vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN1 net3 i vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MP3 o net4 iovdd iovdd sg13_hv_pmos m=1 w=3.9u l=450.00n ng=1
MP2 net3 net4 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
MP1 net4 net3 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
XR0 vss sub / ptap1 r=190.268 A=1.051p Perim=4.1u w=1.025u l=1.025u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_GateLevelUpInv
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_GateLevelUpInv core iovdd ngate pgate vdd vss sub
*.PININFO core:I ngate:O pgate:O iovdd:B vdd:B vss:B
XI1 core iovdd pgate vdd vss sub / sg13g2_LevelUpInv
XI0 core iovdd ngate vdd vss sub / sg13g2_LevelUpInv
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadOut4mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadOut4mA c2p iovdd iovss pad vdd vss sub
*.PININFO c2p:I iovdd:B iovss:B pad:B vdd:B vss:B
XI6 c2p iovdd net2 net1 vdd vss sub / sg13g2_GateLevelUpInv
XI7 net1 iovdd iovss pad sub / sg13g2_Clamp_P2N2D
XI8 net2 iovss pad sub / sg13g2_Clamp_N2N2D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR2 iovss sub / ptap1 r=212.747m A=4.343n Perim=263.6u w=65.9u l=65.9u
XR1 vss sub / ptap1 r=24.125 A=21.902p Perim=18.72u w=4.68u l=4.68u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadOut30mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadOut30mA c2p iovdd iovss pad vdd vss sub
*.PININFO c2p:I iovdd:B iovss:B pad:B vdd:B vss:B
XI6 c2p iovdd net2 net1 vdd vss sub / sg13g2_GateLevelUpInv
XI7 net1 iovdd iovss pad sub / sg13g2_Clamp_P15N15D
XI8 net2 iovss pad sub / sg13g2_Clamp_N15N15D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR1 vss sub / ptap1 r=24.125 A=21.902p Perim=18.72u w=4.68u l=4.68u
XR2 iovss sub / ptap1 r=214.165m A=4.313n Perim=262.7u w=65.675u l=65.675u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadIn
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadIn iovdd iovss p2c pad vdd vss sub
.PININFO p2c:O iovdd:B iovss:B pad:B vdd:B vss:B
XI1 p2c iovdd iovss pad vdd vss sub / sg13g2_LevelDown
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
*XR1 vss sub / ptap1 r=24.69 A=21.252p Perim=18.44u w=4.61u l=4.61u
*XR2 iovss sub / ptap1 r=173.674m A=5.35n Perim=292.58u w=73.145u l=73.145u
XR1 vss sub / ptap1 r=24.69 A=21.981p Perim=107.48u w=4.61u l=4.61u
XR2 iovss sub / ptap1 r=173.674m A=5223.2628p Perim=221.16u w=73.145u l=73.145u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_P8N8D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_P8N8D gate iovdd iovss pad sub
*.PININFO gate:B iovdd:B iovss:B pad:B
XR0 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
MP0 pad gate iovdd iovdd sg13_hv_pmos m=1 w=106.56u l=600.0n ng=16
DD0 gate iovdd dpantenna m=1 w=480n l=480n a=230.4f p=1.92u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_N8N8D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N8N8D gate iovss pad sub
*.PININFO gate:B iovss:B pad:B
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
MN0 pad gate iovss sub sg13_hv_nmos m=1 w=35.2u l=600.0n ng=8
DD0 sub gate dantenna m=1 w=780.00n l=780.00n a=608.400f p=3.12u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadInOut16mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadInOut16mA c2p c2p_en iovdd iovss p2c pad vdd vss sub
*.PININFO c2p:I c2p_en:I p2c:O iovdd:B iovss:B pad:B vdd:B vss:B
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XI0 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI7 net1 iovdd iovss pad sub / sg13g2_Clamp_P8N8D
XI1 p2c iovdd iovss pad vdd vss sub / sg13g2_LevelDown
XI6 net2 iovss pad sub / sg13g2_Clamp_N8N8D
XR1 vss sub / ptap1 r=26.933 A=18.966p Perim=17.42u w=4.355u l=4.355u
XR0 iovss sub / ptap1 r=207.756m A=4.45n Perim=266.84u w=66.71u l=66.71u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadOut16mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadOut16mA c2p iovdd iovss pad vdd vss sub
*.PININFO c2p:I iovdd:B iovss:B pad:B vdd:B vss:B
* TODO: AGAIN?!?!?!
*XI6 c2p iovdda net2 net1 vdd vss sub / sg13g2_GateLevelUpInv
XI6 c2p iovdd net2 net1 vdd vss sub / sg13g2_GateLevelUpInv
XI8 net1 iovdd iovss pad sub / sg13g2_Clamp_P8N8D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI7 net2 iovss pad sub / sg13g2_Clamp_N8N8D
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR1 vss sub / ptap1 r=23.888 A=22.184p Perim=18.84u w=4.71u l=4.71u
XR2 iovss sub / ptap1 r=208.667m A=4.43n Perim=266.24u w=66.56u l=66.56u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadTriOut4mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadTriOut4mA c2p c2p_en iovdd iovss pad vdd vss sub
*.PININFO c2p:I c2p_en:I iovdd:B iovss:B pad:B vdd:B vss:B
XI7 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI8 net2 iovss pad sub / sg13g2_Clamp_N2N2D
XI9 net1 iovdd iovss pad sub / sg13g2_Clamp_P2N2D
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR1 vss sub / ptap1 r=24.567 A=21.391p Perim=18.5u w=4.625u l=4.625u
XR2 iovss sub / ptap1 r=208.667m A=4.43n Perim=266.24u w=66.56u l=66.56u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadTriOut16mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadTriOut16mA c2p c2p_en iovdd iovss pad vdd vss sub
*.PININFO c2p:I c2p_en:I iovdd:B iovss:B pad:B vdd:B vss:B
XI7 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
XI8 net1 iovdd iovss pad sub / sg13g2_Clamp_P8N8D
XI9 net2 iovss pad sub / sg13g2_Clamp_N8N8D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR1 vss sub / ptap1 r=24.897 A=21.022p Perim=18.34u w=4.585u l=4.585u
XR2 iovss sub / ptap1 r=208.211m A=4.44n Perim=266.54u w=66.635u l=66.635u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadTriOut30mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadTriOut30mA c2p c2p_en iovdd iovss pad vdd vss sub
*.PININFO c2p:I c2p_en:I iovdd:B iovss:B pad:B vdd:B vss:B
XI7 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI8 net2 iovss pad sub / sg13g2_Clamp_N15N15D
XI9 net1 iovdd iovss pad sub / sg13g2_Clamp_P15N15D
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR1 vss sub / ptap1 r=24.649 A=21.298p Perim=18.46u w=4.615u l=4.615u
XR2 iovss sub / ptap1 r=208.667m A=4.43n Perim=266.24u w=66.56u l=66.56u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Corner
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Corner iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=35.383 A=13.177p Perim=14.52u w=3.63u l=3.63u
XR0 iovss sub / ptap1 r=93.041m A=10.13n Perim=402.6u w=100.65u l=100.65u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler400
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler400 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=246.192 A=680.625f Perim=3.3u w=825n l=825n
XR0 iovss sub / ptap1 r=6.246 A=114.169p Perim=42.74u w=10.685u l=10.685u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler200
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler200 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=246.192 A=680.625f Perim=3.3u w=825n l=825n
XR0 iovss sub / ptap1 r=14.724 A=40.96p Perim=25.6u w=6.4u l=6.4u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler1000
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler1000 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=162.013 A=1.369p Perim=4.68u w=1.17u l=1.17u
XR0 iovss sub / ptap1 r=2.443 A=328.697p Perim=72.52u w=18.13u l=18.13u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler2000
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler2000 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=101.912 A=2.856p Perim=6.76u w=1.69u l=1.69u
XR0 iovss sub / ptap1 r=1.224 A=695.113p Perim=105.46u w=26.365u l=26.365u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler10000
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler10000 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=32.364 A=14.861p Perim=15.42u w=3.855u l=3.855u
XR0 iovss sub / ptap1 r=253.731m A=3.622n Perim=240.72u w=60.18u l=60.18u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_P20N0D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_P20N0D iovdd iovss pad sub
*.PININFO iovdd:B iovss:B pad:B
MP0 pad net2 iovdd iovdd sg13_hv_pmos m=1 w=266.4u l=600.0n ng=40
*RR0 net2 iovdd 6.768K $SUB=iovdd $[res_rppd] m=1 l=12.9u w=500n ps=180n 
+ trise=0.0 b=0
RR0 iovdd net2 rppd m=1 l=12.9u w=500n
+ trise=0.0 b=0
XR1 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_N20N0D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N20N0D iovss pad sub
*.PININFO iovss:B pad:B
MN0 pad net2 iovss sub sg13_hv_nmos m=1 w=88.000u l=600.0n ng=20
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
*RR1 iovss net2 1.959K $SUB=sub $[res_rppd] m=1 l=3.54u w=500n ps=180n 
+ trise=0.0 b=0
RR1 iovss net2 rppd m=1 l=3.54u w=500n
+ trise=0.0 b=0
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadAnalog
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadAnalog iovdd iovss pad padres vdd vss sub
*.PININFO iovdd:B iovss:B pad:B padres:B vdd:B vss:B
XI9 iovdd iovss pad sub / sg13g2_Clamp_P20N0D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
*** WHYYYYYY. Lets put it like that for now. My god this is annoying
*XI6 padres iovss pad iovdda sub / sg13g2_SecondaryProtection
XI6 padres iovss pad iovdd sub / sg13g2_SecondaryProtection
XI8 iovss pad sub / sg13g2_Clamp_N20N0D
XR1 vss sub / ptap1 r=22.579 A=23.863p Perim=19.54u w=4.885u l=4.885u
XR2 iovss sub / ptap1 r=214.8m A=4.3n Perim=262.3u w=65.575u l=65.575u
.ENDS
.SUBCKT sg13g2_bpd60
.ENDS

.SUBCKT sg13g2_bpd70
.ENDS

.SUBCKT sg13g2_bpd80
.ENDS
*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

.SUBCKT sg13g2_Clamp_N20N0DExt iovss pad sub
*.PININFO iovss:B pad:B
MN0 pad net2 iovss sub sg13_hv_nmos m=1 w=88.000u l=600.0n ng=20
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
*RR1 iovss net2 1.959K $SUB=sub $[res_rppd] m=1 l=3.54u w=500n ps=180n 
+ trise=0.0 b=0
*RR0 net2 iovdd 6.768K $SUB=iovdd $[res_rppd] m=1 l=12.9u w=500n ps=180n 
+ trise=0.0 b=0
RR0 iovdd net2 rppd m=1 l=12.9u w=500n
+ trise=0.0 b=0
.ENDS

.SUBCKT sg13g2_SecondaryProtectionExt core minus pad plus sub
*.PININFO core:B minus:B pad:B plus:B
*RR0 pad core 586.899 $SUB=sub $[res_rppd] m=1 l=2u w=1u ps=180n trise=0.0 b=0
RR0 pad core rppd m=1 l=2u w=1u
DD0 sub core dantenna m=1 w=640n l=3.1u a=1.984p p=7.48u
XR1 minus sub / ptap1 r=46.556 A=9.03p Perim=12.02u w=3.005u l=3.005u
DD1 core plus dpantenna m=1 w=640n l=4.98u a=3.187p p=11.24u
.ENDS

.SUBCKT sg13g2_Clamp_P20N0DExt iovdd iovss pad sub
*.PININFO iovdd:B iovss:B pad:B
MP0 pad net2 iovdd iovdd sg13_hv_pmos m=1 w=266.4u l=600.0n ng=40
RR0 net2 iovdd 6.768K $SUB=iovdd $[res_rppd] m=1 l=12.9u w=500n ps=180n 
+ trise=0.0 b=0
XR1 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
.ENDS

.SUBCKT sg13g2_RCClampInverterExt in iovss out supply sub
*.PININFO in:B iovss:B out:B supply:B
MN1 iovss in iovss sub sg13_hv_nmos m=1 w=126.000u l=9.5u ng=14
MN0 out in iovss sub sg13_hv_nmos m=1 w=108.000u l=500.0n ng=12
XR0 iovss sub / ptap1 r=9.59 A=68.973p Perim=33.22u w=8.305u l=8.305u
MP0 out in supply supply sg13_hv_pmos m=1 w=350.000u l=500.0n ng=50
.ENDS

.SUBCKT sg13g2_RCClampResistorExt pin1 pin2 sub
*.PININFO pin1:B pin2:B
R$274 pin2 pin1 rppd w=1u l=520u ps=0 b=0 m=1
.ENDS

.SUBCKT sg13g2_RCClampResistorExt_Orig pin1 pin2 sub
*.PININFO pin1:B pin2:B
RR29 net15 net16 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR28 net20 net21 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR27 net23 net24 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR24 net17 net18 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR23 net16 net17 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR21 net25 pin2 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR20 net22 net23 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR19 net19 net20 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR17 net24 net25 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR16 net21 net22 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR15 net18 net19 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR14 net5 net6 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR13 net8 net9 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR12 net11 net12 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR11 net14 net15 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR10 net2 net3 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR9 net1 net2 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR8 net13 net14 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR7 net10 net11 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR6 net7 net8 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR5 net4 net5 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR4 net12 net13 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR3 net9 net10 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR2 net6 net7 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR1 net3 net4 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR0 pin1 net1 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
.ENDS

.SUBCKT sg13g2_Clamp_N43N43D4RExt gate pad tie sub
*.PININFO gate:I pad:B tie:B
MN0<1> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<2> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<3> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<4> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<5> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<6> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<7> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<8> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<9> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<10> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<11> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<12> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<13> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<14> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<15> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<16> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<17> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<18> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<19> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<20> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<21> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<22> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<23> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<24> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<25> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<26> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<27> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<28> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<29> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<30> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<31> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<32> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<33> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<34> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<35> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<36> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<37> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<38> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<39> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<40> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<41> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<42> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<43> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<44> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<45> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<46> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<47> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<48> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<49> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<50> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<51> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<52> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<53> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<54> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<55> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<56> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<57> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<58> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<59> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<60> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<61> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<62> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<63> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<64> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<65> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<66> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<67> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<68> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<69> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<70> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<71> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<72> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<73> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<74> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<75> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<76> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<77> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<78> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<79> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<80> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<81> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<82> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<83> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<84> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<85> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<86> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<87> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<88> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<89> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<90> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<91> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<92> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<93> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<94> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<95> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<96> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<97> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<98> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<99> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<100> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<101> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<102> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<103> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<104> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<105> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<106> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<107> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<108> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<109> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<110> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<111> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<112> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<113> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<114> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<115> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<116> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<117> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<118> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<119> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<120> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<121> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<122> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<123> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<124> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<125> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<126> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<127> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<128> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<129> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<130> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<131> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<132> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<133> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<134> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<135> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<136> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<137> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<138> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<139> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<140> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<141> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<142> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<143> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<144> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<145> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<146> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<147> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<148> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<149> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<150> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<151> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<152> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<153> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<154> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<155> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<156> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<157> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<158> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<159> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<160> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<161> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<162> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<163> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<164> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<165> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<166> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<167> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<168> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<169> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<170> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<171> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<172> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
XR0 tie sub / ptap1 r=9.999 A=65.61p Perim=32.4u w=8.1u l=8.1u
DD0 sub gate dantenna m=1 w=480n l=480n a=230.4f p=1.92u
.ENDS

.SUBCKT sg13g2_DCNDiodeExt anode cathode guard sub
*.PININFO anode:B cathode:B guard:B
DD1 sub cathode dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD0 sub cathode dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR0 anode sub / ptap1 r=5.191 A=141.253p Perim=47.54u w=11.885u l=11.885u
.ENDS

.SUBCKT sg13g2_DCPDiodeExt anode cathode guard sub
*.PININFO anode:B cathode:B guard:B
DD1 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD0 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR0 guard sub / ptap1 r=17.289 A=33.524p Perim=23.16u w=5.79u l=5.79u
.ENDS

.SUBCKT sg13g2_IOPadVssExt iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XI1 iovss vss iovss sub / sg13g2_DCNDiodeExt
XI2 vss iovdd iovss sub / sg13g2_DCPDiodeExt
XR1 iovss sub / ptap1 r=174.346m A=5.329n Perim=292u w=73u l=73u
XR0 vss sub / ptap1 r=22.832 A=23.523p Perim=19.4u w=4.85u l=4.85u
.ENDS

.SUBCKT sg13g2_IOPadVddExt iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
* OHH MY GOD
*XI0 net2 vdd iovssa sub / sg13g2_Clamp_N43N43D4RExt
XI0 net2 vdd iovss sub / sg13g2_Clamp_N43N43D4RExt
XI2 vdd net1 sub / sg13g2_RCClampResistorExt
XR1 iovss sub / ptap1 r=456.33m A=1.97n Perim=177.54u w=44.385u l=44.385u
XR0 vss sub / ptap1 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
XI1 net1 iovss net2 vdd sub  / sg13g2_RCClampInverterExt
.ENDS

.SUBCKT sg13g2_IOPadAVDD iovdd iovss pad padres vdd vss sub
*.PININFO iovdd:B iovss:B pad:B padres:B vdd:B vss:B
XI9 iovdd iovss pad sub / sg13g2_Clamp_P20N0DExt
XI3 iovss pad iovdd sub / sg13g2_DCNDiodeExt
XI2 pad iovdd iovss sub / sg13g2_DCPDiodeExt
XI6 padres iovss pad iovdd sub / sg13g2_SecondaryProtectionExt
XI8 iovss pad sub / sg13g2_Clamp_N20N0DExt
XR1 vss sub / ptap1 r=22.579 A=23.863p Perim=19.54u w=4.885u l=4.885u
XR2 iovss sub / ptap1 r=214.8m A=4.3n Perim=262.3u w=65.575u l=65.575u
.ENDS
.SUBCKT sealring
.ENDS
** Created by: circuit_gen.AN2D0
** Cell name: AN2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_AN2D0 a1 a2 vdd vss z
*.PININFO a1:B a2:B vdd:B vss:B z:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.AN2D1
** Cell name: AN2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_AN2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=6.550e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.550e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.AN2D2
** Cell name: AN2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_AN2D2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net10 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_M_u2_0 z net10 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_M_u2_1 z net10 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_M_u3_0 z net10 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_M_u3_1 z net10 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_M_u2 net10 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_M_u1 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.AN2D4
** Cell name: AN2D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_AN2D4 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_0_M_u3 p0 a1 x_u2_0_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_0_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_1_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_2_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_3_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_0_M_u4 x_u2_0_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_1_M_u4 x_u2_1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_1_M_u3 p0 a1 x_u2_1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_0_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_1_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_2_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_3_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_0_M_u2 p0 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_0_M_u1 p0 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_1_M_u2 p0 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_1_M_u1 p0 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.AO21D0
** Cell name: AO21D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_AO21D0 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.AO21D1
** Cell name: AO21D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_AO21D1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.AO21D2
** Cell name: AO21D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_AO21D2 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_0_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_1_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_0_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_1_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.AOI21D0
** Cell name: AOI21D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_AOI21D0 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI7 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI6 zn b vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI5 zn a2 net13 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI4 zn a1 net13 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.AOI21D1
** Cell name: AOI21D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_AOI21D1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI3 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u7 zn b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u4 net13 a2 zn vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3 net13 a1 zn vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ANTENNA
** Cell name: ANTENNA
** Lib name: sg13g2f
.SUBCKT sg13g2f_ANTENNA i vdd vss
*.PININFO i:I vdd:B vss:B
Ddn_1 vss i dantenna m=1 w=1.485u l=970n a=1440.45f
DD0 i vdd dpantenna m=1 w=1.485u l=970n a=1440.45f
.ENDS

** Created by: circuit_gen.BUFFD0
** Cell name: BUFFD0
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD0 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
M_u2_M_u2 net6 i vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.850e-07
M_u2_M_u3 net6 i vdd vdd sg13_lv_pmos l=1.300e-07 w=3.600e-07
.ENDS

** Created by: circuit_gen.BUFFD1
** Cell name: BUFFD1
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD1 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.BUFFD2
** Cell name: BUFFD2
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD2 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_0_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_1_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_0_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_1_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.BUFFD4
** Cell name: BUFFD4
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD4 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_0_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_1_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_2_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_3_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_0_M_u2 p0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_1_M_u2 p0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_0_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_1_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_2_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_3_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_0_M_u3 p0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_1_M_u3 p0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.BUFFD6
** Cell name: BUFFD6
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD6 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u2_M_u2_0 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=1
M_u2_M_u2_1 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=0
M_u3_0_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
M_u3_1_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=0
M_u3_2_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=1
M_u3_3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=0
M_u3_4_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=1
M_u3_5_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=0
M_u2_M_u3_0 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=1
M_u2_M_u3_1 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=0
M_u3_0_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=1
M_u3_1_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
M_u3_2_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=1
M_u3_3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=0
M_u3_4_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=1
M_u3_5_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=0
.ENDS

** Created by: circuit_gen.BUFFD8
** Cell name: BUFFD8
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD8 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI1_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MI2_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.850e-07 $pos=1 $flip=1
M_u2_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
M_u7_0_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
M_u7_1_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
M_u7_2_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
M_u7_3_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
M_u7_4_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
M_u7_5_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=0
M_u7_6_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
M_u7_7_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MI1_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MI2_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=8.050e-07 $pos=1 $flip=1
M_u2_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
M_u7_0_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
M_u7_1_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
M_u7_2_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
M_u7_3_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
M_u7_4_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
M_u7_5_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
M_u7_6_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
M_u7_7_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
.ENDS

** Created by: circuit_gen.BUFFD12
** Cell name: BUFFD12
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD12 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u2_0_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=0 $flip=0
M_u2_1_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=1 $flip=1
M_u2_2_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=2 $flip=0
M_u2_3_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=3 $flip=1
M_u2_4_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=4 $flip=0
MU8_0_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU8_1_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MU8_2_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MU8_3_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=0
MU8_4_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MU8_5_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MU8_6_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=1
MU8_7_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=12 $flip=0
MU8_8_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=13 $flip=1
MU8_9_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=14 $flip=0
MU8_10_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=15 $flip=1
MU8_11_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=16 $flip=0
M_u2_0_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
M_u2_1_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
M_u2_2_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
M_u2_3_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
M_u2_4_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU8_0_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MU8_1_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MU8_2_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MU8_3_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
MU8_4_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
MU8_5_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
MU8_6_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
MU8_7_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=0
MU8_8_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=13 $flip=1
MU8_9_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=14 $flip=0
MU8_10_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=15 $flip=1
MU8_11_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=16 $flip=0
.ENDS

** Created by: circuit_gen.BUFFD16
** Cell name: BUFFD16
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD16 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI6_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07 $pos=0 $flip=1
M_u2_0_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=0
M_u2_1_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
M_u2_2_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=0
M_u2_3_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=1
M_u2_4_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=0
MU8_0_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=1
MU8_1_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=0
MU8_2_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=1
MU8_3_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=0
MU8_4_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=1
MU8_5_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=0
MU8_6_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=12 $flip=1
MU8_7_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=13 $flip=0
MU8_8_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=14 $flip=1
MU8_9_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=15 $flip=0
MU8_10_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=16 $flip=1
MU8_11_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=17 $flip=0
MU8_12_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=18 $flip=1
MU8_13_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=19 $flip=0
MU8_14_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=20 $flip=1
MU8_15_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=21 $flip=0
MI6_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=3.950e-07 $pos=0 $flip=1
M_u2_0_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=0
M_u2_1_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=1
M_u2_2_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
M_u2_3_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=1
M_u2_4_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=0
MU8_0_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=1
MU8_1_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=0
MU8_2_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=1
MU8_3_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=0
MU8_4_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=1
MU8_5_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=0
MU8_6_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=1
MU8_7_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=13 $flip=0
MU8_8_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=14 $flip=1
MU8_9_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=15 $flip=0
MU8_10_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=16 $flip=1
MU8_11_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=17 $flip=0
MU8_12_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=18 $flip=1
MU8_13_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=19 $flip=0
MU8_14_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=20 $flip=1
MU8_15_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=21 $flip=0
.ENDS

** Created by: circuit_gen.DEL0
** Cell name: DEL0
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL0 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI2_M_u2 z net3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU7_M_u2 net3 net5 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU5_M_u2 net5 net9 vss vss sg13_lv_nmos l=1.300e-07 w=4.800e-07
MI1_M_u2 net9 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI2_M_u3 z net3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU7_M_u3 net3 net5 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.040e-06
MU5_M_u3 net5 net9 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u3 net9 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DEL2
** Cell name: DEL2
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL2 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI2_M_u2 z net3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU7_M_u2 net3 net5 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU5_M_u2 net5 net9 vss vss sg13_lv_nmos l=1.300e-07 w=4.800e-07
MI1_M_u2 net9 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI2_M_u3 z net3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU7_M_u3 net3 net5 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.000e-07
MU5_M_u3 net5 net9 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u3 net9 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DEL02
** Cell name: DEL02
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL02 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI17 net3 net21 net27 vss sg13_lv_nmos l=1.300e-07 w=3.350e-07
MI18 net27 net21 vss vss sg13_lv_nmos l=1.300e-07 w=3.350e-07
MI5 net21 net9 net24 vss sg13_lv_nmos l=1.300e-07 w=3.350e-07
MI16 net24 net9 vss vss sg13_lv_nmos l=1.300e-07 w=3.350e-07
MI2_M_u2 z net3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u2 net9 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI15 net27 net21 net3 vdd sg13_lv_pmos l=1.300e-07 w=5.650e-07
MI13 net24 net9 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.650e-07
MI3 vdd net9 net24 vdd sg13_lv_pmos l=1.300e-07 w=5.650e-07
MI14 vdd net21 net27 vdd sg13_lv_pmos l=1.300e-07 w=5.650e-07
MI2_M_u3 z net3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u3 net9 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DEL4
** Cell name: DEL4
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL4 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI2_M_u2 z net13 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU7_M_u2 net13 net11 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU5_M_u2 net11 net9 vss vss sg13_lv_nmos l=1.300e-07 w=4.800e-07
MI1_M_u2 net9 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI2_M_u3 z net13 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU7_M_u3 net13 net11 vdd vdd sg13_lv_pmos l=1.300e-07 w=8.500e-07
MU5_M_u3 net11 net9 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u3 net9 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DEL005
** Cell name: DEL005
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL005 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI12 net3 i net22 vss sg13_lv_nmos l=1.300e-07 w=4.250e-07
MI13 net22 i vss vss sg13_lv_nmos l=1.300e-07 w=4.250e-07
MI2_M_u2 z net3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI10 net3 i net21 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI3 net21 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI2_M_u3 z net3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DEL015
** Cell name: DEL015
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL015 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI11 net27 net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI10 net3 net21 net27 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI5 net21 net9 net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI111 net24 net9 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI2_M_u2 z net3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u2 net9 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8 net27 net21 net3 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI9 vdd net21 net27 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI4 net24 net9 net21 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI3 vdd net9 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI2_M_u3 z net3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u3 net9 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DFCNQD1
** Cell name: DFCNQD1
** Lib name: sg13g2
.SUBCKT sg13g2f_DFCNQD1 cdn cp d q vdd vss
*.PININFO cdn:I cp:I d:I q:O vdd:B vss:B 
Mcpbn incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=0 $flip=0
Mcpbp incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07 $pos=0 $flip=0
Mcpn incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=1 $flip=1
Mcpp incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07 $pos=1 $flip=1
MI4 net52 incpb vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=3 $flip=1
MI7 net85 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07 $pos=3 $flip=1
Mdd0n d0 d net52 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=4 $flip=1
Mdd0p d0 d net85 vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07 $pos=4 $flip=1
MI47 d0 incp net59 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=5 $flip=0
MI45 d0 incpb net98 vdd sg13_lv_pmos l=1.300e-07 w=3.300e-07 $pos=5 $flip=0
MI48 net59 d1 net62 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=6 $flip=0
MI43 net98 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=3.050e-07 $pos=6 $flip=0
Mcdn0n net62 cdn vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=7 $flip=0
Md0d1n d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=8 $flip=1
Mcdn0p net98 cdn vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=8 $flip=0
Mswd1d2n d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=4.900e-07 $pos=9 $flip=0
Mdod1p d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.150e-07 $pos=9 $flip=1
MI23 d2 incpb net57 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=10 $flip=0
Mswd1d2p d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=1.030e-06 $pos=10 $flip=0
MI26 d2 incp net88 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=11 $flip=0
MI24 net57 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=12 $flip=0
MI28 net88 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=12 $flip=0
Mcdn1n net37 cdn vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=13 $flip=1
Mcdn1p d3 cdn vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07 $pos=13 $flip=1
Md2d3n d3 d2 net37 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=14 $flip=1
Md2d3p d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07 $pos=14 $flip=0
Mobp q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06 $pos=15 $flip=1
Mobn q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=16 $flip=1
.ENDS

** Created by: circuit_gen.DFQD1
** Cell name: DFQD1
** Lib name: sg13g2f
.SUBCKT sg13g2f_DFQD1 cp d q vdd vss
*.PININFO cp:I d:I q:O vdd:B vss:B 
MI4 net43 incpb vss vss sg13_lv_nmos l=1.300e-07 w=4.200e-07
MI23 d2 incpb net42 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI5 d0 d net43 vss sg13_lv_nmos l=1.300e-07 w=4.200e-07
MI47 d0 incp net50 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI48 net50 d1 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI24 net42 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI50 d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=3.850e-07
MI32_M_u2 incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI31_M_u2 incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI27_M_u2 q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI53_M_u2 d3 d2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI13_M_u2 d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.700e-07
MI6 d0 d net66 vdd sg13_lv_pmos l=1.300e-07 w=7.500e-07
MI32_M_u3 incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI31_M_u3 incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI27_M_u3 q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI53_M_u3 d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI13_M_u3 d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.500e-07
MI7 net66 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.850e-07
MI52 d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=1.065e-06
MI28 net74 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=3.000e-07
MI26 d2 incp net74 vdd sg13_lv_pmos l=1.300e-07 w=3.000e-07
MI45 d0 incpb net84 vdd sg13_lv_pmos l=1.300e-07 w=3.000e-07
MI43 net84 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=3.000e-07
.ENDS

** Created by: circuit_gen.FILL1
** Cell name: FILL1
** Lib name: sg13g2f
.SUBCKT sg13g2f_FILL1 vdd vss
*.PININFO vdd:B vss:B 
.ENDS

** Created by: circuit_gen.FILL2
** Cell name: FILL2
** Lib name: sg13g2f
.SUBCKT sg13g2f_FILL2 vdd vss
*.PININFO vdd:B vss:B 
.ENDS

** Created by: circuit_gen.FILL4
** Cell name: FILL4
** Lib name: sg13g2f
.SUBCKT sg13g2f_FILL4 vdd vss
*.PININFO vdd:B vss:B 
.ENDS

** Created by: circuit_gen.FILL8
** Cell name: FILL8
** Lib name: sg13g2f
.SUBCKT sg13g2f_FILL8 vdd vss
*.PININFO vdd:B vss:B 
.ENDS

** Created by: circuit_gen.INVD0
** Cell name: INVD0
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD0 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU1_M_u3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.INVD1
** Cell name: INVD1
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD1 i z vss vdd
*.PININFO i:I z:O vss:B vdd:B
M0 z i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M1 z i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.INVD2
** Cell name: INVD2
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD2 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.INVD4
** Cell name: INVD4
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD4 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u2_2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u2_3 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_M_u3_2 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_M_u3_3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.INVD6
** Cell name: INVD6
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD6 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MU1_M_u2_2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MU1_M_u2_3 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MU1_M_u2_4 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU1_M_u2_5 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MU1_M_u3_2 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MU1_M_u3_3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MU1_M_u3_4 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MU1_M_u3_5 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
.ENDS

** Created by: circuit_gen.INVD8
** Cell name: INVD8
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD8 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MU1_M_u2_2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MU1_M_u2_3 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MU1_M_u2_4 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU1_M_u2_5 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU1_M_u2_6 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MU1_M_u2_7 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MU1_M_u3_2 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MU1_M_u3_3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MU1_M_u3_4 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MU1_M_u3_5 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MU1_M_u3_6 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MU1_M_u3_7 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
.ENDS

** Created by: circuit_gen.INVD12
** Cell name: INVD12
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD12 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MU1_M_u2_2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MU1_M_u2_3 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MU1_M_u2_4 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU1_M_u2_5 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU1_M_u2_6 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MU1_M_u2_7 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MU1_M_u2_8 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=0
MU1_M_u2_9 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MU1_M_u2_10 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MU1_M_u2_11 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=1
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MU1_M_u3_2 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MU1_M_u3_3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MU1_M_u3_4 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MU1_M_u3_5 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MU1_M_u3_6 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MU1_M_u3_7 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MU1_M_u3_8 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
MU1_M_u3_9 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
MU1_M_u3_10 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
MU1_M_u3_11 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
.ENDS

** Created by: circuit_gen.INVD16
** Cell name: INVD16
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD16 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MU1_M_u2_2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MU1_M_u2_3 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MU1_M_u2_4 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU1_M_u2_5 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU1_M_u2_6 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MU1_M_u2_7 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MU1_M_u2_8 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=0
MU1_M_u2_9 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MU1_M_u2_10 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MU1_M_u2_11 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=1
MU1_M_u2_12 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=12 $flip=0
MU1_M_u2_13 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=13 $flip=1
MU1_M_u2_14 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=14 $flip=0
MU1_M_u2_15 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=15 $flip=1
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MU1_M_u3_2 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MU1_M_u3_3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MU1_M_u3_4 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MU1_M_u3_5 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MU1_M_u3_6 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MU1_M_u3_7 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MU1_M_u3_8 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
MU1_M_u3_9 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
MU1_M_u3_10 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
MU1_M_u3_11 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
MU1_M_u3_12 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=0
MU1_M_u3_13 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=13 $flip=1
MU1_M_u3_14 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=14 $flip=0
MU1_M_u3_15 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=15 $flip=1
.ENDS

** Created by: circuit_gen.MUX2D0
** Cell name: MUX2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_MUX2D0 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI16_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI17_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI16_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI17_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.MUX2D1
** Cell name: MUX2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_MUX2D1 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.200e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=8.400e-07
.ENDS

** Created by: circuit_gen.MUX2D2
** Cell name: MUX2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_MUX2D2 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.200e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU29_0_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU29_1_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU29_0_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU29_1_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.MUX2D4
** Cell name: MUX2D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_MUX2D4 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI21_M_u3 net24 s net28 vss sg13_lv_nmos l=1.300e-07 w=6.200e-07
MU7_M_u3 net16 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=5.350e-07
MI20_0_M_u2 net24 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI20_1_M_u2 net24 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI19_0_M_u2 net16 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.200e-07
MI19_1_M_u2 net16 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.200e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU29_0_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU29_1_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU29_2_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU29_3_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI21_M_u2 net24 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU7_M_u2 net16 s net28 vdd sg13_lv_pmos l=1.300e-07 w=1.095e-06
MI20_0_M_u3 net24 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI20_1_M_u3 net24 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI19_0_M_u3 net16 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI19_1_M_u3 net16 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU29_0_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU29_1_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU29_2_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU29_3_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ND2D0
** Cell name: ND2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND2D0 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI0_M_u3 zn a1 xi0_net6 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI0_M_u4 xi0_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI0_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI0_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.ND2D1
** Cell name: ND2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u3 zn a1 xi1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u4 xi1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ND2D2
** Cell name: ND2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND2D2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MU3_0_M_u3 zn a1 xu3_0_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU3_0_M_u4 xu3_0_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU3_1_M_u4 xu3_1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU3_1_M_u3 zn a1 xu3_1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU3_0_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU3_0_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU3_1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU3_1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ND2D4
** Cell name: ND2D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND2D4 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_0_M_u3 zn a1 xi1_0_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_0_M_u4 xi1_0_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_1_M_u4 xi1_1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_1_M_u3 zn a1 xi1_1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_2_M_u4 xi1_2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_2_M_u3 zn a1 xi1_2_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_3_M_u4 xi1_3_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_3_M_u3 zn a1 xi1_3_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_0_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_0_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_2_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_2_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_3_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_3_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ND3D0
** Cell name: ND3D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND3D0 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI2_M_u4 zn a1 xi2_net10 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u5 xi2_net10 a2 xi2_net13 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u6 xi2_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI2_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI2_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.ND3D1
** Cell name: ND3D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND3D1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 xi1_net10 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u5 xi1_net10 a2 xi1_net13 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u6 xi1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ND3D2
** Cell name: ND3D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND3D2 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI0_0_M_u4 zn a1 xi0_0_net10 vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_0_M_u5 xi0_0_net10 a2 xi0_0_net13 vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_0_M_u6 xi0_0_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_1_M_u4 zn a1 xi0_1_net10 vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_1_M_u5 xi0_1_net10 a2 xi0_1_net13 vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_1_M_u6 xi0_1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_0_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0_0_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0_0_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0_1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0_1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0_1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.NR2D0
** Cell name: NR2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR2D0 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.NR2D1
** Cell name: NR2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.NR2D2
** Cell name: NR2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR2D2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_0_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=1
MI1_0_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=0
MI1_1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
MI1_1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=0
MI1_0_M_u1 xi1_0_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=1
MI1_0_M_u2 zn a1 xi1_0_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MI1_1_M_u2 zn a1 xi1_1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MI1_1_M_u1 xi1_1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
.ENDS

** Created by: circuit_gen.NR2D4
** Cell name: NR2D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR2D4 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI6_0 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=1
MI15_0 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=0
MI15_1 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
MI6_2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=0
MI6_3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=1
MI15_2 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=0
MI15_3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=1
MI6_1 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=0
MI27_0 net26_0_ a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=1
MI28_0 zn a1 net26_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MI28_1 zn a1 net26_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MI27_1 net26_1_ a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
MI27_2 net26_2_ a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=1
MI28_2 zn a1 net26_2_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MI28_3 zn a1 net26_3_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MI27_3 net26_3_ a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=0
.ENDS

** Created by: circuit_gen.NR3D0
** Cell name: NR3D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR3D0 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI0 net28 a2 net25 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u1 net25 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1 zn a1 net28 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.NR3D1
** Cell name: NR3D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR3D1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=1
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=0
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
M_u1_0 net34_0_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=1
MI4_0 net37_0_ a2 net34_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MI5_0 zn a1 net37_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=1
MI5_1 zn a1 net37_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
MI4_1 net37_1_ a2 net34_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
M_u1_1 net34_1_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=0
.ENDS

** Created by: circuit_gen.NR3D2
** Cell name: NR3D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR3D2 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4_0 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
M_u4_1 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=0
MI6_0 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=1
MI6_1 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=0
MI7_0 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MI7_1 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
M_u1_0 net34 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
M_u1_1 net34 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
M_u1_2 net34 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
M_u1_3 net34 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MI22_0 net31 a2 net34 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=1
MI22_1 net31 a2 net34 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=0
MI22_2 net31 a2 net34 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=1
MI22_3 net31 a2 net34 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=0
MI23_0 zn a1 net31 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
MI23_1 zn a1 net31 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
MI23_2 zn a1 net31 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
MI23_3 zn a1 net31 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=0
.ENDS

** Created by: circuit_gen.NR3D4
** Cell name: NR3D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR3D4 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI0_M_u4_0 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=1
MI0_M_u4_1 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=0
MI0_M_u4_2 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=1
MI0_M_u4_3 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=0
MI0_M_u5_0 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=12 $flip=1
MI0_M_u5_1 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=13 $flip=0
MI0_M_u5_2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=14 $flip=1
MI0_M_u5_3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=15 $flip=0
MI0_M_u6_0 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=17 $flip=1
MI0_M_u6_1 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=18 $flip=0
MI0_M_u6_2 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=19 $flip=1
MI0_M_u6_3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=20 $flip=0
MI0_M_u1_0 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MI0_M_u1_1 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MI0_M_u1_2 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MI0_M_u1_3 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MI0_M_u1_4 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MI0_M_u1_5 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MI0_M_u1_6 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MI0_M_u1_7 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MI0_M_u2_0 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=1
MI0_M_u2_1 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=0
MI0_M_u2_2 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=1
MI0_M_u2_3 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=0
MI0_M_u2_4 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=1
MI0_M_u2_5 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=13 $flip=0
MI0_M_u2_6 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=14 $flip=1
MI0_M_u2_7 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=15 $flip=0
MI0_M_u3_0 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=17 $flip=1
MI0_M_u3_1 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=18 $flip=0
MI0_M_u3_2 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=19 $flip=1
MI0_M_u3_3 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=20 $flip=0
MI0_M_u3_4 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=21 $flip=1
MI0_M_u3_5 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=22 $flip=0
MI0_M_u3_6 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=23 $flip=1
MI0_M_u3_7 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=24 $flip=0
.ENDS

** Created by: circuit_gen.OA21D1
** Cell name: OA21D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_OA21D1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OA21D2
** Cell name: OA21D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_OA21D2 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_0_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_1_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_0_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_1_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OAI21D0
** Cell name: OAI21D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_OAI21D0 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.OAI21D1
** Cell name: OAI21D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_OAI21D1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OAI211D0
** Cell name: OAI211D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_OAI211D0 a1 a2 b c vdd vss zn
*.PININFO a1:I a2:I b:I c:I zn:O vdd:B vss:B 
MI8 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI9 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u2 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI7 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI6 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI5 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI4 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u12 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.OAI211D1
** Cell name: OAI211D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_OAI211D1 a1 a2 b c vdd vss zn
*.PININFO a1:I a2:I b:I c:I zn:O vdd:B vss:B 
MI2 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI3 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u11 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u12 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OAI211D4
** Cell name: OAI211D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_OAI211D4 a1 a2 b c vdd vss zn
*.PININFO a1:I a2:I b:I c:I zn:O vdd:B vss:B 
MI13_0 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MI13_1 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MI13_2 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MI13_3 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MI14_0 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MI14_1 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MI14_2 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MI14_3 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MI2_0 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MI2_1 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MI2_2 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=1
MI2_3 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=12 $flip=0
MI12_0 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=13 $flip=0
MI12_1 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=14 $flip=1
MI12_2 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=15 $flip=0
MI12_3 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=16 $flip=1
MI11_0 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=1
MI11_1 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=0
MI11_2 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=1
MI11_3 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
MI9_0 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MI9_1 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MI9_2 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MI9_3 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
M_u12_0 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
M_u12_1 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
M_u12_2 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
M_u12_3 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=0
MI8_0 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=13 $flip=1
MI8_1 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=14 $flip=0
MI8_2 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=15 $flip=1
MI8_3 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=16 $flip=0
.ENDS

** Created by: circuit_gen.OR2D0
** Cell name: OR2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_OR2D0 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.OR2D1
** Cell name: OR2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_OR2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=6.550e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=6.550e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.550e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OR2D2
** Cell name: OR2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_OR2D2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_0_M_u2 z net9 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_1_M_u2 z net9 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u7_M_u4 net9 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u3 net9 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u2 net9 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_0_M_u3 z net9 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_1_M_u3 z net9 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OR2D4
** Cell name: OR2D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_OR2D4 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_0_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_1_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_2_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_3_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u7_0_M_u4 p0 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_0_M_u3 p0 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_1_M_u4 p0 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_1_M_u3 p0 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_0_M_u2 p0 a1 x_u7_0_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_0_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_1_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_2_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_3_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u7_0_M_u1 x_u7_0_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u7_1_M_u1 x_u7_1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u7_1_M_u2 p0 a1 x_u7_1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.TAPCELL
** Cell name: TAPCELL
** Lib name: sg13g2f
.SUBCKT sg13g2f_TAPCELL vdd vss
*.PININFO vdd:B vss:B 
.ENDS

** Created by: circuit_gen.TIEH
** Cell name: TIEH
** Lib name: sg13g2f
.SUBCKT sg13g2f_TIEH vdd vss z
*.PININFO z:O vdd:B vss:B 
M_u2 net6 net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u1 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.TIEL
** Cell name: TIEL
** Lib name: sg13g2f
.SUBCKT sg13g2f_TIEL vdd vss zn
*.PININFO zn:O vdd:B vss:B 
M_u2 zn net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u1 net6 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.XNR2D0
** Cell name: XNR2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_XNR2D0 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI2_M_u3 net28 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI0_M_u3 net6 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI1_M_u2 net28 net6 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
M_u2_M_u2 net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI2_M_u2 net28 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
MI0_M_u2 net6 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
MI1_M_u3 net28 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
M_u2_M_u3 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
.ENDS

** Created by: circuit_gen.XNR2D1
** Cell name: XNR2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_XNR2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.XNR2D2
** Cell name: XNR2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_XNR2D2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u4_0_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u4_1_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u4_0_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u4_1_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.XOR2D0
** Cell name: XOR2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_XOR2D0 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI5_M_u3 net25 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
M_u6_M_u3 net4 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI6_M_u2 net25 net4 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI1_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u4_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI5_M_u2 net25 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
M_u6_M_u2 net4 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
MI6_M_u3 net25 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
MI1_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u4_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI2_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
.ENDS

** Created by: circuit_gen.XOR2D1
** Cell name: XOR2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_XOR2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI4_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI4_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.XOR2D2
** Cell name: XOR2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_XOR2D2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI4_0_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI4_1_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI4_0_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI4_1_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS
** Cell name: SARADC_CELL_INVX0_ASSW
** Lib name: sg13g2f
.SUBCKT SARADC_CELL_INVX0_ASSW i vdd vss zn vnw vpw
*.PININFO i:B zn:B vdd:B vss:B 
MU1_M_u2 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU1_M_u3 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS
** Cell name: SARADC_CELL_INVX16_ASCAP
** Lib name: sg13g2f
.SUBCKT SARADC_CELL_INVX16_ASCAP i vdd vss zn vnw vpw
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MU1_M_u2_1 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MU1_M_u2_2 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MU1_M_u2_3 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MU1_M_u2_4 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU1_M_u2_5 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU1_M_u2_6 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MU1_M_u2_7 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MU1_M_u2_8 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=0
MU1_M_u2_9 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MU1_M_u2_10 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MU1_M_u2_11 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=1
MU1_M_u3_0 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MU1_M_u3_1 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MU1_M_u3_2 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MU1_M_u3_3 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MU1_M_u3_4 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MU1_M_u3_5 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MU1_M_u3_6 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MU1_M_u3_7 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MU1_M_u3_8 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
MU1_M_u3_9 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
MU1_M_u3_10 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
MU1_M_u3_11 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
.ENDS
** Cell name: SARADC_FILLTIE2
** Lib name: sg13g2f
.SUBCKT SARADC_FILLTIE2 vdd vss
*.PININFO vdd:B vss:B 
.ENDS
** Cell name: SARADC_FILL1
.SUBCKT SARADC_FILL1 vdd vss
*.PININFO vdd:B vss:B 
.ENDS
** Cell name: SARADC_FILL1_NOPOWER
.SUBCKT SARADC_FILL1_NOPOWER
.ENDS
* CDL Netlist generated by OpenROAD

*.BUSDELIMITER [

.SUBCKT SARADC AVDD CLK GO RESULT[0] RESULT[1] RESULT[2] RESULT[3]
+ RESULT[4] RST SAMPLE VALID VDD VIN VIP VREFH VREFL VSS
Xanalog/buflogic.conv.cmpbegin.ccmpbuf1.impl analog/buflogic.conv.cmpbegin.CCMPNR
+ AVDD VSS analog/buflogic.conv.cmpbegin.CCMPNR1 sg13g2f_BUFFD8
Xanalog/buflogic.conv.cmpbegin.ccmpbuf2.impl analog/buflogic.conv.cmpbegin.CCMPNR1
+ AVDD VSS analog/buflogic.CMP sg13g2f_BUFFD16
Xanalog/buflogic.conv.cmpbegin.ccmpnor.impl SAMPLE CLKBUF
+ VALID AVDD VSS analog/buflogic.conv.cmpbegin.CCMPNR sg13g2f_NR3D4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.ibuf16.impl RESULTN\[1\]
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.ln1.impl analog/buflogic.conv.re2cr\[1\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.ln2.impl analog/buflogic.conv.re2cr\[1\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zbuf.impl analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD3
+ AVDD VSS analog/CRH\[0\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_1.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_1.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_2.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_2.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_3.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_3.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.znbuf.impl analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD3
+ AVDD VSS analog/CRHB\[0\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_1.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_1.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_2.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_2.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_3.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_3.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.ibuf16.impl RESULT[1]
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.ln1.impl analog/buflogic.conv.re2cr\[1\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.ln2.impl analog/buflogic.conv.re2cr\[1\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zbuf.impl analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD3
+ AVDD VSS analog/CRL\[0\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_1.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_1.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_2.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_2.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_3.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_3.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.znbuf.impl analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD3
+ AVDD VSS analog/CRLB\[0\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_1.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_1.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_2.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_2.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_3.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_3.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.ibuf16.impl RESULTN\[2\]
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.ln1.impl analog/buflogic.conv.re2cr\[2\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.ln2.impl analog/buflogic.conv.re2cr\[2\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zbuf.impl analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD3
+ AVDD VSS analog/CRH\[1\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_1.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_1.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_2.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_2.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_3.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_3.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.znbuf.impl analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD3
+ AVDD VSS analog/CRHB\[1\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_1.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_1.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_2.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_2.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_3.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_3.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.ibuf16.impl RESULT[2]
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.ln1.impl analog/buflogic.conv.re2cr\[2\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.ln2.impl analog/buflogic.conv.re2cr\[2\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zbuf.impl analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD3
+ AVDD VSS analog/CRL\[1\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_1.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_1.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_2.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_2.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_3.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_3.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.znbuf.impl analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD3
+ AVDD VSS analog/CRLB\[1\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_1.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_1.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_2.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_2.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_3.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_3.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.ibuf16.impl RESULTN\[3\]
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.ln1.impl analog/buflogic.conv.re2cr\[3\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.ln2.impl analog/buflogic.conv.re2cr\[3\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zbuf.impl analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD3
+ AVDD VSS analog/CRH\[2\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_1.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_1.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_2.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_2.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_3.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_3.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.znbuf.impl analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD3
+ AVDD VSS analog/CRHB\[2\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_1.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_1.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_2.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_2.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_3.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_3.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.ibuf16.impl RESULT[3]
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.ln1.impl analog/buflogic.conv.re2cr\[3\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.ln2.impl analog/buflogic.conv.re2cr\[3\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zbuf.impl analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD3
+ AVDD VSS analog/CRL\[2\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_1.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_1.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_2.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_2.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_3.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_3.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.znbuf.impl analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD3
+ AVDD VSS analog/CRLB\[2\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_1.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_1.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_2.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_2.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_3.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_3.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.ibuf16.impl RESULTN\[4\]
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.ln1.impl analog/buflogic.conv.re2cr\[4\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.ln2.impl analog/buflogic.conv.re2cr\[4\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zbuf.impl analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD3
+ AVDD VSS analog/CRH\[3\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_1.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_1.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_2.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_2.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_3.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_3.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.znbuf.impl analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD3
+ AVDD VSS analog/CRHB\[3\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_1.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_1.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_2.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_2.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_3.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_3.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.ibuf16.impl RESULT[4]
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.ln1.impl analog/buflogic.conv.re2cr\[4\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.ln2.impl analog/buflogic.conv.re2cr\[4\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zbuf.impl analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD3
+ AVDD VSS analog/CRL\[3\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_1.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_1.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_2.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_2.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_3.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_3.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.znbuf.impl analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD3
+ AVDD VSS analog/CRLB\[3\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_1.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_1.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_2.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_2.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_3.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_3.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.smpcs.choldb.impl analog/buflogic.HOLD
+ AVDD VSS analog/buflogic.conv.smpcs.CHOLDB sg13g2f_INVD8
Xanalog/buflogic.conv.smpcs.choldb1.impl analog/buflogic.conv.smpcs.CHOLDB
+ AVDD VSS analog/buflogic.conv.smpcs.CHOLDB1 sg13g2f_BUFFD8
Xanalog/buflogic.conv.smpcs.clkbuf.impl clknet_1_0__leaf_CLK_regs
+ AVDD VSS CLKBUF sg13g2f_BUFFD16
Xanalog/buflogic.conv.smpcs.clkbufd1.impl1 CLKBUF AVDD VSS
+ analog/buflogic.conv.smpcs.clkbufd1.Z1 sg13g2f_DEL4
Xanalog/buflogic.conv.smpcs.clkbufd1.impl2 analog/buflogic.conv.smpcs.clkbufd1.Z1
+ AVDD VSS analog/buflogic.conv.smpcs.CLKBUFD1 sg13g2f_BUFFD4
Xanalog/buflogic.conv.smpcs.clkbufd2.impl1 analog/buflogic.conv.smpcs.CLKBUFD1
+ AVDD VSS analog/buflogic.conv.smpcs.clkbufd2.Z1 sg13g2f_DEL4
Xanalog/buflogic.conv.smpcs.clkbufd2.impl2 analog/buflogic.conv.smpcs.clkbufd2.Z1
+ AVDD VSS analog/buflogic.conv.smpcs.CLKBUFD2 sg13g2f_BUFFD4
Xanalog/buflogic.conv.smpcs.clkbufd3.impl1 analog/buflogic.conv.smpcs.CLKBUFD2
+ AVDD VSS analog/buflogic.conv.smpcs.clkbufd3.Z1 sg13g2f_DEL4
Xanalog/buflogic.conv.smpcs.clkbufd3.impl2 analog/buflogic.conv.smpcs.clkbufd3.Z1
+ AVDD VSS analog/buflogic.conv.smpcs.CLKBUFD3 sg13g2f_BUFFD4
Xanalog/buflogic.conv.smpcs.cpreand.impl analog/buflogic.conv.smpcs.CHOLDB1
+ analog/buflogic.conv.smpcs.CLKBUFD3 AVDD VSS analog/buflogic.PRE
+ sg13g2f_AN2D4
Xanalog/buflogic.conv.smpcs.invsmp.impl SAMPLE AVDD VSS analog/buflogic.HOLD
+ sg13g2f_INVD8
Xanalog/buflogic.lnbuf_ccmp.del4.impl1 analog/buflogic.CMP
+ AVDD VSS analog/buflogic.lnbuf_ccmp.del4.Z1 sg13g2f_DEL4
Xanalog/buflogic.lnbuf_ccmp.del4.impl2 analog/buflogic.lnbuf_ccmp.del4.Z1
+ AVDD VSS analog/buflogic.lnbuf_ccmp.ID sg13g2f_BUFFD4
Xanalog/buflogic.lnbuf_ccmp.deland.impl analog/buflogic.CMP
+ analog/buflogic.lnbuf_ccmp.ID AVDD VSS analog/buflogic.lnbuf_ccmp.IP
+ sg13g2f_AN2D4
Xanalog/buflogic.lnbuf_ccmp.delbuf16.impl analog/buflogic.lnbuf_ccmp.IP
+ AVDD VSS analog/CCMP sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_ccmp.ln1.impl analog/buflogic.CMP AVDD
+ VSS analog/buflogic.lnbuf_ccmp.IL sg13g2f_INVD6
Xanalog/buflogic.lnbuf_ccmp.ln2.impl analog/buflogic.lnbuf_ccmp.IL
+ AVDD VSS analog/buflogic.CMP sg13g2f_INVD6
Xanalog/buflogic.lnbuf_ccmp.lnbbuf16.impl analog/buflogic.lnbuf_ccmp.ILBUF
+ AVDD VSS analog/CCMPB sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_ccmp.lnbbuf4.impl analog/buflogic.lnbuf_ccmp.IL
+ AVDD VSS analog/buflogic.lnbuf_ccmp.ILBUF sg13g2f_BUFFD4
Xanalog/buflogic.lnbuf_chold.ibuf16.impl analog/buflogic.HOLD
+ AVDD VSS analog/buflogic.lnbuf_chold.N3 sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_chold.ln1.impl analog/buflogic.lnbuf_chold.N3
+ AVDD VSS analog/buflogic.lnbuf_chold.N2 sg13g2f_INVD8
Xanalog/buflogic.lnbuf_chold.ln2.impl analog/buflogic.lnbuf_chold.N2
+ AVDD VSS analog/buflogic.lnbuf_chold.N3 sg13g2f_INVD8
Xanalog/buflogic.lnbuf_chold.zbuf16_1.impl analog/buflogic.lnbuf_chold.N1
+ AVDD VSS analog/CHOLD sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_chold.zbuf16_2.impl analog/buflogic.lnbuf_chold.N1
+ AVDD VSS analog/CHOLD sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_chold.zbuf8.impl analog/buflogic.lnbuf_chold.N3
+ AVDD VSS analog/buflogic.lnbuf_chold.N1 sg13g2f_BUFFD8
Xanalog/buflogic.lnbuf_chold.znbuf16_1.impl analog/buflogic.lnbuf_chold.N2
+ AVDD VSS analog/CHOLDB sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_chold.znbuf16_2.impl analog/buflogic.lnbuf_chold.N2
+ AVDD VSS analog/CHOLDB sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_cpre.ibuf16.impl analog/buflogic.PRE
+ AVDD VSS analog/buflogic.lnbuf_cpre.N3 sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_cpre.ln1.impl analog/buflogic.lnbuf_cpre.N3
+ AVDD VSS analog/buflogic.lnbuf_cpre.N2 sg13g2f_INVD8
Xanalog/buflogic.lnbuf_cpre.ln2.impl analog/buflogic.lnbuf_cpre.N2
+ AVDD VSS analog/buflogic.lnbuf_cpre.N3 sg13g2f_INVD8
Xanalog/buflogic.lnbuf_cpre.zbuf16_1.impl analog/buflogic.lnbuf_cpre.N1
+ AVDD VSS analog/CPRE sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_cpre.zbuf16_2.impl analog/buflogic.lnbuf_cpre.N1
+ AVDD VSS analog/CPRE sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_cpre.zbuf8.impl analog/buflogic.lnbuf_cpre.N3
+ AVDD VSS analog/buflogic.lnbuf_cpre.N1 sg13g2f_BUFFD8
Xanalog/buflogic.lnbuf_cpre.znbuf16_1.impl analog/buflogic.lnbuf_cpre.N2
+ AVDD VSS analog/CPREB sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_cpre.znbuf16_2.impl analog/buflogic.lnbuf_cpre.N2
+ AVDD VSS analog/CPREB sg13g2f_BUFFD16
Xanalog/cmp.buf_n0.impl analog/cmp.OUTNp AVDD VSS analog/cmp.OUTNpb
+ sg13g2f_BUFFD0
Xanalog/cmp.buf_n1.impl analog/cmp.OUTNpb AVDD VSS analog/cmp.OUTN
+ sg13g2f_BUFFD2
Xanalog/cmp.buf_p0.impl analog/cmp.OUTPp AVDD VSS analog/cmp.OUTPpb
+ sg13g2f_BUFFD0
Xanalog/cmp.buf_p1.impl analog/cmp.OUTPpb AVDD VSS CMPO sg13g2f_BUFFD2
Xanalog/cmp.n2p.impl analog/cmp.OUTNp analog/CCMP AVDD VSS
+ analog/cmp.OUTPp sg13g2f_ND2D2
Xanalog/cmp.p2n.impl analog/cmp.OUTPp analog/CCMP AVDD VSS
+ analog/cmp.OUTNp sg13g2f_ND2D2
Xanalog/cmp.vn_cmp.impl_0 analog/CCMPB analog/VOUTL analog/CCMP
+ analog/cmp.OUTNp AVDD VSS analog/cmp.OUTPp sg13g2f_OAI211D4
Xanalog/cmp.vn_cmp.impl_1 analog/CCMPB analog/VOUTL analog/CCMP
+ analog/cmp.OUTNp AVDD VSS analog/cmp.OUTPp sg13g2f_OAI211D4
Xanalog/cmp.vn_cmp.impl_2 analog/CCMPB analog/VOUTL analog/CCMP
+ analog/cmp.OUTNp AVDD VSS analog/cmp.OUTPp sg13g2f_OAI211D4
Xanalog/cmp.vn_cmp.impl_3 analog/CCMPB analog/VOUTL analog/CCMP
+ analog/cmp.OUTNp AVDD VSS analog/cmp.OUTPp sg13g2f_OAI211D4
Xanalog/cmp.vp_cmp.impl_0 analog/CCMPB analog/VOUTH analog/CCMP
+ analog/cmp.OUTPp AVDD VSS analog/cmp.OUTNp sg13g2f_OAI211D4
Xanalog/cmp.vp_cmp.impl_1 analog/CCMPB analog/VOUTH analog/CCMP
+ analog/cmp.OUTPp AVDD VSS analog/cmp.OUTNp sg13g2f_OAI211D4
Xanalog/cmp.vp_cmp.impl_2 analog/CCMPB analog/VOUTH analog/CCMP
+ analog/cmp.OUTPp AVDD VSS analog/cmp.OUTNp sg13g2f_OAI211D4
Xanalog/cmp.vp_cmp.impl_3 analog/CCMPB analog/VOUTH analog/CCMP
+ analog/cmp.OUTPp AVDD VSS analog/cmp.OUTNp sg13g2f_OAI211D4
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VOUTH analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VOUTH
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VOUTH
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VOUTH analog/dummy_h.dummy\[0\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VOUTL analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VOUTL
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VOUTL
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VOUTL analog/dummy_h.dummy\[0\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VREF
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VREF analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VREF analog/dummy_h.dummy\[0\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VREF
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VOUTH analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VOUTH
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VOUTH
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VOUTH analog/dummy_h.dummy\[10\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VOUTL analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VOUTL
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VOUTL
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VOUTL analog/dummy_h.dummy\[10\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VREF
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VREF analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VREF analog/dummy_h.dummy\[10\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VREF
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VOUTH analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VOUTH
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VOUTH
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VOUTH analog/dummy_h.dummy\[11\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VOUTL analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VOUTL
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VOUTL
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VOUTL analog/dummy_h.dummy\[11\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VREF
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VREF analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VREF analog/dummy_h.dummy\[11\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VREF
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VOUTH analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VOUTH
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VOUTH
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VOUTH analog/dummy_h.dummy\[12\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VOUTL analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VOUTL
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VOUTL
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VOUTL analog/dummy_h.dummy\[12\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VREF
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VREF analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VREF analog/dummy_h.dummy\[12\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VREF
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VOUTH analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VOUTH
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VOUTH
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VOUTH analog/dummy_h.dummy\[13\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VOUTL analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VOUTL
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VOUTL
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VOUTL analog/dummy_h.dummy\[13\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VREF
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VREF analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VREF analog/dummy_h.dummy\[13\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VREF
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VOUTH analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VOUTH
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VOUTH
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VOUTH analog/dummy_h.dummy\[14\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VOUTL analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VOUTL
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VOUTL
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VOUTL analog/dummy_h.dummy\[14\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VREF
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VREF analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VREF analog/dummy_h.dummy\[14\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VREF
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VOUTH analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VOUTH
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VOUTH
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VOUTH analog/dummy_h.dummy\[15\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VOUTL analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VOUTL
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VOUTL
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VOUTL analog/dummy_h.dummy\[15\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VREF
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VREF analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VREF analog/dummy_h.dummy\[15\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VREF
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VOUTH analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VOUTH
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VOUTH
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VOUTH analog/dummy_h.dummy\[16\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VOUTL analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VOUTL
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VOUTL
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VOUTL analog/dummy_h.dummy\[16\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VREF
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VREF analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VREF analog/dummy_h.dummy\[16\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VREF
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VOUTH analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VOUTH
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VOUTH
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VOUTH analog/dummy_h.dummy\[17\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VOUTL analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VOUTL
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VOUTL
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VOUTL analog/dummy_h.dummy\[17\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VREF
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VREF analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VREF analog/dummy_h.dummy\[17\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VREF
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VOUTH analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VOUTH
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VOUTH
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VOUTH analog/dummy_h.dummy\[18\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VOUTL analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VOUTL
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VOUTL
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VOUTL analog/dummy_h.dummy\[18\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VREF
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VREF analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VREF analog/dummy_h.dummy\[18\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VREF
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VOUTH analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VOUTH
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VOUTH
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VOUTH analog/dummy_h.dummy\[19\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VOUTL analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VOUTL
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VOUTL
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VOUTL analog/dummy_h.dummy\[19\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VREF
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VREF analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VREF analog/dummy_h.dummy\[19\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VREF
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VOUTH analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VOUTH
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VOUTH
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VOUTH analog/dummy_h.dummy\[1\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VOUTL analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VOUTL
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VOUTL
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VOUTL analog/dummy_h.dummy\[1\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VREF
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VREF analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VREF analog/dummy_h.dummy\[1\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VREF
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VOUTH analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VOUTH
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VOUTH
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VOUTH analog/dummy_h.dummy\[20\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VOUTL analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VOUTL
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VOUTL
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VOUTL analog/dummy_h.dummy\[20\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VREF
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VREF analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VREF analog/dummy_h.dummy\[20\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VREF
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VOUTH analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VOUTH
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VOUTH
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VOUTH analog/dummy_h.dummy\[21\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VOUTL analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VOUTL
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VOUTL
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VOUTL analog/dummy_h.dummy\[21\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VREF
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VREF analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VREF analog/dummy_h.dummy\[21\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VREF
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VOUTH analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VOUTH
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VOUTH
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VOUTH analog/dummy_h.dummy\[22\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VOUTL analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VOUTL
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VOUTL
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VOUTL analog/dummy_h.dummy\[22\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VREF
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VREF analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VREF analog/dummy_h.dummy\[22\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VREF
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VOUTH analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VOUTH
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VOUTH
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VOUTH analog/dummy_h.dummy\[23\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VOUTL analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VOUTL
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VOUTL
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VOUTL analog/dummy_h.dummy\[23\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VREF
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VREF analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VREF analog/dummy_h.dummy\[23\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VREF
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VOUTH analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VOUTH
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VOUTH
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VOUTH analog/dummy_h.dummy\[24\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VOUTL analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VOUTL
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VOUTL
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VOUTL analog/dummy_h.dummy\[24\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VREF
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VREF analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VREF analog/dummy_h.dummy\[24\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VREF
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VOUTH analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VOUTH
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VOUTH
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VOUTH analog/dummy_h.dummy\[25\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VOUTL analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VOUTL
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VOUTL
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VOUTL analog/dummy_h.dummy\[25\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VREF
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VREF analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VREF analog/dummy_h.dummy\[25\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VREF
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VOUTH analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VOUTH
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VOUTH
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VOUTH analog/dummy_h.dummy\[26\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VOUTL analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VOUTL
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VOUTL
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VOUTL analog/dummy_h.dummy\[26\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VREF
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VREF analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VREF analog/dummy_h.dummy\[26\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VREF
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VOUTH analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VOUTH
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VOUTH
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VOUTH analog/dummy_h.dummy\[27\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VOUTL analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VOUTL
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VOUTL
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VOUTL analog/dummy_h.dummy\[27\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VREF
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VREF analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VREF analog/dummy_h.dummy\[27\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VREF
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VOUTH analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VOUTH
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VOUTH
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VOUTH analog/dummy_h.dummy\[2\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VOUTL analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VOUTL
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VOUTL
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VOUTL analog/dummy_h.dummy\[2\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VREF
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VREF analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VREF analog/dummy_h.dummy\[2\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VREF
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VOUTH analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VOUTH
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VOUTH
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VOUTH analog/dummy_h.dummy\[3\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VOUTL analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VOUTL
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VOUTL
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VOUTL analog/dummy_h.dummy\[3\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VREF
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VREF analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VREF analog/dummy_h.dummy\[3\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VREF
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VOUTH analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VOUTH
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VOUTH
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VOUTH analog/dummy_h.dummy\[4\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VOUTL analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VOUTL
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VOUTL
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VOUTL analog/dummy_h.dummy\[4\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VREF
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VREF analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VREF analog/dummy_h.dummy\[4\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VREF
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VOUTH analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VOUTH
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VOUTH
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VOUTH analog/dummy_h.dummy\[5\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VOUTL analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VOUTL
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VOUTL
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VOUTL analog/dummy_h.dummy\[5\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VREF
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VREF analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VREF analog/dummy_h.dummy\[5\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VREF
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VOUTH analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VOUTH
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VOUTH
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VOUTH analog/dummy_h.dummy\[6\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VOUTL analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VOUTL
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VOUTL
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VOUTL analog/dummy_h.dummy\[6\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VREF
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VREF analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VREF analog/dummy_h.dummy\[6\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VREF
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VOUTH analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VOUTH
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VOUTH
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VOUTH analog/dummy_h.dummy\[7\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VOUTL analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VOUTL
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VOUTL
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VOUTL analog/dummy_h.dummy\[7\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VREF
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VREF analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VREF analog/dummy_h.dummy\[7\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VREF
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VOUTH analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VOUTH
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VOUTH
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VOUTH analog/dummy_h.dummy\[8\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VOUTL analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VOUTL
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VOUTL
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VOUTL analog/dummy_h.dummy\[8\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VREF
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VREF analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VREF analog/dummy_h.dummy\[8\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VREF
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VOUTH analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VOUTH
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VOUTH
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VOUTH analog/dummy_h.dummy\[9\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VOUTL analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VOUTL
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VOUTL
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VOUTL analog/dummy_h.dummy\[9\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VREF
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VREF analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VREF analog/dummy_h.dummy\[9\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VREF
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.tieh.impl AVDD VSS analog/dummy_h.dummy\[0\].dummy.CRHB
+ sg13g2f_TIEH
Xanalog/dummy_h.tiel.impl AVDD VSS analog/dummy_h.dummy\[0\].dummy.CRH
+ sg13g2f_TIEL
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VOUTH analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VOUTH
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VOUTH
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VOUTH analog/dummy_l.dummy\[0\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VOUTL analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VOUTL
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VOUTL
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VOUTL analog/dummy_l.dummy\[0\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VREF
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VREF analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VREF analog/dummy_l.dummy\[0\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VREF
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VOUTH analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VOUTH
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VOUTH
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VOUTH analog/dummy_l.dummy\[10\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VOUTL analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VOUTL
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VOUTL
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VOUTL analog/dummy_l.dummy\[10\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VREF
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VREF analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VREF analog/dummy_l.dummy\[10\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VREF
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VOUTH analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VOUTH
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VOUTH
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VOUTH analog/dummy_l.dummy\[11\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VOUTL analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VOUTL
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VOUTL
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VOUTL analog/dummy_l.dummy\[11\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VREF
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VREF analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VREF analog/dummy_l.dummy\[11\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VREF
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VOUTH analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VOUTH
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VOUTH
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VOUTH analog/dummy_l.dummy\[12\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VOUTL analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VOUTL
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VOUTL
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VOUTL analog/dummy_l.dummy\[12\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VREF
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VREF analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VREF analog/dummy_l.dummy\[12\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VREF
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VOUTH analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VOUTH
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VOUTH
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VOUTH analog/dummy_l.dummy\[13\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VOUTL analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VOUTL
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VOUTL
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VOUTL analog/dummy_l.dummy\[13\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VREF
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VREF analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VREF analog/dummy_l.dummy\[13\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VREF
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VOUTH analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VOUTH
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VOUTH
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VOUTH analog/dummy_l.dummy\[14\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VOUTL analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VOUTL
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VOUTL
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VOUTL analog/dummy_l.dummy\[14\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VREF
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VREF analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VREF analog/dummy_l.dummy\[14\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VREF
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VOUTH analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VOUTH
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VOUTH
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VOUTH analog/dummy_l.dummy\[15\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VOUTL analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VOUTL
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VOUTL
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VOUTL analog/dummy_l.dummy\[15\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VREF
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VREF analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VREF analog/dummy_l.dummy\[15\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VREF
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VOUTH analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VOUTH
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VOUTH
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VOUTH analog/dummy_l.dummy\[16\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VOUTL analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VOUTL
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VOUTL
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VOUTL analog/dummy_l.dummy\[16\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VREF
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VREF analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VREF analog/dummy_l.dummy\[16\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VREF
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VOUTH analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VOUTH
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VOUTH
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VOUTH analog/dummy_l.dummy\[17\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VOUTL analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VOUTL
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VOUTL
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VOUTL analog/dummy_l.dummy\[17\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VREF
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VREF analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VREF analog/dummy_l.dummy\[17\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VREF
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VOUTH analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VOUTH
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VOUTH
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VOUTH analog/dummy_l.dummy\[18\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VOUTL analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VOUTL
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VOUTL
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VOUTL analog/dummy_l.dummy\[18\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VREF
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VREF analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VREF analog/dummy_l.dummy\[18\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VREF
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VOUTH analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VOUTH
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VOUTH
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VOUTH analog/dummy_l.dummy\[19\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VOUTL analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VOUTL
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VOUTL
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VOUTL analog/dummy_l.dummy\[19\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VREF
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VREF analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VREF analog/dummy_l.dummy\[19\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VREF
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VOUTH analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VOUTH
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VOUTH
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VOUTH analog/dummy_l.dummy\[1\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VOUTL analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VOUTL
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VOUTL
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VOUTL analog/dummy_l.dummy\[1\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VREF
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VREF analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VREF analog/dummy_l.dummy\[1\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VREF
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VOUTH analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VOUTH
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VOUTH
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VOUTH analog/dummy_l.dummy\[20\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VOUTL analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VOUTL
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VOUTL
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VOUTL analog/dummy_l.dummy\[20\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VREF
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VREF analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VREF analog/dummy_l.dummy\[20\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VREF
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VOUTH analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VOUTH
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VOUTH
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VOUTH analog/dummy_l.dummy\[21\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VOUTL analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VOUTL
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VOUTL
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VOUTL analog/dummy_l.dummy\[21\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VREF
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VREF analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VREF analog/dummy_l.dummy\[21\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VREF
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VOUTH analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VOUTH
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VOUTH
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VOUTH analog/dummy_l.dummy\[22\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VOUTL analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VOUTL
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VOUTL
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VOUTL analog/dummy_l.dummy\[22\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VREF
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VREF analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VREF analog/dummy_l.dummy\[22\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VREF
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VOUTH analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VOUTH
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VOUTH
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VOUTH analog/dummy_l.dummy\[23\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VOUTL analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VOUTL
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VOUTL
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VOUTL analog/dummy_l.dummy\[23\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VREF
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VREF analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VREF analog/dummy_l.dummy\[23\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VREF
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VOUTH analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VOUTH
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VOUTH
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VOUTH analog/dummy_l.dummy\[24\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VOUTL analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VOUTL
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VOUTL
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VOUTL analog/dummy_l.dummy\[24\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VREF
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VREF analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VREF analog/dummy_l.dummy\[24\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VREF
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VOUTH analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VOUTH
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VOUTH
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VOUTH analog/dummy_l.dummy\[25\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VOUTL analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VOUTL
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VOUTL
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VOUTL analog/dummy_l.dummy\[25\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VREF
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VREF analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VREF analog/dummy_l.dummy\[25\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VREF
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VOUTH analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VOUTH
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VOUTH
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VOUTH analog/dummy_l.dummy\[26\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VOUTL analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VOUTL
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VOUTL
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VOUTL analog/dummy_l.dummy\[26\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VREF
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VREF analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VREF analog/dummy_l.dummy\[26\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VREF
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VOUTH analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VOUTH
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VOUTH
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VOUTH analog/dummy_l.dummy\[27\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VOUTL analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VOUTL
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VOUTL
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VOUTL analog/dummy_l.dummy\[27\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VREF
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VREF analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VREF analog/dummy_l.dummy\[27\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VREF
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VOUTH analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VOUTH
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VOUTH
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VOUTH analog/dummy_l.dummy\[2\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VOUTL analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VOUTL
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VOUTL
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VOUTL analog/dummy_l.dummy\[2\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VREF
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VREF analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VREF analog/dummy_l.dummy\[2\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VREF
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VOUTH analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VOUTH
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VOUTH
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VOUTH analog/dummy_l.dummy\[3\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VOUTL analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VOUTL
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VOUTL
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VOUTL analog/dummy_l.dummy\[3\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VREF
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VREF analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VREF analog/dummy_l.dummy\[3\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VREF
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VOUTH analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VOUTH
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VOUTH
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VOUTH analog/dummy_l.dummy\[4\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VOUTL analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VOUTL
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VOUTL
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VOUTL analog/dummy_l.dummy\[4\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VREF
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VREF analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VREF analog/dummy_l.dummy\[4\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VREF
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VOUTH analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VOUTH
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VOUTH
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VOUTH analog/dummy_l.dummy\[5\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VOUTL analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VOUTL
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VOUTL
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VOUTL analog/dummy_l.dummy\[5\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VREF
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VREF analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VREF analog/dummy_l.dummy\[5\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VREF
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VOUTH analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VOUTH
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VOUTH
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VOUTH analog/dummy_l.dummy\[6\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VOUTL analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VOUTL
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VOUTL
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VOUTL analog/dummy_l.dummy\[6\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VREF
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VREF analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VREF analog/dummy_l.dummy\[6\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VREF
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VOUTH analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VOUTH
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VOUTH
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VOUTH analog/dummy_l.dummy\[7\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VOUTL analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VOUTL
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VOUTL
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VOUTL analog/dummy_l.dummy\[7\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VREF
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VREF analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VREF analog/dummy_l.dummy\[7\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VREF
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VOUTH analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VOUTH
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VOUTH
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VOUTH analog/dummy_l.dummy\[8\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VOUTL analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VOUTL
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VOUTL
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VOUTL analog/dummy_l.dummy\[8\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VREF
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VREF analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VREF analog/dummy_l.dummy\[8\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VREF
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VOUTH analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VOUTH
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VOUTH
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VOUTH analog/dummy_l.dummy\[9\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VOUTL analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VOUTL
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VOUTL
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VOUTL analog/dummy_l.dummy\[9\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VREF
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VREF analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VREF analog/dummy_l.dummy\[9\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VREF
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.tieh.impl AVDD VSS analog/dummy_l.dummy\[0\].dummy.CRHB
+ sg13g2f_TIEH
Xanalog/dummy_l.tiel.impl AVDD VSS analog/dummy_l.dummy\[0\].dummy.CRH
+ sg13g2f_TIEL
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[0\] analog/LSB_H_VSH\[1\] analog/VOUTH analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[0\] analog/VOUTH analog/LSB_H_VSH\[1\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[0\] analog/VOUTH analog/LSB_H_VSH\[1\] analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[0\] analog/LSB_H_VSH\[1\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[0\] analog/LSB_H_VSH\[1\] analog/VOUTL analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[0\] analog/VOUTL analog/LSB_H_VSH\[1\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[0\] analog/VOUTL analog/LSB_H_VSH\[1\] analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[0\] analog/LSB_H_VSH\[1\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[1\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[1\] VREFH analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[1\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[1\] analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[1\] analog/LSB_H_VSH\[2\] analog/VOUTH analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[1\] analog/VOUTH analog/LSB_H_VSH\[2\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[1\] analog/VOUTH analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[1\] analog/LSB_H_VSH\[2\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[1\] analog/LSB_H_VSH\[2\] analog/VOUTH analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[1\] analog/VOUTH analog/LSB_H_VSH\[2\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[1\] analog/VOUTH analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[1\] analog/LSB_H_VSH\[2\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[1\] analog/LSB_H_VSH\[2\] analog/VOUTL analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[1\] analog/VOUTL analog/LSB_H_VSH\[2\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[1\] analog/VOUTL analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[1\] analog/LSB_H_VSH\[2\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[1\] analog/LSB_H_VSH\[2\] analog/VOUTL analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[1\] analog/VOUTL analog/LSB_H_VSH\[2\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[1\] analog/VOUTL analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[1\] analog/LSB_H_VSH\[2\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[2\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[2\] VREFH analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[2\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[2\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[2\] VREFH analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[2\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[12\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[13\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[14\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[15\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[16\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[17\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[18\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[19\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[20\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[21\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[22\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[23\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[3\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[3\] VREFH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[3\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[3\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[3\] VREFH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[3\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[3\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[3\] VREFH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[3\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[3\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[3\] VREFH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[3\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[12\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[13\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[14\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[15\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[16\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[17\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[18\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[19\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[20\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[21\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[22\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[23\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[24\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[25\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[26\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[27\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[28\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[29\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[30\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[31\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[32\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[33\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[34\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[35\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[36\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[37\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[38\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[39\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[40\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[41\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[42\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[43\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[44\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[45\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[46\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[47\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/lsb_cdac_h.cdac_unit.CRH analog/LSB_H_VSH\[0\] analog/VOUTH
+ analog/LSB_H_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/lsb_cdac_h.cdac_unit.CRH analog/VOUTH analog/LSB_H_VSH\[0\]
+ analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/lsb_cdac_h.cdac_unit.CRHB analog/VOUTH analog/LSB_H_VSH\[0\]
+ analog/LSB_H_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/lsb_cdac_h.cdac_unit.CRHB analog/LSB_H_VSH\[0\] analog/VOUTH
+ analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/lsb_cdac_h.cdac_unit.CRH analog/LSB_H_VSH\[0\] analog/VOUTL
+ analog/LSB_H_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/lsb_cdac_h.cdac_unit.CRH analog/VOUTL analog/LSB_H_VSH\[0\]
+ analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/lsb_cdac_h.cdac_unit.CRHB analog/VOUTL analog/LSB_H_VSH\[0\]
+ analog/LSB_H_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/lsb_cdac_h.cdac_unit.CRHB analog/LSB_H_VSH\[0\] analog/VOUTL
+ analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap\[0\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.cap\[1\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.cap\[2\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.cap\[3\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.cap\[4\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.cap\[5\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[0\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[0\] VREFH analog/LSB_H_VSH\[0\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[0\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[0\] analog/LSB_H_VSH\[0\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.tieh.impl AVDD VSS analog/lsb_cdac_h.cdac_unit.CRHB
+ sg13g2f_TIEH
Xanalog/lsb_cdac_h.tiel.impl AVDD VSS analog/lsb_cdac_h.cdac_unit.CRH
+ sg13g2f_TIEL
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[0\] analog/LSB_L_VSH\[1\] analog/VOUTL analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[0\] analog/VOUTL analog/LSB_L_VSH\[1\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[0\] analog/VOUTL analog/LSB_L_VSH\[1\] analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[0\] analog/LSB_L_VSH\[1\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[0\] analog/LSB_L_VSH\[1\] analog/VOUTH analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[0\] analog/VOUTH analog/LSB_L_VSH\[1\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[0\] analog/VOUTH analog/LSB_L_VSH\[1\] analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[0\] analog/LSB_L_VSH\[1\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[1\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[1\] VREFL analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[1\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[1\] analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[1\] analog/LSB_L_VSH\[2\] analog/VOUTL analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[1\] analog/VOUTL analog/LSB_L_VSH\[2\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[1\] analog/VOUTL analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[1\] analog/LSB_L_VSH\[2\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[1\] analog/LSB_L_VSH\[2\] analog/VOUTL analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[1\] analog/VOUTL analog/LSB_L_VSH\[2\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[1\] analog/VOUTL analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[1\] analog/LSB_L_VSH\[2\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[1\] analog/LSB_L_VSH\[2\] analog/VOUTH analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[1\] analog/VOUTH analog/LSB_L_VSH\[2\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[1\] analog/VOUTH analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[1\] analog/LSB_L_VSH\[2\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[1\] analog/LSB_L_VSH\[2\] analog/VOUTH analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[1\] analog/VOUTH analog/LSB_L_VSH\[2\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[1\] analog/VOUTH analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[1\] analog/LSB_L_VSH\[2\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[2\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[2\] VREFL analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[2\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[2\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[2\] VREFL analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[2\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[12\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[13\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[14\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[15\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[16\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[17\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[18\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[19\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[20\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[21\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[22\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[23\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[3\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[3\] VREFL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[3\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[3\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[3\] VREFL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[3\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[3\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[3\] VREFL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[3\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[3\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[3\] VREFL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[3\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[12\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[13\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[14\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[15\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[16\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[17\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[18\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[19\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[20\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[21\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[22\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[23\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[24\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[25\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[26\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[27\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[28\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[29\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[30\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[31\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[32\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[33\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[34\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[35\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[36\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[37\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[38\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[39\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[40\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[41\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[42\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[43\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[44\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[45\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[46\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[47\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/lsb_cdac_l.cdac_unit.CRH analog/LSB_L_VSH\[0\] analog/VOUTL
+ analog/LSB_L_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/lsb_cdac_l.cdac_unit.CRH analog/VOUTL analog/LSB_L_VSH\[0\]
+ analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/lsb_cdac_l.cdac_unit.CRHB analog/VOUTL analog/LSB_L_VSH\[0\]
+ analog/LSB_L_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/lsb_cdac_l.cdac_unit.CRHB analog/LSB_L_VSH\[0\] analog/VOUTL
+ analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/lsb_cdac_l.cdac_unit.CRH analog/LSB_L_VSH\[0\] analog/VOUTH
+ analog/LSB_L_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/lsb_cdac_l.cdac_unit.CRH analog/VOUTH analog/LSB_L_VSH\[0\]
+ analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/lsb_cdac_l.cdac_unit.CRHB analog/VOUTH analog/LSB_L_VSH\[0\]
+ analog/LSB_L_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/lsb_cdac_l.cdac_unit.CRHB analog/LSB_L_VSH\[0\] analog/VOUTH
+ analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap\[0\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.cap\[1\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.cap\[2\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.cap\[3\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.cap\[4\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.cap\[5\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[0\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[0\] VREFL analog/LSB_L_VSH\[0\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[0\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[0\] analog/LSB_L_VSH\[0\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.tieh.impl AVDD VSS analog/lsb_cdac_l.cdac_unit.CRHB
+ sg13g2f_TIEH
Xanalog/lsb_cdac_l.tiel.impl AVDD VSS analog/lsb_cdac_l.cdac_unit.CRH
+ sg13g2f_TIEL
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap\[0\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[10\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[11\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[12\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[13\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[14\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[15\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[16\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[17\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[18\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[19\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[1\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[20\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[21\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[22\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[23\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[24\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[25\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[26\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[27\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[28\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[29\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[2\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[30\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[31\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[32\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[33\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[34\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[35\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[36\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[37\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[38\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[39\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[3\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[40\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[41\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[42\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[43\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[44\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[45\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[46\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[47\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[48\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[49\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[4\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[50\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[51\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[52\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[53\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[54\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[55\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[56\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[57\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[58\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[59\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[5\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[60\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[61\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[62\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[63\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[64\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[65\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[66\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[67\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[68\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[69\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[6\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[70\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[71\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[72\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[73\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[74\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[75\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[76\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[77\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[78\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[79\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[7\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[80\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[81\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[82\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[83\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[84\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[85\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[86\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[87\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[88\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[89\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[8\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[90\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[91\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[92\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[93\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[94\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[95\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[9\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.tieh.impl AVDD VSS analog/msb_cdac_h.cdac_unit.CRLB
+ sg13g2f_TIEH
Xanalog/msb_cdac_h.tiel.impl AVDD VSS analog/msb_cdac_h.cdac_unit.CRL
+ sg13g2f_TIEL
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap\[0\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[10\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[11\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[12\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[13\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[14\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[15\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[16\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[17\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[18\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[19\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[1\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[20\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[21\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[22\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[23\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[24\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[25\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[26\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[27\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[28\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[29\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[2\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[30\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[31\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[32\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[33\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[34\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[35\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[36\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[37\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[38\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[39\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[3\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[40\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[41\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[42\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[43\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[44\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[45\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[46\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[47\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[48\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[49\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[4\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[50\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[51\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[52\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[53\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[54\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[55\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[56\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[57\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[58\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[59\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[5\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[60\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[61\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[62\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[63\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[64\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[65\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[66\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[67\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[68\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[69\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[6\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[70\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[71\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[72\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[73\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[74\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[75\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[76\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[77\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[78\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[79\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[7\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[80\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[81\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[82\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[83\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[84\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[85\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[86\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[87\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[88\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[89\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[8\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[90\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[91\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[92\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[93\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[94\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[95\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[9\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.tieh.impl AVDD VSS analog/msb_cdac_l.cdac_unit.CRLB
+ sg13g2f_TIEH
Xanalog/msb_cdac_l.tiel.impl AVDD VSS analog/msb_cdac_l.cdac_unit.CRL
+ sg13g2f_TIEL
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz1 analog/CPRE
+ analog/VOUTH analog/VOUTL analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2 analog/CPRE
+ analog/VOUTL analog/VOUTH analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz1 analog/CPREB
+ analog/VOUTL analog/VOUTH analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz2 analog/CPREB
+ analog/VOUTH analog/VOUTL analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz1 analog/CPRE
+ analog/VOUTH analog/VOUTL analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2 analog/CPRE
+ analog/VOUTL analog/VOUTH analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz1 analog/CPREB
+ analog/VOUTL analog/VOUTH analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz2 analog/CPREB
+ analog/VOUTH analog/VOUTL analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgn_lz1 analog/CPRE
+ analog/VOUTH analog/VOUTL analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgn_lz2 analog/CPRE
+ analog/VOUTL analog/VOUTH analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz1 analog/CPREB
+ analog/VOUTL analog/VOUTH analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz2 analog/CPREB
+ analog/VOUTH analog/VOUTL analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xdigital/ins_051_ digital/state\[1\] digital/ins_017_ VSS
+ VDD sg13g2f_INVD1
Xdigital/ins_052_ digital/state\[0\] digital/ins_018_ VSS
+ VDD sg13g2f_INVD1
Xdigital/ins_053_ digital/mask\[0\] digital/ins_019_ VSS VDD
+ sg13g2f_INVD1
Xdigital/ins_054_ digital/mask\[1\] digital/ins_020_ VSS VDD
+ sg13g2f_INVD1
Xdigital/ins_055_ digital/mask\[2\] digital/ins_021_ VSS VDD
+ sg13g2f_INVD1
Xdigital/ins_056_ digital/mask\[3\] digital/ins_022_ VSS VDD
+ sg13g2f_INVD1
Xdigital/ins_057_ digital/mask\[4\] digital/ins_023_ VSS VDD
+ sg13g2f_INVD1
Xdigital/ins_058_ RST digital/ins_024_ VSS VDD sg13g2f_INVD1
Xdigital/ins_059_ RESULT[0] digital/ins_025_ VSS VDD sg13g2f_INVD1
Xdigital/ins_060_ RESULT[1] digital/ins_026_ VSS VDD sg13g2f_INVD1
Xdigital/ins_061_ RESULT[2] digital/ins_027_ VSS VDD sg13g2f_INVD1
Xdigital/ins_062_ RESULT[3] digital/ins_028_ VSS VDD sg13g2f_INVD1
Xdigital/ins_063_ RESULT[4] digital/ins_029_ VSS VDD sg13g2f_INVD1
Xdigital/ins_064_ digital/state\[1\] digital/ins_018_ RST
+ VDD VSS digital/ins_030_ sg13g2f_AOI21D1
Xdigital/ins_065_ digital/state\[1\] digital/ins_018_ RST
+ VDD VSS digital/ins_031_ sg13g2f_AO21D1
Xdigital/ins_066_ RST CMPO VDD VSS digital/ins_032_ sg13g2f_NR2D1
Xdigital/ins_067_ digital/mask\[0\] digital/ins_032_ RESULTN\[0\]
+ VDD VSS digital/ins_033_ sg13g2f_AO21D1
Xdigital/ins_068_ digital/ins_031_ digital/ins_033_ VDD VSS
+ digital/ins_000_ sg13g2f_AN2D1
Xdigital/ins_069_ digital/mask\[1\] digital/ins_032_ RESULTN\[1\]
+ VDD VSS digital/ins_034_ sg13g2f_AO21D1
Xdigital/ins_070_ digital/ins_031_ digital/ins_034_ VDD VSS
+ digital/ins_001_ sg13g2f_AN2D1
Xdigital/ins_071_ digital/mask\[2\] digital/ins_032_ RESULTN\[2\]
+ VDD VSS digital/ins_035_ sg13g2f_AO21D1
Xdigital/ins_072_ digital/ins_031_ digital/ins_035_ VDD VSS
+ digital/ins_002_ sg13g2f_AN2D1
Xdigital/ins_073_ digital/mask\[3\] digital/ins_032_ RESULTN\[3\]
+ VDD VSS digital/ins_036_ sg13g2f_AO21D1
Xdigital/ins_074_ digital/ins_031_ digital/ins_036_ VDD VSS
+ digital/ins_003_ sg13g2f_AN2D1
Xdigital/ins_075_ digital/mask\[4\] digital/ins_032_ RESULTN\[4\]
+ VDD VSS digital/ins_037_ sg13g2f_AO21D1
Xdigital/ins_076_ digital/ins_031_ digital/ins_037_ VDD VSS
+ digital/ins_004_ sg13g2f_AN2D1
Xdigital/ins_077_ digital/state\[1\] digital/ins_018_ digital/ins_024_
+ VDD VSS digital/ins_038_ sg13g2f_ND3D1
Xdigital/ins_078_ digital/ins_017_ digital/state\[0\] VDD
+ VSS SAMPLE sg13g2f_AN2D1
Xdigital/ins_079_ digital/ins_017_ digital/state\[0\] digital/ins_024_
+ VDD VSS digital/ins_039_ sg13g2f_ND3D1
Xdigital/ins_080_ digital/state\[1\] digital/state\[0\] VDD
+ VSS digital/ins_040_ sg13g2f_XNR2D1
Xdigital/ins_081_ RST digital/ins_040_ VDD VSS digital/ins_011_
+ sg13g2f_NR2D1
Xdigital/ins_082_ RST digital/ins_040_ digital/mask\[0\] VDD
+ VSS digital/ins_041_ sg13g2f_OAI21D1
Xdigital/ins_083_ digital/ins_020_ digital/ins_038_ digital/ins_041_
+ VDD VSS digital/ins_005_ sg13g2f_OAI21D1
Xdigital/ins_084_ RST digital/ins_040_ digital/mask\[1\] VDD
+ VSS digital/ins_042_ sg13g2f_OAI21D1
Xdigital/ins_085_ digital/ins_021_ digital/ins_038_ digital/ins_042_
+ VDD VSS digital/ins_006_ sg13g2f_OAI21D1
Xdigital/ins_086_ RST digital/ins_040_ digital/mask\[2\] VDD
+ VSS digital/ins_043_ sg13g2f_OAI21D1
Xdigital/ins_087_ digital/ins_022_ digital/ins_038_ digital/ins_043_
+ VDD VSS digital/ins_007_ sg13g2f_OAI21D1
Xdigital/ins_088_ RST digital/ins_040_ digital/mask\[3\] VDD
+ VSS digital/ins_044_ sg13g2f_OAI21D1
Xdigital/ins_089_ digital/ins_023_ digital/ins_038_ digital/ins_044_
+ VDD VSS digital/ins_008_ sg13g2f_OAI21D1
Xdigital/ins_090_ digital/ins_023_ digital/ins_011_ digital/ins_039_
+ VDD VSS digital/ins_009_ sg13g2f_OAI21D1
Xdigital/ins_091_ digital/ins_024_ GO digital/ins_040_ VDD
+ VSS digital/ins_045_ sg13g2f_ND3D1
Xdigital/ins_092_ digital/ins_019_ digital/ins_038_ digital/ins_045_
+ VDD VSS digital/ins_010_ sg13g2f_OAI21D1
Xdigital/ins_093_ digital/mask\[0\] digital/ins_024_ CMPO
+ VDD VSS digital/ins_046_ sg13g2f_ND3D1
Xdigital/ins_094_ digital/ins_025_ digital/ins_046_ digital/ins_030_
+ VDD VSS digital/ins_012_ sg13g2f_AOI21D1
Xdigital/ins_095_ digital/mask\[1\] digital/ins_024_ CMPO
+ VDD VSS digital/ins_047_ sg13g2f_ND3D1
Xdigital/ins_096_ digital/ins_026_ digital/ins_047_ digital/ins_030_
+ VDD VSS digital/ins_013_ sg13g2f_AOI21D1
Xdigital/ins_097_ digital/mask\[2\] digital/ins_024_ CMPO
+ VDD VSS digital/ins_048_ sg13g2f_ND3D1
Xdigital/ins_098_ digital/ins_027_ digital/ins_048_ digital/ins_030_
+ VDD VSS digital/ins_014_ sg13g2f_AOI21D1
Xdigital/ins_099_ digital/mask\[3\] digital/ins_024_ CMPO
+ VDD VSS digital/ins_049_ sg13g2f_ND3D1
Xdigital/ins_100_ digital/ins_028_ digital/ins_049_ digital/ins_030_
+ VDD VSS digital/ins_015_ sg13g2f_AOI21D1
Xdigital/ins_101_ digital/mask\[4\] digital/ins_024_ CMPO
+ VDD VSS digital/ins_050_ sg13g2f_ND3D1
Xdigital/ins_102_ digital/ins_029_ digital/ins_050_ digital/ins_030_
+ VDD VSS digital/ins_016_ sg13g2f_AOI21D1
Xdigital/ins_103_ digital/state\[1\] digital/state\[0\] VDD
+ VSS VALID sg13g2f_AN2D1
Xdigital/ins_104_ clknet_leaf_2_CLK digital/ins_000_ RESULTN\[0\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_105_ clknet_leaf_2_CLK digital/ins_001_ RESULTN\[1\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_106_ clknet_leaf_2_CLK digital/ins_002_ RESULTN\[2\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_107_ clknet_leaf_0_CLK digital/ins_003_ RESULTN\[3\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_108_ clknet_leaf_2_CLK digital/ins_004_ RESULTN\[4\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_109_ clknet_leaf_1_CLK digital/ins_005_ digital/mask\[0\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_110_ clknet_leaf_1_CLK digital/ins_006_ digital/mask\[1\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_111_ clknet_leaf_0_CLK digital/ins_007_ digital/mask\[2\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_112_ clknet_1_1__leaf_CLK digital/ins_008_ digital/mask\[3\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_113_ clknet_leaf_3_CLK digital/ins_009_ digital/mask\[4\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_114_ clknet_leaf_0_CLK digital/ins_010_ digital/state\[0\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_115_ clknet_leaf_0_CLK digital/ins_011_ digital/state\[1\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_116_ clknet_leaf_3_CLK digital/ins_012_ RESULT[0]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_117_ clknet_leaf_1_CLK digital/ins_013_ RESULT[1]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_118_ clknet_leaf_1_CLK digital/ins_014_ RESULT[2]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_119_ clknet_leaf_3_CLK digital/ins_015_ RESULT[3]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_120_ clknet_leaf_3_CLK digital/ins_016_ RESULT[4]
+ VDD VSS sg13g2f_DFQD1
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit_0_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit_0_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_0_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_0_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_1_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_1_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_2_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_2_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_3_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_3_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_4_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_4_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_5_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_5_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_6_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_6_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_7_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_7_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_8_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_8_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_9_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_9_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_10_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_10_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_11_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_11_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_12_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_12_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_13_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_13_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_14_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_14_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_15_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_15_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz2_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz2_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_7_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz2_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz2_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_7_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgn_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgn_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz2_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz2_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/sw_vouth2voutl_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_7_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_7_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/sw_vouth2voutl_SW_TAPBB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/sw_vouth2voutl_SW_TAPAA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit_0_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit_0_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_0_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_0_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_1_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_1_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_2_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_2_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_3_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_3_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_4_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_4_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_5_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_5_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_6_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_6_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_7_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_7_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_8_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_8_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_9_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_9_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_10_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_10_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_11_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_11_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_12_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_12_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_13_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_13_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_14_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_14_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_15_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_15_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xtapcell_up_inst_1 AVDD VSS sg13g2f_TAPCELL
Xtapcell_dw_inst_1 AVDD VSS sg13g2f_TAPCELL
Xtapcell_up_inst_3 AVDD VSS sg13g2f_TAPCELL
Xtapcell_dw_inst_3 AVDD VSS sg13g2f_TAPCELL
Xtapcell_up_inst_7 AVDD VSS sg13g2f_TAPCELL
Xtapcell_dw_inst_7 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_25_ANALOG_2_Left_0 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_26_ANALOG_2_Left_1 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_27_ANALOG_2_Left_2 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_22_ANALOG_Left_3 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_23_ANALOG_Left_4 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_24_ANALOG_Left_5 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_25_ANALOG_2_Right_6 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_22_ANALOG_Right_7 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_23_ANALOG_Right_8 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_24_ANALOG_Right_9 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_26_ANALOG_2_Right_10 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_27_ANALOG_2_Right_11 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_28_ANALOG_Right_12 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_29_ANALOG_Right_13 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_30_ANALOG_Right_14 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_28_ANALOG_Left_15 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_29_ANALOG_Left_16 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_30_ANALOG_Left_17 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_52_2_Right_18 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_51_2_Right_19 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_50_2_Right_20 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_49_2_Right_21 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_48_2_Right_22 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_47_2_Right_23 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_46_2_Right_24 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_45_2_Right_25 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_44_2_Right_26 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_43_2_Right_27 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_42_2_Right_28 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_41_2_Right_29 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_40_2_Right_30 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_39_2_Right_31 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_38_2_Right_32 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_37_2_Right_33 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_36_2_Right_34 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_35_2_Right_35 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_34_2_Right_36 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_33_2_Right_37 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_32_2_Right_38 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_31_2_Right_39 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_30_2_Right_40 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_29_2_Right_41 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_28_2_Right_42 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_27_2_Right_43 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_26_2_Right_44 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_25_2_Right_45 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_24_2_Right_46 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_23_2_Right_47 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_22_2_Right_48 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_21_2_Right_49 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_20_2_Right_50 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_19_2_Right_51 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_18_2_Right_52 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_17_2_Right_53 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_16_2_Right_54 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_15_2_Right_55 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_14_2_Right_56 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_13_2_Right_57 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_12_2_Right_58 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_11_2_Right_59 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_10_2_Right_60 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_9_2_Right_61 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_8_2_Right_62 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_7_2_Right_63 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_6_2_Right_64 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_5_2_Right_65 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_4_2_Right_66 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_3_2_Right_67 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_2_2_Right_68 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_1_2_Right_69 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_0_2_Right_70 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_52_2_Left_71 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_51_2_Left_72 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_50_2_Left_73 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_49_2_Left_74 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_48_2_Left_75 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_47_2_Left_76 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_46_2_Left_77 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_45_2_Left_78 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_44_2_Left_79 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_43_2_Left_80 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_42_2_Left_81 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_41_2_Left_82 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_40_2_Left_83 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_39_2_Left_84 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_38_2_Left_85 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_37_2_Left_86 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_36_2_Left_87 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_35_2_Left_88 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_34_2_Left_89 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_33_2_Left_90 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_32_2_Left_91 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_31_2_Left_92 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_30_2_Left_93 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_29_2_Left_94 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_28_2_Left_95 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_27_2_Left_96 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_26_2_Left_97 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_25_2_Left_98 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_24_2_Left_99 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_23_2_Left_100 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_22_2_Left_101 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_21_2_Left_102 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_20_2_Left_103 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_19_2_Left_104 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_18_2_Left_105 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_17_2_Left_106 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_16_2_Left_107 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_15_2_Left_108 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_14_2_Left_109 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_13_2_Left_110 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_12_2_Left_111 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_11_2_Left_112 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_10_2_Left_113 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_9_2_Left_114 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_8_2_Left_115 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_7_2_Left_116 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_6_2_Left_117 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_5_2_Left_118 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_4_2_Left_119 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_3_2_Left_120 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_2_2_Left_121 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_1_2_Left_122 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_0_2_Left_123 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_25_ANALOG_2_124 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_25_ANALOG_2_125 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_25_ANALOG_2_126 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_25_ANALOG_2_127 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_128 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_129 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_130 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_131 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_132 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_133 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_134 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_135 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_136 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_137 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_138 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_23_ANALOG_139 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_23_ANALOG_140 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_23_ANALOG_141 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_23_ANALOG_142 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_23_ANALOG_143 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_144 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_145 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_146 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_147 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_148 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_149 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_150 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_151 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_152 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_153 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_154 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_26_ANALOG_2_155 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_26_ANALOG_2_156 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_26_ANALOG_2_157 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_26_ANALOG_2_158 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_27_ANALOG_2_159 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_27_ANALOG_2_160 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_27_ANALOG_2_161 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_162 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_163 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_164 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_165 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_166 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_167 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_168 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_169 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_170 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_171 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_172 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_29_ANALOG_173 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_29_ANALOG_174 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_29_ANALOG_175 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_29_ANALOG_176 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_29_ANALOG_177 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_178 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_179 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_180 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_181 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_182 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_183 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_184 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_185 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_186 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_187 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_188 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_52_2_189 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_50_2_190 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_48_2_191 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_46_2_192 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_44_2_193 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_42_2_194 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_40_2_195 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_38_2_196 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_36_2_197 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_34_2_198 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_32_2_199 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_2_200 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_2_201 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_26_2_202 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_2_203 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_2_204 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_20_2_205 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_18_2_206 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_16_2_207 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_14_2_208 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_12_2_209 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_10_2_210 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_8_2_211 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_6_2_212 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_4_2_213 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_2_2_214 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_0_2_215 VDD VSS sg13g2f_TAPCELL
Xclkbuf_regs_0_CLK CLK VDD VSS CLK_regs sg13g2f_BUFFD1
Xclkbuf_leaf_0_CLK clknet_1_1__leaf_CLK VDD VSS clknet_leaf_0_CLK
+ sg13g2f_BUFFD1
Xclkbuf_leaf_1_CLK clknet_1_1__leaf_CLK VDD VSS clknet_leaf_1_CLK
+ sg13g2f_BUFFD1
Xclkbuf_leaf_2_CLK clknet_1_0__leaf_CLK VDD VSS clknet_leaf_2_CLK
+ sg13g2f_BUFFD1
Xclkbuf_leaf_3_CLK clknet_1_0__leaf_CLK VDD VSS clknet_leaf_3_CLK
+ sg13g2f_BUFFD1
Xclkbuf_0_CLK CLK VDD VSS clknet_0_CLK sg13g2f_BUFFD1
Xclkbuf_1_0__f_CLK clknet_0_CLK VDD VSS clknet_1_0__leaf_CLK
+ sg13g2f_BUFFD1
Xclkbuf_1_1__f_CLK clknet_0_CLK VDD VSS clknet_1_1__leaf_CLK
+ sg13g2f_BUFFD1
Xclkload0 clknet_1_0__leaf_CLK _unconnected_0 VSS VDD sg13g2f_INVD1
Xclkbuf_0_CLK_regs CLK_regs VDD VSS clknet_0_CLK_regs sg13g2f_BUFFD1
Xclkbuf_1_0__f_CLK_regs clknet_0_CLK_regs VDD VSS clknet_1_0__leaf_CLK_regs
+ sg13g2f_BUFFD1
XFILLER_0_1390 VDD VSS sg13g2f_FILL8
XFILLER_0_1398 VDD VSS sg13g2f_FILL8
XFILLER_0_1406 VDD VSS sg13g2f_FILL8
XFILLER_0_1414 VDD VSS sg13g2f_FILL8
XFILLER_0_1422 VDD VSS sg13g2f_FILL8
XFILLER_0_1430 VDD VSS sg13g2f_FILL8
XFILLER_0_1438 VDD VSS sg13g2f_FILL8
XFILLER_0_1446 VDD VSS sg13g2f_FILL8
XFILLER_0_1454 VDD VSS sg13g2f_FILL8
XFILLER_0_1462 VDD VSS sg13g2f_FILL8
XFILLER_0_1470 VDD VSS sg13g2f_FILL8
XFILLER_0_1478 VDD VSS sg13g2f_FILL8
XFILLER_0_1486 VDD VSS sg13g2f_FILL8
XFILLER_0_1494 VDD VSS sg13g2f_FILL1
XFILLER_0_1502 VDD VSS sg13g2f_FILL8
XFILLER_0_1510 VDD VSS sg13g2f_FILL8
XFILLER_0_1518 VDD VSS sg13g2f_FILL8
XFILLER_0_1526 VDD VSS sg13g2f_FILL8
XFILLER_0_1534 VDD VSS sg13g2f_FILL8
XFILLER_0_1542 VDD VSS sg13g2f_FILL8
XFILLER_0_1550 VDD VSS sg13g2f_FILL1
XFILLER_1_1390 VDD VSS sg13g2f_FILL8
XFILLER_1_1398 VDD VSS sg13g2f_FILL8
XFILLER_1_1406 VDD VSS sg13g2f_FILL8
XFILLER_1_1414 VDD VSS sg13g2f_FILL8
XFILLER_1_1422 VDD VSS sg13g2f_FILL8
XFILLER_1_1430 VDD VSS sg13g2f_FILL8
XFILLER_1_1438 VDD VSS sg13g2f_FILL8
XFILLER_1_1446 VDD VSS sg13g2f_FILL8
XFILLER_1_1454 VDD VSS sg13g2f_FILL8
XFILLER_1_1462 VDD VSS sg13g2f_FILL8
XFILLER_1_1470 VDD VSS sg13g2f_FILL8
XFILLER_1_1478 VDD VSS sg13g2f_FILL8
XFILLER_1_1486 VDD VSS sg13g2f_FILL8
XFILLER_1_1494 VDD VSS sg13g2f_FILL8
XFILLER_1_1502 VDD VSS sg13g2f_FILL8
XFILLER_1_1510 VDD VSS sg13g2f_FILL4
XFILLER_1_1514 VDD VSS sg13g2f_FILL1
XFILLER_1_1526 VDD VSS sg13g2f_FILL8
XFILLER_1_1534 VDD VSS sg13g2f_FILL8
XFILLER_1_1542 VDD VSS sg13g2f_FILL8
XFILLER_1_1550 VDD VSS sg13g2f_FILL1
XFILLER_2_1390 VDD VSS sg13g2f_FILL8
XFILLER_2_1398 VDD VSS sg13g2f_FILL8
XFILLER_2_1406 VDD VSS sg13g2f_FILL8
XFILLER_2_1414 VDD VSS sg13g2f_FILL8
XFILLER_2_1422 VDD VSS sg13g2f_FILL8
XFILLER_2_1430 VDD VSS sg13g2f_FILL8
XFILLER_2_1438 VDD VSS sg13g2f_FILL8
XFILLER_2_1446 VDD VSS sg13g2f_FILL8
XFILLER_2_1454 VDD VSS sg13g2f_FILL8
XFILLER_2_1462 VDD VSS sg13g2f_FILL8
XFILLER_2_1470 VDD VSS sg13g2f_FILL8
XFILLER_2_1478 VDD VSS sg13g2f_FILL8
XFILLER_2_1486 VDD VSS sg13g2f_FILL8
XFILLER_2_1494 VDD VSS sg13g2f_FILL4
XFILLER_2_1505 VDD VSS sg13g2f_FILL8
XFILLER_2_1513 VDD VSS sg13g2f_FILL8
XFILLER_2_1521 VDD VSS sg13g2f_FILL8
XFILLER_2_1529 VDD VSS sg13g2f_FILL8
XFILLER_2_1537 VDD VSS sg13g2f_FILL8
XFILLER_2_1545 VDD VSS sg13g2f_FILL4
XFILLER_2_1549 VDD VSS sg13g2f_FILL2
XFILLER_3_1390 VDD VSS sg13g2f_FILL8
XFILLER_3_1398 VDD VSS sg13g2f_FILL8
XFILLER_3_1406 VDD VSS sg13g2f_FILL8
XFILLER_3_1414 VDD VSS sg13g2f_FILL8
XFILLER_3_1422 VDD VSS sg13g2f_FILL8
XFILLER_3_1430 VDD VSS sg13g2f_FILL8
XFILLER_3_1438 VDD VSS sg13g2f_FILL8
XFILLER_3_1446 VDD VSS sg13g2f_FILL8
XFILLER_3_1454 VDD VSS sg13g2f_FILL8
XFILLER_3_1462 VDD VSS sg13g2f_FILL8
XFILLER_3_1470 VDD VSS sg13g2f_FILL8
XFILLER_3_1478 VDD VSS sg13g2f_FILL8
XFILLER_3_1486 VDD VSS sg13g2f_FILL8
XFILLER_3_1494 VDD VSS sg13g2f_FILL8
XFILLER_3_1502 VDD VSS sg13g2f_FILL2
XFILLER_3_1504 VDD VSS sg13g2f_FILL1
XFILLER_3_1537 VDD VSS sg13g2f_FILL8
XFILLER_3_1545 VDD VSS sg13g2f_FILL4
XFILLER_3_1549 VDD VSS sg13g2f_FILL2
XFILLER_4_1390 VDD VSS sg13g2f_FILL8
XFILLER_4_1398 VDD VSS sg13g2f_FILL8
XFILLER_4_1406 VDD VSS sg13g2f_FILL8
XFILLER_4_1414 VDD VSS sg13g2f_FILL8
XFILLER_4_1422 VDD VSS sg13g2f_FILL8
XFILLER_4_1430 VDD VSS sg13g2f_FILL8
XFILLER_4_1438 VDD VSS sg13g2f_FILL8
XFILLER_4_1446 VDD VSS sg13g2f_FILL8
XFILLER_4_1454 VDD VSS sg13g2f_FILL8
XFILLER_4_1462 VDD VSS sg13g2f_FILL8
XFILLER_4_1470 VDD VSS sg13g2f_FILL8
XFILLER_4_1478 VDD VSS sg13g2f_FILL8
XFILLER_4_1486 VDD VSS sg13g2f_FILL8
XFILLER_4_1494 VDD VSS sg13g2f_FILL4
XFILLER_4_1505 VDD VSS sg13g2f_FILL8
XFILLER_4_1513 VDD VSS sg13g2f_FILL2
XFILLER_4_1515 VDD VSS sg13g2f_FILL1
XFILLER_4_1527 VDD VSS sg13g2f_FILL8
XFILLER_4_1535 VDD VSS sg13g2f_FILL8
XFILLER_4_1543 VDD VSS sg13g2f_FILL8
XFILLER_5_1390 VDD VSS sg13g2f_FILL8
XFILLER_5_1398 VDD VSS sg13g2f_FILL8
XFILLER_5_1406 VDD VSS sg13g2f_FILL8
XFILLER_5_1414 VDD VSS sg13g2f_FILL8
XFILLER_5_1422 VDD VSS sg13g2f_FILL8
XFILLER_5_1430 VDD VSS sg13g2f_FILL8
XFILLER_5_1438 VDD VSS sg13g2f_FILL8
XFILLER_5_1446 VDD VSS sg13g2f_FILL8
XFILLER_5_1454 VDD VSS sg13g2f_FILL8
XFILLER_5_1462 VDD VSS sg13g2f_FILL8
XFILLER_5_1470 VDD VSS sg13g2f_FILL8
XFILLER_5_1478 VDD VSS sg13g2f_FILL8
XFILLER_5_1486 VDD VSS sg13g2f_FILL8
XFILLER_5_1494 VDD VSS sg13g2f_FILL4
XFILLER_5_1498 VDD VSS sg13g2f_FILL2
XFILLER_5_1500 VDD VSS sg13g2f_FILL1
XFILLER_5_1543 VDD VSS sg13g2f_FILL8
XFILLER_6_1390 VDD VSS sg13g2f_FILL8
XFILLER_6_1398 VDD VSS sg13g2f_FILL8
XFILLER_6_1406 VDD VSS sg13g2f_FILL8
XFILLER_6_1414 VDD VSS sg13g2f_FILL8
XFILLER_6_1422 VDD VSS sg13g2f_FILL8
XFILLER_6_1430 VDD VSS sg13g2f_FILL8
XFILLER_6_1438 VDD VSS sg13g2f_FILL8
XFILLER_6_1446 VDD VSS sg13g2f_FILL8
XFILLER_6_1454 VDD VSS sg13g2f_FILL8
XFILLER_6_1462 VDD VSS sg13g2f_FILL8
XFILLER_6_1470 VDD VSS sg13g2f_FILL8
XFILLER_6_1478 VDD VSS sg13g2f_FILL8
XFILLER_6_1486 VDD VSS sg13g2f_FILL8
XFILLER_6_1494 VDD VSS sg13g2f_FILL4
XFILLER_6_1547 VDD VSS sg13g2f_FILL4
XFILLER_7_1390 VDD VSS sg13g2f_FILL8
XFILLER_7_1398 VDD VSS sg13g2f_FILL8
XFILLER_7_1406 VDD VSS sg13g2f_FILL8
XFILLER_7_1414 VDD VSS sg13g2f_FILL8
XFILLER_7_1422 VDD VSS sg13g2f_FILL8
XFILLER_7_1430 VDD VSS sg13g2f_FILL8
XFILLER_7_1438 VDD VSS sg13g2f_FILL8
XFILLER_7_1446 VDD VSS sg13g2f_FILL8
XFILLER_7_1454 VDD VSS sg13g2f_FILL8
XFILLER_7_1462 VDD VSS sg13g2f_FILL8
XFILLER_7_1470 VDD VSS sg13g2f_FILL8
XFILLER_7_1478 VDD VSS sg13g2f_FILL8
XFILLER_7_1486 VDD VSS sg13g2f_FILL8
XFILLER_7_1494 VDD VSS sg13g2f_FILL8
XFILLER_7_1502 VDD VSS sg13g2f_FILL8
XFILLER_7_1510 VDD VSS sg13g2f_FILL8
XFILLER_7_1518 VDD VSS sg13g2f_FILL8
XFILLER_7_1526 VDD VSS sg13g2f_FILL8
XFILLER_7_1534 VDD VSS sg13g2f_FILL8
XFILLER_7_1542 VDD VSS sg13g2f_FILL8
XFILLER_7_1550 VDD VSS sg13g2f_FILL1
XFILLER_8_1390 VDD VSS sg13g2f_FILL8
XFILLER_8_1398 VDD VSS sg13g2f_FILL8
XFILLER_8_1406 VDD VSS sg13g2f_FILL8
XFILLER_8_1414 VDD VSS sg13g2f_FILL8
XFILLER_8_1422 VDD VSS sg13g2f_FILL8
XFILLER_8_1430 VDD VSS sg13g2f_FILL8
XFILLER_8_1438 VDD VSS sg13g2f_FILL8
XFILLER_8_1446 VDD VSS sg13g2f_FILL8
XFILLER_8_1454 VDD VSS sg13g2f_FILL8
XFILLER_8_1462 VDD VSS sg13g2f_FILL8
XFILLER_8_1470 VDD VSS sg13g2f_FILL8
XFILLER_8_1478 VDD VSS sg13g2f_FILL8
XFILLER_8_1486 VDD VSS sg13g2f_FILL8
XFILLER_8_1494 VDD VSS sg13g2f_FILL4
XFILLER_8_1547 VDD VSS sg13g2f_FILL4
XFILLER_9_1390 VDD VSS sg13g2f_FILL8
XFILLER_9_1398 VDD VSS sg13g2f_FILL8
XFILLER_9_1406 VDD VSS sg13g2f_FILL8
XFILLER_9_1414 VDD VSS sg13g2f_FILL8
XFILLER_9_1422 VDD VSS sg13g2f_FILL8
XFILLER_9_1430 VDD VSS sg13g2f_FILL8
XFILLER_9_1438 VDD VSS sg13g2f_FILL8
XFILLER_9_1446 VDD VSS sg13g2f_FILL8
XFILLER_9_1454 VDD VSS sg13g2f_FILL8
XFILLER_9_1462 VDD VSS sg13g2f_FILL8
XFILLER_9_1470 VDD VSS sg13g2f_FILL8
XFILLER_9_1478 VDD VSS sg13g2f_FILL8
XFILLER_9_1486 VDD VSS sg13g2f_FILL8
XFILLER_9_1494 VDD VSS sg13g2f_FILL8
XFILLER_9_1502 VDD VSS sg13g2f_FILL8
XFILLER_9_1510 VDD VSS sg13g2f_FILL8
XFILLER_9_1518 VDD VSS sg13g2f_FILL8
XFILLER_9_1526 VDD VSS sg13g2f_FILL8
XFILLER_9_1534 VDD VSS sg13g2f_FILL8
XFILLER_9_1542 VDD VSS sg13g2f_FILL8
XFILLER_9_1550 VDD VSS sg13g2f_FILL1
XFILLER_10_1390 VDD VSS sg13g2f_FILL8
XFILLER_10_1398 VDD VSS sg13g2f_FILL8
XFILLER_10_1406 VDD VSS sg13g2f_FILL8
XFILLER_10_1414 VDD VSS sg13g2f_FILL8
XFILLER_10_1422 VDD VSS sg13g2f_FILL8
XFILLER_10_1430 VDD VSS sg13g2f_FILL8
XFILLER_10_1438 VDD VSS sg13g2f_FILL8
XFILLER_10_1446 VDD VSS sg13g2f_FILL8
XFILLER_10_1454 VDD VSS sg13g2f_FILL8
XFILLER_10_1462 VDD VSS sg13g2f_FILL8
XFILLER_10_1470 VDD VSS sg13g2f_FILL8
XFILLER_10_1478 VDD VSS sg13g2f_FILL8
XFILLER_10_1486 VDD VSS sg13g2f_FILL8
XFILLER_10_1494 VDD VSS sg13g2f_FILL4
XFILLER_10_1538 VDD VSS sg13g2f_FILL8
XFILLER_10_1546 VDD VSS sg13g2f_FILL4
XFILLER_10_1550 VDD VSS sg13g2f_FILL1
XFILLER_11_1390 VDD VSS sg13g2f_FILL8
XFILLER_11_1398 VDD VSS sg13g2f_FILL8
XFILLER_11_1406 VDD VSS sg13g2f_FILL8
XFILLER_11_1414 VDD VSS sg13g2f_FILL8
XFILLER_11_1422 VDD VSS sg13g2f_FILL8
XFILLER_11_1430 VDD VSS sg13g2f_FILL8
XFILLER_11_1438 VDD VSS sg13g2f_FILL8
XFILLER_11_1446 VDD VSS sg13g2f_FILL8
XFILLER_11_1454 VDD VSS sg13g2f_FILL8
XFILLER_11_1462 VDD VSS sg13g2f_FILL8
XFILLER_11_1470 VDD VSS sg13g2f_FILL8
XFILLER_11_1478 VDD VSS sg13g2f_FILL4
XFILLER_11_1482 VDD VSS sg13g2f_FILL2
XFILLER_11_1484 VDD VSS sg13g2f_FILL1
XFILLER_11_1548 VDD VSS sg13g2f_FILL2
XFILLER_11_1550 VDD VSS sg13g2f_FILL1
XFILLER_12_1390 VDD VSS sg13g2f_FILL8
XFILLER_12_1398 VDD VSS sg13g2f_FILL8
XFILLER_12_1406 VDD VSS sg13g2f_FILL8
XFILLER_12_1414 VDD VSS sg13g2f_FILL8
XFILLER_12_1422 VDD VSS sg13g2f_FILL8
XFILLER_12_1430 VDD VSS sg13g2f_FILL8
XFILLER_12_1438 VDD VSS sg13g2f_FILL8
XFILLER_12_1446 VDD VSS sg13g2f_FILL8
XFILLER_12_1454 VDD VSS sg13g2f_FILL8
XFILLER_12_1462 VDD VSS sg13g2f_FILL8
XFILLER_12_1470 VDD VSS sg13g2f_FILL8
XFILLER_12_1478 VDD VSS sg13g2f_FILL8
XFILLER_12_1486 VDD VSS sg13g2f_FILL8
XFILLER_12_1494 VDD VSS sg13g2f_FILL4
XFILLER_12_1505 VDD VSS sg13g2f_FILL4
XFILLER_12_1536 VDD VSS sg13g2f_FILL2
XFILLER_12_1538 VDD VSS sg13g2f_FILL1
XFILLER_12_1547 VDD VSS sg13g2f_FILL4
XFILLER_13_1390 VDD VSS sg13g2f_FILL8
XFILLER_13_1398 VDD VSS sg13g2f_FILL8
XFILLER_13_1406 VDD VSS sg13g2f_FILL8
XFILLER_13_1414 VDD VSS sg13g2f_FILL8
XFILLER_13_1422 VDD VSS sg13g2f_FILL8
XFILLER_13_1430 VDD VSS sg13g2f_FILL8
XFILLER_13_1438 VDD VSS sg13g2f_FILL8
XFILLER_13_1446 VDD VSS sg13g2f_FILL8
XFILLER_13_1454 VDD VSS sg13g2f_FILL8
XFILLER_13_1462 VDD VSS sg13g2f_FILL8
XFILLER_13_1470 VDD VSS sg13g2f_FILL8
XFILLER_13_1478 VDD VSS sg13g2f_FILL8
XFILLER_13_1486 VDD VSS sg13g2f_FILL8
XFILLER_13_1494 VDD VSS sg13g2f_FILL4
XFILLER_13_1498 VDD VSS sg13g2f_FILL2
XFILLER_13_1542 VDD VSS sg13g2f_FILL8
XFILLER_13_1550 VDD VSS sg13g2f_FILL1
XFILLER_14_1390 VDD VSS sg13g2f_FILL8
XFILLER_14_1398 VDD VSS sg13g2f_FILL8
XFILLER_14_1406 VDD VSS sg13g2f_FILL8
XFILLER_14_1414 VDD VSS sg13g2f_FILL8
XFILLER_14_1422 VDD VSS sg13g2f_FILL8
XFILLER_14_1430 VDD VSS sg13g2f_FILL8
XFILLER_14_1438 VDD VSS sg13g2f_FILL8
XFILLER_14_1446 VDD VSS sg13g2f_FILL8
XFILLER_14_1454 VDD VSS sg13g2f_FILL8
XFILLER_14_1462 VDD VSS sg13g2f_FILL8
XFILLER_14_1470 VDD VSS sg13g2f_FILL8
XFILLER_14_1478 VDD VSS sg13g2f_FILL4
XFILLER_14_1482 VDD VSS sg13g2f_FILL2
XFILLER_14_1484 VDD VSS sg13g2f_FILL1
XFILLER_14_1547 VDD VSS sg13g2f_FILL4
XFILLER_15_1390 VDD VSS sg13g2f_FILL8
XFILLER_15_1398 VDD VSS sg13g2f_FILL8
XFILLER_15_1406 VDD VSS sg13g2f_FILL8
XFILLER_15_1414 VDD VSS sg13g2f_FILL8
XFILLER_15_1422 VDD VSS sg13g2f_FILL8
XFILLER_15_1430 VDD VSS sg13g2f_FILL8
XFILLER_15_1438 VDD VSS sg13g2f_FILL8
XFILLER_15_1446 VDD VSS sg13g2f_FILL8
XFILLER_15_1454 VDD VSS sg13g2f_FILL8
XFILLER_15_1462 VDD VSS sg13g2f_FILL8
XFILLER_15_1470 VDD VSS sg13g2f_FILL8
XFILLER_15_1478 VDD VSS sg13g2f_FILL8
XFILLER_15_1486 VDD VSS sg13g2f_FILL8
XFILLER_15_1494 VDD VSS sg13g2f_FILL8
XFILLER_15_1502 VDD VSS sg13g2f_FILL8
XFILLER_15_1510 VDD VSS sg13g2f_FILL4
XFILLER_15_1525 VDD VSS sg13g2f_FILL8
XFILLER_15_1533 VDD VSS sg13g2f_FILL8
XFILLER_15_1541 VDD VSS sg13g2f_FILL8
XFILLER_15_1549 VDD VSS sg13g2f_FILL2
XFILLER_16_1390 VDD VSS sg13g2f_FILL8
XFILLER_16_1398 VDD VSS sg13g2f_FILL8
XFILLER_16_1406 VDD VSS sg13g2f_FILL8
XFILLER_16_1414 VDD VSS sg13g2f_FILL8
XFILLER_16_1422 VDD VSS sg13g2f_FILL8
XFILLER_16_1430 VDD VSS sg13g2f_FILL8
XFILLER_16_1438 VDD VSS sg13g2f_FILL8
XFILLER_16_1446 VDD VSS sg13g2f_FILL8
XFILLER_16_1454 VDD VSS sg13g2f_FILL8
XFILLER_16_1462 VDD VSS sg13g2f_FILL8
XFILLER_16_1470 VDD VSS sg13g2f_FILL8
XFILLER_16_1478 VDD VSS sg13g2f_FILL8
XFILLER_16_1486 VDD VSS sg13g2f_FILL8
XFILLER_16_1494 VDD VSS sg13g2f_FILL4
XFILLER_16_1547 VDD VSS sg13g2f_FILL4
XFILLER_17_1390 VDD VSS sg13g2f_FILL8
XFILLER_17_1398 VDD VSS sg13g2f_FILL8
XFILLER_17_1406 VDD VSS sg13g2f_FILL8
XFILLER_17_1414 VDD VSS sg13g2f_FILL8
XFILLER_17_1422 VDD VSS sg13g2f_FILL8
XFILLER_17_1430 VDD VSS sg13g2f_FILL8
XFILLER_17_1438 VDD VSS sg13g2f_FILL8
XFILLER_17_1446 VDD VSS sg13g2f_FILL8
XFILLER_17_1454 VDD VSS sg13g2f_FILL8
XFILLER_17_1462 VDD VSS sg13g2f_FILL8
XFILLER_17_1470 VDD VSS sg13g2f_FILL8
XFILLER_17_1478 VDD VSS sg13g2f_FILL8
XFILLER_17_1486 VDD VSS sg13g2f_FILL8
XFILLER_17_1494 VDD VSS sg13g2f_FILL8
XFILLER_17_1502 VDD VSS sg13g2f_FILL8
XFILLER_17_1510 VDD VSS sg13g2f_FILL8
XFILLER_17_1518 VDD VSS sg13g2f_FILL8
XFILLER_17_1526 VDD VSS sg13g2f_FILL8
XFILLER_17_1534 VDD VSS sg13g2f_FILL8
XFILLER_17_1542 VDD VSS sg13g2f_FILL8
XFILLER_17_1550 VDD VSS sg13g2f_FILL1
XFILLER_18_1390 VDD VSS sg13g2f_FILL8
XFILLER_18_1398 VDD VSS sg13g2f_FILL8
XFILLER_18_1406 VDD VSS sg13g2f_FILL8
XFILLER_18_1414 VDD VSS sg13g2f_FILL8
XFILLER_18_1422 VDD VSS sg13g2f_FILL8
XFILLER_18_1430 VDD VSS sg13g2f_FILL8
XFILLER_18_1438 VDD VSS sg13g2f_FILL8
XFILLER_18_1446 VDD VSS sg13g2f_FILL8
XFILLER_18_1454 VDD VSS sg13g2f_FILL8
XFILLER_18_1462 VDD VSS sg13g2f_FILL8
XFILLER_18_1470 VDD VSS sg13g2f_FILL8
XFILLER_18_1478 VDD VSS sg13g2f_FILL8
XFILLER_18_1486 VDD VSS sg13g2f_FILL8
XFILLER_18_1494 VDD VSS sg13g2f_FILL4
XFILLER_18_1505 VDD VSS sg13g2f_FILL8
XFILLER_18_1513 VDD VSS sg13g2f_FILL8
XFILLER_18_1521 VDD VSS sg13g2f_FILL8
XFILLER_18_1529 VDD VSS sg13g2f_FILL8
XFILLER_18_1537 VDD VSS sg13g2f_FILL8
XFILLER_18_1545 VDD VSS sg13g2f_FILL4
XFILLER_18_1549 VDD VSS sg13g2f_FILL2
XFILLER_19_1390 VDD VSS sg13g2f_FILL8
XFILLER_19_1398 VDD VSS sg13g2f_FILL8
XFILLER_19_1406 VDD VSS sg13g2f_FILL8
XFILLER_19_1414 VDD VSS sg13g2f_FILL8
XFILLER_19_1422 VDD VSS sg13g2f_FILL8
XFILLER_19_1430 VDD VSS sg13g2f_FILL8
XFILLER_19_1438 VDD VSS sg13g2f_FILL8
XFILLER_19_1446 VDD VSS sg13g2f_FILL8
XFILLER_19_1454 VDD VSS sg13g2f_FILL8
XFILLER_19_1462 VDD VSS sg13g2f_FILL8
XFILLER_19_1470 VDD VSS sg13g2f_FILL8
XFILLER_19_1478 VDD VSS sg13g2f_FILL8
XFILLER_19_1486 VDD VSS sg13g2f_FILL8
XFILLER_19_1494 VDD VSS sg13g2f_FILL1
XFILLER_19_1530 VDD VSS sg13g2f_FILL8
XFILLER_19_1538 VDD VSS sg13g2f_FILL8
XFILLER_19_1546 VDD VSS sg13g2f_FILL4
XFILLER_19_1550 VDD VSS sg13g2f_FILL1
XFILLER_20_1390 VDD VSS sg13g2f_FILL8
XFILLER_20_1398 VDD VSS sg13g2f_FILL8
XFILLER_20_1406 VDD VSS sg13g2f_FILL8
XFILLER_20_1414 VDD VSS sg13g2f_FILL8
XFILLER_20_1422 VDD VSS sg13g2f_FILL8
XFILLER_20_1430 VDD VSS sg13g2f_FILL8
XFILLER_20_1438 VDD VSS sg13g2f_FILL8
XFILLER_20_1446 VDD VSS sg13g2f_FILL8
XFILLER_20_1454 VDD VSS sg13g2f_FILL8
XFILLER_20_1462 VDD VSS sg13g2f_FILL8
XFILLER_20_1470 VDD VSS sg13g2f_FILL8
XFILLER_20_1478 VDD VSS sg13g2f_FILL1
XFILLER_20_1505 VDD VSS sg13g2f_FILL2
XFILLER_20_1507 VDD VSS sg13g2f_FILL1
XFILLER_20_1538 VDD VSS sg13g2f_FILL8
XFILLER_20_1546 VDD VSS sg13g2f_FILL4
XFILLER_20_1550 VDD VSS sg13g2f_FILL1
XFILLER_21_1390 VDD VSS sg13g2f_FILL8
XFILLER_21_1398 VDD VSS sg13g2f_FILL8
XFILLER_21_1406 VDD VSS sg13g2f_FILL8
XFILLER_21_1414 VDD VSS sg13g2f_FILL8
XFILLER_21_1422 VDD VSS sg13g2f_FILL8
XFILLER_21_1430 VDD VSS sg13g2f_FILL8
XFILLER_21_1438 VDD VSS sg13g2f_FILL8
XFILLER_21_1446 VDD VSS sg13g2f_FILL8
XFILLER_21_1454 VDD VSS sg13g2f_FILL8
XFILLER_21_1462 VDD VSS sg13g2f_FILL8
XFILLER_21_1470 VDD VSS sg13g2f_FILL8
XFILLER_21_1478 VDD VSS sg13g2f_FILL8
XFILLER_21_1486 VDD VSS sg13g2f_FILL8
XFILLER_21_1494 VDD VSS sg13g2f_FILL8
XFILLER_21_1502 VDD VSS sg13g2f_FILL8
XFILLER_21_1510 VDD VSS sg13g2f_FILL8
XFILLER_21_1518 VDD VSS sg13g2f_FILL8
XFILLER_21_1526 VDD VSS sg13g2f_FILL8
XFILLER_21_1534 VDD VSS sg13g2f_FILL8
XFILLER_21_1542 VDD VSS sg13g2f_FILL8
XFILLER_21_1550 VDD VSS sg13g2f_FILL1
XFILLER_22_7 AVDD VSS sg13g2f_FILL4
XFILLER_22_11 AVDD VSS sg13g2f_FILL1
XFILLER_22_47 AVDD VSS sg13g2f_FILL1
XFILLER_22_119 AVDD VSS sg13g2f_FILL8
XFILLER_22_127 AVDD VSS sg13g2f_FILL8
XFILLER_22_135 AVDD VSS sg13g2f_FILL8
XFILLER_22_143 AVDD VSS sg13g2f_FILL8
XFILLER_22_151 AVDD VSS sg13g2f_FILL8
XFILLER_22_159 AVDD VSS sg13g2f_FILL8
XFILLER_22_167 AVDD VSS sg13g2f_FILL8
XFILLER_22_175 AVDD VSS sg13g2f_FILL8
XFILLER_22_183 AVDD VSS sg13g2f_FILL8
XFILLER_22_191 AVDD VSS sg13g2f_FILL8
XFILLER_22_199 AVDD VSS sg13g2f_FILL8
XFILLER_22_207 AVDD VSS sg13g2f_FILL8
XFILLER_22_215 AVDD VSS sg13g2f_FILL8
XFILLER_22_223 AVDD VSS sg13g2f_FILL1
XFILLER_22_231 AVDD VSS sg13g2f_FILL8
XFILLER_22_239 AVDD VSS sg13g2f_FILL8
XFILLER_22_247 AVDD VSS sg13g2f_FILL8
XFILLER_22_255 AVDD VSS sg13g2f_FILL8
XFILLER_22_263 AVDD VSS sg13g2f_FILL8
XFILLER_22_271 AVDD VSS sg13g2f_FILL8
XFILLER_22_279 AVDD VSS sg13g2f_FILL8
XFILLER_22_287 AVDD VSS sg13g2f_FILL8
XFILLER_22_295 AVDD VSS sg13g2f_FILL8
XFILLER_22_303 AVDD VSS sg13g2f_FILL8
XFILLER_22_311 AVDD VSS sg13g2f_FILL8
XFILLER_22_319 AVDD VSS sg13g2f_FILL8
XFILLER_22_327 AVDD VSS sg13g2f_FILL8
XFILLER_22_335 AVDD VSS sg13g2f_FILL1
XFILLER_22_343 AVDD VSS sg13g2f_FILL8
XFILLER_22_351 AVDD VSS sg13g2f_FILL8
XFILLER_22_359 AVDD VSS sg13g2f_FILL8
XFILLER_22_367 AVDD VSS sg13g2f_FILL8
XFILLER_22_375 AVDD VSS sg13g2f_FILL8
XFILLER_22_383 AVDD VSS sg13g2f_FILL1
XFILLER_22_455 AVDD VSS sg13g2f_FILL8
XFILLER_22_463 AVDD VSS sg13g2f_FILL8
XFILLER_22_471 AVDD VSS sg13g2f_FILL8
XFILLER_22_479 AVDD VSS sg13g2f_FILL8
XFILLER_22_487 AVDD VSS sg13g2f_FILL8
XFILLER_22_495 AVDD VSS sg13g2f_FILL8
XFILLER_22_503 AVDD VSS sg13g2f_FILL8
XFILLER_22_511 AVDD VSS sg13g2f_FILL8
XFILLER_22_519 AVDD VSS sg13g2f_FILL8
XFILLER_22_527 AVDD VSS sg13g2f_FILL8
XFILLER_22_535 AVDD VSS sg13g2f_FILL8
XFILLER_22_543 AVDD VSS sg13g2f_FILL8
XFILLER_22_551 AVDD VSS sg13g2f_FILL8
XFILLER_22_559 AVDD VSS sg13g2f_FILL1
XFILLER_22_567 AVDD VSS sg13g2f_FILL8
XFILLER_22_575 AVDD VSS sg13g2f_FILL8
XFILLER_22_583 AVDD VSS sg13g2f_FILL8
XFILLER_22_591 AVDD VSS sg13g2f_FILL8
XFILLER_22_599 AVDD VSS sg13g2f_FILL8
XFILLER_22_607 AVDD VSS sg13g2f_FILL8
XFILLER_22_615 AVDD VSS sg13g2f_FILL8
XFILLER_22_623 AVDD VSS sg13g2f_FILL8
XFILLER_22_631 AVDD VSS sg13g2f_FILL8
XFILLER_22_639 AVDD VSS sg13g2f_FILL8
XFILLER_22_647 AVDD VSS sg13g2f_FILL8
XFILLER_22_655 AVDD VSS sg13g2f_FILL8
XFILLER_22_663 AVDD VSS sg13g2f_FILL8
XFILLER_22_671 AVDD VSS sg13g2f_FILL1
XFILLER_22_679 AVDD VSS sg13g2f_FILL8
XFILLER_22_687 AVDD VSS sg13g2f_FILL8
XFILLER_22_695 AVDD VSS sg13g2f_FILL8
XFILLER_22_703 AVDD VSS sg13g2f_FILL8
XFILLER_22_711 AVDD VSS sg13g2f_FILL8
XFILLER_22_719 AVDD VSS sg13g2f_FILL8
XFILLER_22_727 AVDD VSS sg13g2f_FILL8
XFILLER_22_735 AVDD VSS sg13g2f_FILL8
XFILLER_22_743 AVDD VSS sg13g2f_FILL8
XFILLER_22_751 AVDD VSS sg13g2f_FILL8
XFILLER_22_759 AVDD VSS sg13g2f_FILL8
XFILLER_22_767 AVDD VSS sg13g2f_FILL8
XFILLER_22_775 AVDD VSS sg13g2f_FILL8
XFILLER_22_783 AVDD VSS sg13g2f_FILL1
XFILLER_22_791 AVDD VSS sg13g2f_FILL8
XFILLER_22_799 AVDD VSS sg13g2f_FILL8
XFILLER_22_807 AVDD VSS sg13g2f_FILL8
XFILLER_22_815 AVDD VSS sg13g2f_FILL8
XFILLER_22_823 AVDD VSS sg13g2f_FILL8
XFILLER_22_831 AVDD VSS sg13g2f_FILL8
XFILLER_22_839 AVDD VSS sg13g2f_FILL8
XFILLER_22_847 AVDD VSS sg13g2f_FILL8
XFILLER_22_855 AVDD VSS sg13g2f_FILL8
XFILLER_22_863 AVDD VSS sg13g2f_FILL8
XFILLER_22_871 AVDD VSS sg13g2f_FILL8
XFILLER_22_879 AVDD VSS sg13g2f_FILL8
XFILLER_22_887 AVDD VSS sg13g2f_FILL8
XFILLER_22_895 AVDD VSS sg13g2f_FILL1
XFILLER_22_903 AVDD VSS sg13g2f_FILL8
XFILLER_22_911 AVDD VSS sg13g2f_FILL8
XFILLER_22_919 AVDD VSS sg13g2f_FILL8
XFILLER_22_927 AVDD VSS sg13g2f_FILL8
XFILLER_22_935 AVDD VSS sg13g2f_FILL8
XFILLER_22_943 AVDD VSS sg13g2f_FILL8
XFILLER_22_951 AVDD VSS sg13g2f_FILL8
XFILLER_22_959 AVDD VSS sg13g2f_FILL8
XFILLER_22_967 AVDD VSS sg13g2f_FILL8
XFILLER_22_975 AVDD VSS sg13g2f_FILL8
XFILLER_22_983 AVDD VSS sg13g2f_FILL8
XFILLER_22_991 AVDD VSS sg13g2f_FILL8
XFILLER_22_999 AVDD VSS sg13g2f_FILL8
XFILLER_22_1007 AVDD VSS sg13g2f_FILL1
XFILLER_22_1015 AVDD VSS sg13g2f_FILL8
XFILLER_22_1023 AVDD VSS sg13g2f_FILL8
XFILLER_22_1031 AVDD VSS sg13g2f_FILL8
XFILLER_22_1039 AVDD VSS sg13g2f_FILL8
XFILLER_22_1047 AVDD VSS sg13g2f_FILL8
XFILLER_22_1055 AVDD VSS sg13g2f_FILL8
XFILLER_22_1063 AVDD VSS sg13g2f_FILL8
XFILLER_22_1071 AVDD VSS sg13g2f_FILL8
XFILLER_22_1079 AVDD VSS sg13g2f_FILL8
XFILLER_22_1087 AVDD VSS sg13g2f_FILL8
XFILLER_22_1095 AVDD VSS sg13g2f_FILL8
XFILLER_22_1103 AVDD VSS sg13g2f_FILL8
XFILLER_22_1111 AVDD VSS sg13g2f_FILL8
XFILLER_22_1119 AVDD VSS sg13g2f_FILL1
XFILLER_22_1127 AVDD VSS sg13g2f_FILL8
XFILLER_22_1135 AVDD VSS sg13g2f_FILL4
XFILLER_22_1139 AVDD VSS sg13g2f_FILL2
XFILLER_22_1152 AVDD VSS sg13g2f_FILL8
XFILLER_22_1160 AVDD VSS sg13g2f_FILL8
XFILLER_22_1168 AVDD VSS sg13g2f_FILL8
XFILLER_22_1176 AVDD VSS sg13g2f_FILL8
XFILLER_22_1184 AVDD VSS sg13g2f_FILL8
XFILLER_22_1192 AVDD VSS sg13g2f_FILL8
XFILLER_22_1200 AVDD VSS sg13g2f_FILL8
XFILLER_22_1208 AVDD VSS sg13g2f_FILL8
XFILLER_22_1216 AVDD VSS sg13g2f_FILL8
XFILLER_22_1224 AVDD VSS sg13g2f_FILL8
XFILLER_22_1239 AVDD VSS sg13g2f_FILL8
XFILLER_22_1247 AVDD VSS sg13g2f_FILL8
XFILLER_22_1255 AVDD VSS sg13g2f_FILL8
XFILLER_22_1263 AVDD VSS sg13g2f_FILL4
XFILLER_22_1267 AVDD VSS sg13g2f_FILL1
XFILLER_22_1390 VDD VSS sg13g2f_FILL8
XFILLER_22_1398 VDD VSS sg13g2f_FILL8
XFILLER_22_1406 VDD VSS sg13g2f_FILL8
XFILLER_22_1414 VDD VSS sg13g2f_FILL8
XFILLER_22_1422 VDD VSS sg13g2f_FILL8
XFILLER_22_1430 VDD VSS sg13g2f_FILL8
XFILLER_22_1438 VDD VSS sg13g2f_FILL8
XFILLER_22_1446 VDD VSS sg13g2f_FILL8
XFILLER_22_1454 VDD VSS sg13g2f_FILL8
XFILLER_22_1462 VDD VSS sg13g2f_FILL8
XFILLER_22_1470 VDD VSS sg13g2f_FILL8
XFILLER_22_1478 VDD VSS sg13g2f_FILL8
XFILLER_22_1486 VDD VSS sg13g2f_FILL8
XFILLER_22_1494 VDD VSS sg13g2f_FILL4
XFILLER_22_1547 VDD VSS sg13g2f_FILL4
XFILLER_23_7 AVDD VSS sg13g2f_FILL4
XFILLER_23_11 AVDD VSS sg13g2f_FILL1
XFILLER_23_58 AVDD VSS sg13g2f_FILL4
XFILLER_23_126 AVDD VSS sg13g2f_FILL8
XFILLER_23_134 AVDD VSS sg13g2f_FILL8
XFILLER_23_142 AVDD VSS sg13g2f_FILL8
XFILLER_23_150 AVDD VSS sg13g2f_FILL8
XFILLER_23_158 AVDD VSS sg13g2f_FILL8
XFILLER_23_166 AVDD VSS sg13g2f_FILL8
XFILLER_23_174 AVDD VSS sg13g2f_FILL8
XFILLER_23_182 AVDD VSS sg13g2f_FILL8
XFILLER_23_190 AVDD VSS sg13g2f_FILL8
XFILLER_23_198 AVDD VSS sg13g2f_FILL8
XFILLER_23_206 AVDD VSS sg13g2f_FILL8
XFILLER_23_214 AVDD VSS sg13g2f_FILL8
XFILLER_23_222 AVDD VSS sg13g2f_FILL8
XFILLER_23_230 AVDD VSS sg13g2f_FILL1
XFILLER_23_238 AVDD VSS sg13g2f_FILL8
XFILLER_23_246 AVDD VSS sg13g2f_FILL8
XFILLER_23_254 AVDD VSS sg13g2f_FILL8
XFILLER_23_262 AVDD VSS sg13g2f_FILL8
XFILLER_23_270 AVDD VSS sg13g2f_FILL8
XFILLER_23_278 AVDD VSS sg13g2f_FILL8
XFILLER_23_286 AVDD VSS sg13g2f_FILL8
XFILLER_23_294 AVDD VSS sg13g2f_FILL8
XFILLER_23_302 AVDD VSS sg13g2f_FILL8
XFILLER_23_310 AVDD VSS sg13g2f_FILL8
XFILLER_23_318 AVDD VSS sg13g2f_FILL8
XFILLER_23_326 AVDD VSS sg13g2f_FILL8
XFILLER_23_334 AVDD VSS sg13g2f_FILL8
XFILLER_23_342 AVDD VSS sg13g2f_FILL8
XFILLER_23_350 AVDD VSS sg13g2f_FILL8
XFILLER_23_358 AVDD VSS sg13g2f_FILL8
XFILLER_23_366 AVDD VSS sg13g2f_FILL8
XFILLER_23_374 AVDD VSS sg13g2f_FILL8
XFILLER_23_382 AVDD VSS sg13g2f_FILL8
XFILLER_23_390 AVDD VSS sg13g2f_FILL4
XFILLER_23_394 AVDD VSS sg13g2f_FILL1
XFILLER_23_459 AVDD VSS sg13g2f_FILL2
XFILLER_23_461 AVDD VSS sg13g2f_FILL1
XFILLER_23_469 AVDD VSS sg13g2f_FILL8
XFILLER_23_477 AVDD VSS sg13g2f_FILL8
XFILLER_23_485 AVDD VSS sg13g2f_FILL8
XFILLER_23_493 AVDD VSS sg13g2f_FILL8
XFILLER_23_501 AVDD VSS sg13g2f_FILL8
XFILLER_23_509 AVDD VSS sg13g2f_FILL8
XFILLER_23_517 AVDD VSS sg13g2f_FILL8
XFILLER_23_525 AVDD VSS sg13g2f_FILL8
XFILLER_23_533 AVDD VSS sg13g2f_FILL8
XFILLER_23_541 AVDD VSS sg13g2f_FILL8
XFILLER_23_549 AVDD VSS sg13g2f_FILL8
XFILLER_23_557 AVDD VSS sg13g2f_FILL1
XFILLER_23_622 AVDD VSS sg13g2f_FILL8
XFILLER_23_630 AVDD VSS sg13g2f_FILL8
XFILLER_23_638 AVDD VSS sg13g2f_FILL8
XFILLER_23_646 AVDD VSS sg13g2f_FILL8
XFILLER_23_654 AVDD VSS sg13g2f_FILL8
XFILLER_23_662 AVDD VSS sg13g2f_FILL8
XFILLER_23_670 AVDD VSS sg13g2f_FILL8
XFILLER_23_678 AVDD VSS sg13g2f_FILL8
XFILLER_23_686 AVDD VSS sg13g2f_FILL4
XFILLER_23_690 AVDD VSS sg13g2f_FILL2
XFILLER_23_692 AVDD VSS sg13g2f_FILL1
XFILLER_23_700 AVDD VSS sg13g2f_FILL8
XFILLER_23_708 AVDD VSS sg13g2f_FILL8
XFILLER_23_716 AVDD VSS sg13g2f_FILL8
XFILLER_23_724 AVDD VSS sg13g2f_FILL8
XFILLER_23_732 AVDD VSS sg13g2f_FILL8
XFILLER_23_740 AVDD VSS sg13g2f_FILL8
XFILLER_23_748 AVDD VSS sg13g2f_FILL8
XFILLER_23_756 AVDD VSS sg13g2f_FILL8
XFILLER_23_764 AVDD VSS sg13g2f_FILL8
XFILLER_23_772 AVDD VSS sg13g2f_FILL8
XFILLER_23_780 AVDD VSS sg13g2f_FILL8
XFILLER_23_788 AVDD VSS sg13g2f_FILL8
XFILLER_23_796 AVDD VSS sg13g2f_FILL8
XFILLER_23_804 AVDD VSS sg13g2f_FILL8
XFILLER_23_812 AVDD VSS sg13g2f_FILL8
XFILLER_23_820 AVDD VSS sg13g2f_FILL8
XFILLER_23_828 AVDD VSS sg13g2f_FILL8
XFILLER_23_836 AVDD VSS sg13g2f_FILL8
XFILLER_23_844 AVDD VSS sg13g2f_FILL8
XFILLER_23_868 AVDD VSS sg13g2f_FILL8
XFILLER_23_876 AVDD VSS sg13g2f_FILL4
XFILLER_23_905 AVDD VSS sg13g2f_FILL8
XFILLER_23_913 AVDD VSS sg13g2f_FILL8
XFILLER_23_921 AVDD VSS sg13g2f_FILL2
XFILLER_23_923 AVDD VSS sg13g2f_FILL1
XFILLER_23_931 AVDD VSS sg13g2f_FILL8
XFILLER_23_939 AVDD VSS sg13g2f_FILL8
XFILLER_23_947 AVDD VSS sg13g2f_FILL8
XFILLER_23_955 AVDD VSS sg13g2f_FILL8
XFILLER_23_963 AVDD VSS sg13g2f_FILL8
XFILLER_23_971 AVDD VSS sg13g2f_FILL8
XFILLER_23_979 AVDD VSS sg13g2f_FILL8
XFILLER_23_987 AVDD VSS sg13g2f_FILL8
XFILLER_23_995 AVDD VSS sg13g2f_FILL8
XFILLER_23_1003 AVDD VSS sg13g2f_FILL8
XFILLER_23_1011 AVDD VSS sg13g2f_FILL8
XFILLER_23_1019 AVDD VSS sg13g2f_FILL2
XFILLER_23_1021 AVDD VSS sg13g2f_FILL1
XFILLER_23_1038 AVDD VSS sg13g2f_FILL8
XFILLER_23_1110 AVDD VSS sg13g2f_FILL8
XFILLER_23_1118 AVDD VSS sg13g2f_FILL8
XFILLER_23_1126 AVDD VSS sg13g2f_FILL8
XFILLER_23_1150 AVDD VSS sg13g2f_FILL4
XFILLER_23_1154 AVDD VSS sg13g2f_FILL1
XFILLER_23_1162 AVDD VSS sg13g2f_FILL8
XFILLER_23_1170 AVDD VSS sg13g2f_FILL8
XFILLER_23_1178 AVDD VSS sg13g2f_FILL8
XFILLER_23_1186 AVDD VSS sg13g2f_FILL8
XFILLER_23_1194 AVDD VSS sg13g2f_FILL8
XFILLER_23_1202 AVDD VSS sg13g2f_FILL8
XFILLER_23_1210 AVDD VSS sg13g2f_FILL8
XFILLER_23_1218 AVDD VSS sg13g2f_FILL8
XFILLER_23_1226 AVDD VSS sg13g2f_FILL8
XFILLER_23_1234 AVDD VSS sg13g2f_FILL8
XFILLER_23_1242 AVDD VSS sg13g2f_FILL8
XFILLER_23_1250 AVDD VSS sg13g2f_FILL8
XFILLER_23_1258 AVDD VSS sg13g2f_FILL8
XFILLER_23_1266 AVDD VSS sg13g2f_FILL2
XFILLER_23_1390 VDD VSS sg13g2f_FILL8
XFILLER_23_1398 VDD VSS sg13g2f_FILL8
XFILLER_23_1406 VDD VSS sg13g2f_FILL8
XFILLER_23_1414 VDD VSS sg13g2f_FILL8
XFILLER_23_1422 VDD VSS sg13g2f_FILL8
XFILLER_23_1430 VDD VSS sg13g2f_FILL8
XFILLER_23_1438 VDD VSS sg13g2f_FILL8
XFILLER_23_1446 VDD VSS sg13g2f_FILL8
XFILLER_23_1454 VDD VSS sg13g2f_FILL8
XFILLER_23_1462 VDD VSS sg13g2f_FILL8
XFILLER_23_1470 VDD VSS sg13g2f_FILL8
XFILLER_23_1478 VDD VSS sg13g2f_FILL8
XFILLER_23_1486 VDD VSS sg13g2f_FILL8
XFILLER_23_1494 VDD VSS sg13g2f_FILL8
XFILLER_23_1502 VDD VSS sg13g2f_FILL1
XFILLER_23_1545 VDD VSS sg13g2f_FILL4
XFILLER_23_1549 VDD VSS sg13g2f_FILL2
XFILLER_24_7 AVDD VSS sg13g2f_FILL4
XFILLER_24_11 AVDD VSS sg13g2f_FILL1
XFILLER_24_119 AVDD VSS sg13g2f_FILL8
XFILLER_24_127 AVDD VSS sg13g2f_FILL8
XFILLER_24_135 AVDD VSS sg13g2f_FILL8
XFILLER_24_143 AVDD VSS sg13g2f_FILL8
XFILLER_24_151 AVDD VSS sg13g2f_FILL8
XFILLER_24_159 AVDD VSS sg13g2f_FILL8
XFILLER_24_167 AVDD VSS sg13g2f_FILL8
XFILLER_24_175 AVDD VSS sg13g2f_FILL8
XFILLER_24_183 AVDD VSS sg13g2f_FILL8
XFILLER_24_191 AVDD VSS sg13g2f_FILL8
XFILLER_24_199 AVDD VSS sg13g2f_FILL8
XFILLER_24_207 AVDD VSS sg13g2f_FILL8
XFILLER_24_215 AVDD VSS sg13g2f_FILL8
XFILLER_24_223 AVDD VSS sg13g2f_FILL1
XFILLER_24_247 AVDD VSS sg13g2f_FILL8
XFILLER_24_255 AVDD VSS sg13g2f_FILL8
XFILLER_24_263 AVDD VSS sg13g2f_FILL8
XFILLER_24_271 AVDD VSS sg13g2f_FILL8
XFILLER_24_279 AVDD VSS sg13g2f_FILL8
XFILLER_24_287 AVDD VSS sg13g2f_FILL8
XFILLER_24_295 AVDD VSS sg13g2f_FILL8
XFILLER_24_303 AVDD VSS sg13g2f_FILL8
XFILLER_24_311 AVDD VSS sg13g2f_FILL8
XFILLER_24_319 AVDD VSS sg13g2f_FILL8
XFILLER_24_327 AVDD VSS sg13g2f_FILL8
XFILLER_24_335 AVDD VSS sg13g2f_FILL1
XFILLER_24_343 AVDD VSS sg13g2f_FILL8
XFILLER_24_351 AVDD VSS sg13g2f_FILL1
XFILLER_24_374 AVDD VSS sg13g2f_FILL8
XFILLER_24_382 AVDD VSS sg13g2f_FILL2
XFILLER_24_455 AVDD VSS sg13g2f_FILL8
XFILLER_24_463 AVDD VSS sg13g2f_FILL8
XFILLER_24_471 AVDD VSS sg13g2f_FILL8
XFILLER_24_479 AVDD VSS sg13g2f_FILL8
XFILLER_24_487 AVDD VSS sg13g2f_FILL8
XFILLER_24_495 AVDD VSS sg13g2f_FILL8
XFILLER_24_503 AVDD VSS sg13g2f_FILL8
XFILLER_24_511 AVDD VSS sg13g2f_FILL8
XFILLER_24_519 AVDD VSS sg13g2f_FILL8
XFILLER_24_527 AVDD VSS sg13g2f_FILL8
XFILLER_24_535 AVDD VSS sg13g2f_FILL8
XFILLER_24_543 AVDD VSS sg13g2f_FILL8
XFILLER_24_551 AVDD VSS sg13g2f_FILL8
XFILLER_24_559 AVDD VSS sg13g2f_FILL1
XFILLER_24_567 AVDD VSS sg13g2f_FILL8
XFILLER_24_575 AVDD VSS sg13g2f_FILL8
XFILLER_24_583 AVDD VSS sg13g2f_FILL8
XFILLER_24_591 AVDD VSS sg13g2f_FILL8
XFILLER_24_599 AVDD VSS sg13g2f_FILL8
XFILLER_24_607 AVDD VSS sg13g2f_FILL8
XFILLER_24_615 AVDD VSS sg13g2f_FILL8
XFILLER_24_623 AVDD VSS sg13g2f_FILL8
XFILLER_24_631 AVDD VSS sg13g2f_FILL8
XFILLER_24_639 AVDD VSS sg13g2f_FILL8
XFILLER_24_647 AVDD VSS sg13g2f_FILL8
XFILLER_24_655 AVDD VSS sg13g2f_FILL8
XFILLER_24_663 AVDD VSS sg13g2f_FILL8
XFILLER_24_671 AVDD VSS sg13g2f_FILL1
XFILLER_24_679 AVDD VSS sg13g2f_FILL2
XFILLER_24_681 AVDD VSS sg13g2f_FILL1
XFILLER_24_746 AVDD VSS sg13g2f_FILL8
XFILLER_24_754 AVDD VSS sg13g2f_FILL8
XFILLER_24_762 AVDD VSS sg13g2f_FILL8
XFILLER_24_770 AVDD VSS sg13g2f_FILL8
XFILLER_24_778 AVDD VSS sg13g2f_FILL4
XFILLER_24_782 AVDD VSS sg13g2f_FILL2
XFILLER_24_855 AVDD VSS sg13g2f_FILL8
XFILLER_24_863 AVDD VSS sg13g2f_FILL8
XFILLER_24_871 AVDD VSS sg13g2f_FILL8
XFILLER_24_879 AVDD VSS sg13g2f_FILL1
XFILLER_24_928 AVDD VSS sg13g2f_FILL2
XFILLER_24_994 AVDD VSS sg13g2f_FILL8
XFILLER_24_1002 AVDD VSS sg13g2f_FILL4
XFILLER_24_1006 AVDD VSS sg13g2f_FILL2
XFILLER_24_1101 AVDD VSS sg13g2f_FILL4
XFILLER_24_1105 AVDD VSS sg13g2f_FILL2
XFILLER_24_1118 AVDD VSS sg13g2f_FILL2
XFILLER_24_1127 AVDD VSS sg13g2f_FILL1
XFILLER_24_1153 AVDD VSS sg13g2f_FILL4
XFILLER_24_1198 AVDD VSS sg13g2f_FILL8
XFILLER_24_1206 AVDD VSS sg13g2f_FILL8
XFILLER_24_1214 AVDD VSS sg13g2f_FILL8
XFILLER_24_1222 AVDD VSS sg13g2f_FILL8
XFILLER_24_1230 AVDD VSS sg13g2f_FILL2
XFILLER_24_1239 AVDD VSS sg13g2f_FILL8
XFILLER_24_1247 AVDD VSS sg13g2f_FILL8
XFILLER_24_1255 AVDD VSS sg13g2f_FILL8
XFILLER_24_1263 AVDD VSS sg13g2f_FILL4
XFILLER_24_1267 AVDD VSS sg13g2f_FILL1
XFILLER_24_1398 VDD VSS sg13g2f_FILL8
XFILLER_24_1406 VDD VSS sg13g2f_FILL8
XFILLER_24_1414 VDD VSS sg13g2f_FILL8
XFILLER_24_1422 VDD VSS sg13g2f_FILL8
XFILLER_24_1430 VDD VSS sg13g2f_FILL8
XFILLER_24_1438 VDD VSS sg13g2f_FILL8
XFILLER_24_1446 VDD VSS sg13g2f_FILL8
XFILLER_24_1454 VDD VSS sg13g2f_FILL8
XFILLER_24_1462 VDD VSS sg13g2f_FILL8
XFILLER_24_1470 VDD VSS sg13g2f_FILL8
XFILLER_24_1478 VDD VSS sg13g2f_FILL8
XFILLER_24_1486 VDD VSS sg13g2f_FILL8
XFILLER_24_1494 VDD VSS sg13g2f_FILL4
XFILLER_24_1513 VDD VSS sg13g2f_FILL8
XFILLER_24_1521 VDD VSS sg13g2f_FILL8
XFILLER_24_1529 VDD VSS sg13g2f_FILL8
XFILLER_24_1537 VDD VSS sg13g2f_FILL8
XFILLER_24_1545 VDD VSS sg13g2f_FILL4
XFILLER_24_1549 VDD VSS sg13g2f_FILL2
XFILLER_25_151 AVDD VSS sg13g2f_FILL8
XFILLER_25_159 AVDD VSS sg13g2f_FILL8
XFILLER_25_167 AVDD VSS sg13g2f_FILL8
XFILLER_25_175 AVDD VSS sg13g2f_FILL4
XFILLER_25_179 AVDD VSS sg13g2f_FILL1
XFILLER_25_205 AVDD VSS sg13g2f_FILL8
XFILLER_25_238 AVDD VSS sg13g2f_FILL8
XFILLER_25_246 AVDD VSS sg13g2f_FILL8
XFILLER_25_254 AVDD VSS sg13g2f_FILL8
XFILLER_25_262 AVDD VSS sg13g2f_FILL2
XFILLER_25_289 AVDD VSS sg13g2f_FILL8
XFILLER_25_297 AVDD VSS sg13g2f_FILL8
XFILLER_25_305 AVDD VSS sg13g2f_FILL8
XFILLER_25_313 AVDD VSS sg13g2f_FILL4
XFILLER_25_317 AVDD VSS sg13g2f_FILL2
XFILLER_25_319 AVDD VSS sg13g2f_FILL1
XFILLER_25_336 AVDD VSS sg13g2f_FILL2
XFILLER_25_368 AVDD VSS sg13g2f_FILL4
XFILLER_25_372 AVDD VSS sg13g2f_FILL2
XFILLER_25_374 AVDD VSS sg13g2f_FILL1
XFILLER_25_382 AVDD VSS sg13g2f_FILL2
XFILLER_25_427 AVDD VSS sg13g2f_FILL4
XFILLER_25_431 AVDD VSS sg13g2f_FILL2
XFILLER_25_433 AVDD VSS sg13g2f_FILL1
XFILLER_25_498 AVDD VSS sg13g2f_FILL8
XFILLER_25_506 AVDD VSS sg13g2f_FILL8
XFILLER_25_514 AVDD VSS sg13g2f_FILL8
XFILLER_25_522 AVDD VSS sg13g2f_FILL8
XFILLER_25_530 AVDD VSS sg13g2f_FILL8
XFILLER_25_538 AVDD VSS sg13g2f_FILL2
XFILLER_25_540 AVDD VSS sg13g2f_FILL1
XFILLER_25_605 AVDD VSS sg13g2f_FILL1
XFILLER_25_613 AVDD VSS sg13g2f_FILL8
XFILLER_25_621 AVDD VSS sg13g2f_FILL8
XFILLER_25_629 AVDD VSS sg13g2f_FILL2
XFILLER_25_631 AVDD VSS sg13g2f_FILL1
XFILLER_25_665 AVDD VSS sg13g2f_FILL8
XFILLER_25_673 AVDD VSS sg13g2f_FILL2
XFILLER_25_675 AVDD VSS sg13g2f_FILL1
XFILLER_25_740 AVDD VSS sg13g2f_FILL8
XFILLER_25_748 AVDD VSS sg13g2f_FILL8
XFILLER_25_820 AVDD VSS sg13g2f_FILL1
XFILLER_25_844 AVDD VSS sg13g2f_FILL1
XFILLER_25_870 AVDD VSS sg13g2f_FILL8
XFILLER_25_878 AVDD VSS sg13g2f_FILL2
XFILLER_25_960 AVDD VSS sg13g2f_FILL4
XFILLER_25_964 AVDD VSS sg13g2f_FILL1
XFILLER_25_986 AVDD VSS sg13g2f_FILL8
XFILLER_25_994 AVDD VSS sg13g2f_FILL8
XFILLER_25_1002 AVDD VSS sg13g2f_FILL8
XFILLER_25_1010 AVDD VSS sg13g2f_FILL4
XFILLER_25_1014 AVDD VSS sg13g2f_FILL2
XFILLER_25_1041 AVDD VSS sg13g2f_FILL2
XFILLER_25_1116 AVDD VSS sg13g2f_FILL8
XFILLER_25_1124 AVDD VSS sg13g2f_FILL4
XFILLER_25_1139 AVDD VSS sg13g2f_FILL2
XFILLER_25_1141 AVDD VSS sg13g2f_FILL1
XFILLER_25_1206 AVDD VSS sg13g2f_FILL8
XFILLER_25_1214 AVDD VSS sg13g2f_FILL8
XFILLER_25_1222 AVDD VSS sg13g2f_FILL8
XFILLER_25_1230 AVDD VSS sg13g2f_FILL8
XFILLER_25_1238 AVDD VSS sg13g2f_FILL8
XFILLER_25_1246 AVDD VSS sg13g2f_FILL8
XFILLER_25_1254 AVDD VSS sg13g2f_FILL8
XFILLER_25_1262 AVDD VSS sg13g2f_FILL4
XFILLER_25_1266 AVDD VSS sg13g2f_FILL2
XFILLER_25_1390 VDD VSS sg13g2f_FILL8
XFILLER_25_1398 VDD VSS sg13g2f_FILL8
XFILLER_25_1406 VDD VSS sg13g2f_FILL8
XFILLER_25_1414 VDD VSS sg13g2f_FILL8
XFILLER_25_1422 VDD VSS sg13g2f_FILL8
XFILLER_25_1430 VDD VSS sg13g2f_FILL8
XFILLER_25_1438 VDD VSS sg13g2f_FILL8
XFILLER_25_1446 VDD VSS sg13g2f_FILL8
XFILLER_25_1454 VDD VSS sg13g2f_FILL8
XFILLER_25_1462 VDD VSS sg13g2f_FILL8
XFILLER_25_1470 VDD VSS sg13g2f_FILL8
XFILLER_25_1478 VDD VSS sg13g2f_FILL8
XFILLER_25_1486 VDD VSS sg13g2f_FILL8
XFILLER_25_1494 VDD VSS sg13g2f_FILL8
XFILLER_25_1502 VDD VSS sg13g2f_FILL8
XFILLER_25_1510 VDD VSS sg13g2f_FILL4
XFILLER_25_1514 VDD VSS sg13g2f_FILL2
XFILLER_25_1535 VDD VSS sg13g2f_FILL8
XFILLER_25_1543 VDD VSS sg13g2f_FILL8
XFILLER_26_405 AVDD VSS sg13g2f_FILL4
XFILLER_26_409 AVDD VSS sg13g2f_FILL1
XFILLER_26_497 AVDD VSS sg13g2f_FILL8
XFILLER_26_505 AVDD VSS sg13g2f_FILL2
XFILLER_26_507 AVDD VSS sg13g2f_FILL1
XFILLER_26_524 AVDD VSS sg13g2f_FILL8
XFILLER_26_532 AVDD VSS sg13g2f_FILL1
XFILLER_26_622 AVDD VSS sg13g2f_FILL8
XFILLER_26_630 AVDD VSS sg13g2f_FILL8
XFILLER_26_638 AVDD VSS sg13g2f_FILL2
XFILLER_26_656 AVDD VSS sg13g2f_FILL1
XFILLER_26_744 AVDD VSS sg13g2f_FILL8
XFILLER_26_752 AVDD VSS sg13g2f_FILL4
XFILLER_26_772 AVDD VSS sg13g2f_FILL1
XFILLER_26_846 AVDD VSS sg13g2f_FILL4
XFILLER_26_850 AVDD VSS sg13g2f_FILL1
XFILLER_26_870 AVDD VSS sg13g2f_FILL8
XFILLER_26_878 AVDD VSS sg13g2f_FILL2
XFILLER_26_937 AVDD VSS sg13g2f_FILL4
XFILLER_26_970 AVDD VSS sg13g2f_FILL8
XFILLER_26_994 AVDD VSS sg13g2f_FILL8
XFILLER_26_1002 AVDD VSS sg13g2f_FILL8
XFILLER_26_1010 AVDD VSS sg13g2f_FILL8
XFILLER_26_1099 AVDD VSS sg13g2f_FILL8
XFILLER_26_1107 AVDD VSS sg13g2f_FILL8
XFILLER_26_1115 AVDD VSS sg13g2f_FILL8
XFILLER_26_1123 AVDD VSS sg13g2f_FILL8
XFILLER_26_1131 AVDD VSS sg13g2f_FILL4
XFILLER_26_1135 AVDD VSS sg13g2f_FILL2
XFILLER_26_1162 AVDD VSS sg13g2f_FILL2
XFILLER_26_1190 AVDD VSS sg13g2f_FILL8
XFILLER_26_1198 AVDD VSS sg13g2f_FILL4
XFILLER_26_1202 AVDD VSS sg13g2f_FILL2
XFILLER_26_1406 VDD VSS sg13g2f_FILL8
XFILLER_26_1414 VDD VSS sg13g2f_FILL8
XFILLER_26_1422 VDD VSS sg13g2f_FILL8
XFILLER_26_1430 VDD VSS sg13g2f_FILL8
XFILLER_26_1438 VDD VSS sg13g2f_FILL8
XFILLER_26_1446 VDD VSS sg13g2f_FILL8
XFILLER_26_1454 VDD VSS sg13g2f_FILL8
XFILLER_26_1462 VDD VSS sg13g2f_FILL8
XFILLER_26_1470 VDD VSS sg13g2f_FILL8
XFILLER_26_1478 VDD VSS sg13g2f_FILL4
XFILLER_26_1496 VDD VSS sg13g2f_FILL2
XFILLER_26_1547 VDD VSS sg13g2f_FILL4
XFILLER_27_430 AVDD VSS sg13g2f_FILL4
XFILLER_27_498 AVDD VSS sg13g2f_FILL8
XFILLER_27_506 AVDD VSS sg13g2f_FILL2
XFILLER_27_513 AVDD VSS sg13g2f_FILL4
XFILLER_27_613 AVDD VSS sg13g2f_FILL8
XFILLER_27_621 AVDD VSS sg13g2f_FILL8
XFILLER_27_629 AVDD VSS sg13g2f_FILL2
XFILLER_27_631 AVDD VSS sg13g2f_FILL1
XFILLER_27_665 AVDD VSS sg13g2f_FILL1
XFILLER_27_746 AVDD VSS sg13g2f_FILL8
XFILLER_27_754 AVDD VSS sg13g2f_FILL2
XFILLER_27_831 AVDD VSS sg13g2f_FILL4
XFILLER_27_835 AVDD VSS sg13g2f_FILL2
XFILLER_27_860 AVDD VSS sg13g2f_FILL8
XFILLER_27_868 AVDD VSS sg13g2f_FILL8
XFILLER_27_876 AVDD VSS sg13g2f_FILL4
XFILLER_27_880 AVDD VSS sg13g2f_FILL2
XFILLER_27_907 AVDD VSS sg13g2f_FILL8
XFILLER_27_915 AVDD VSS sg13g2f_FILL2
XFILLER_27_917 AVDD VSS sg13g2f_FILL1
XFILLER_27_987 AVDD VSS sg13g2f_FILL8
XFILLER_27_995 AVDD VSS sg13g2f_FILL8
XFILLER_27_1003 AVDD VSS sg13g2f_FILL4
XFILLER_27_1007 AVDD VSS sg13g2f_FILL2
XFILLER_27_1020 AVDD VSS sg13g2f_FILL2
XFILLER_27_1022 AVDD VSS sg13g2f_FILL1
XFILLER_27_1066 AVDD VSS sg13g2f_FILL2
XFILLER_27_1118 AVDD VSS sg13g2f_FILL8
XFILLER_27_1126 AVDD VSS sg13g2f_FILL2
XFILLER_27_1192 AVDD VSS sg13g2f_FILL8
XFILLER_27_1200 AVDD VSS sg13g2f_FILL8
XFILLER_27_1208 AVDD VSS sg13g2f_FILL8
XFILLER_27_1216 AVDD VSS sg13g2f_FILL8
XFILLER_27_1224 AVDD VSS sg13g2f_FILL8
XFILLER_27_1232 AVDD VSS sg13g2f_FILL8
XFILLER_27_1240 AVDD VSS sg13g2f_FILL8
XFILLER_27_1248 AVDD VSS sg13g2f_FILL8
XFILLER_27_1256 AVDD VSS sg13g2f_FILL8
XFILLER_27_1264 AVDD VSS sg13g2f_FILL4
XFILLER_27_1390 VDD VSS sg13g2f_FILL8
XFILLER_27_1398 VDD VSS sg13g2f_FILL8
XFILLER_27_1406 VDD VSS sg13g2f_FILL8
XFILLER_27_1414 VDD VSS sg13g2f_FILL8
XFILLER_27_1422 VDD VSS sg13g2f_FILL8
XFILLER_27_1430 VDD VSS sg13g2f_FILL8
XFILLER_27_1438 VDD VSS sg13g2f_FILL8
XFILLER_27_1446 VDD VSS sg13g2f_FILL8
XFILLER_27_1454 VDD VSS sg13g2f_FILL8
XFILLER_27_1462 VDD VSS sg13g2f_FILL8
XFILLER_27_1470 VDD VSS sg13g2f_FILL4
XFILLER_27_1516 VDD VSS sg13g2f_FILL8
XFILLER_27_1524 VDD VSS sg13g2f_FILL8
XFILLER_27_1532 VDD VSS sg13g2f_FILL8
XFILLER_27_1540 VDD VSS sg13g2f_FILL8
XFILLER_27_1548 VDD VSS sg13g2f_FILL2
XFILLER_27_1550 VDD VSS sg13g2f_FILL1
XFILLER_28_7 AVDD VSS sg13g2f_FILL4
XFILLER_28_11 AVDD VSS sg13g2f_FILL2
XFILLER_28_124 AVDD VSS sg13g2f_FILL8
XFILLER_28_132 AVDD VSS sg13g2f_FILL4
XFILLER_28_136 AVDD VSS sg13g2f_FILL2
XFILLER_28_138 AVDD VSS sg13g2f_FILL1
XFILLER_28_155 AVDD VSS sg13g2f_FILL2
XFILLER_28_190 AVDD VSS sg13g2f_FILL8
XFILLER_28_198 AVDD VSS sg13g2f_FILL8
XFILLER_28_206 AVDD VSS sg13g2f_FILL8
XFILLER_28_214 AVDD VSS sg13g2f_FILL8
XFILLER_28_222 AVDD VSS sg13g2f_FILL2
XFILLER_28_231 AVDD VSS sg13g2f_FILL8
XFILLER_28_239 AVDD VSS sg13g2f_FILL8
XFILLER_28_247 AVDD VSS sg13g2f_FILL8
XFILLER_28_255 AVDD VSS sg13g2f_FILL8
XFILLER_28_263 AVDD VSS sg13g2f_FILL8
XFILLER_28_271 AVDD VSS sg13g2f_FILL8
XFILLER_28_279 AVDD VSS sg13g2f_FILL8
XFILLER_28_287 AVDD VSS sg13g2f_FILL4
XFILLER_28_291 AVDD VSS sg13g2f_FILL2
XFILLER_28_293 AVDD VSS sg13g2f_FILL1
XFILLER_28_305 AVDD VSS sg13g2f_FILL8
XFILLER_28_313 AVDD VSS sg13g2f_FILL8
XFILLER_28_321 AVDD VSS sg13g2f_FILL8
XFILLER_28_329 AVDD VSS sg13g2f_FILL4
XFILLER_28_333 AVDD VSS sg13g2f_FILL2
XFILLER_28_335 AVDD VSS sg13g2f_FILL1
XFILLER_28_343 AVDD VSS sg13g2f_FILL4
XFILLER_28_374 AVDD VSS sg13g2f_FILL8
XFILLER_28_382 AVDD VSS sg13g2f_FILL2
XFILLER_28_455 AVDD VSS sg13g2f_FILL8
XFILLER_28_463 AVDD VSS sg13g2f_FILL1
XFILLER_28_496 AVDD VSS sg13g2f_FILL8
XFILLER_28_504 AVDD VSS sg13g2f_FILL8
XFILLER_28_512 AVDD VSS sg13g2f_FILL8
XFILLER_28_520 AVDD VSS sg13g2f_FILL4
XFILLER_28_567 AVDD VSS sg13g2f_FILL4
XFILLER_28_571 AVDD VSS sg13g2f_FILL2
XFILLER_28_573 AVDD VSS sg13g2f_FILL1
XFILLER_28_593 AVDD VSS sg13g2f_FILL4
XFILLER_28_597 AVDD VSS sg13g2f_FILL1
XFILLER_28_617 AVDD VSS sg13g2f_FILL8
XFILLER_28_625 AVDD VSS sg13g2f_FILL4
XFILLER_28_629 AVDD VSS sg13g2f_FILL2
XFILLER_28_631 AVDD VSS sg13g2f_FILL1
XFILLER_28_643 AVDD VSS sg13g2f_FILL8
XFILLER_28_651 AVDD VSS sg13g2f_FILL2
XFILLER_28_653 AVDD VSS sg13g2f_FILL1
XFILLER_28_670 AVDD VSS sg13g2f_FILL2
XFILLER_28_743 AVDD VSS sg13g2f_FILL8
XFILLER_28_751 AVDD VSS sg13g2f_FILL4
XFILLER_28_755 AVDD VSS sg13g2f_FILL1
XFILLER_28_778 AVDD VSS sg13g2f_FILL4
XFILLER_28_782 AVDD VSS sg13g2f_FILL2
XFILLER_28_791 AVDD VSS sg13g2f_FILL8
XFILLER_28_799 AVDD VSS sg13g2f_FILL4
XFILLER_28_803 AVDD VSS sg13g2f_FILL2
XFILLER_28_805 AVDD VSS sg13g2f_FILL1
XFILLER_28_870 AVDD VSS sg13g2f_FILL8
XFILLER_28_878 AVDD VSS sg13g2f_FILL2
XFILLER_28_891 AVDD VSS sg13g2f_FILL4
XFILLER_28_895 AVDD VSS sg13g2f_FILL1
XFILLER_28_914 AVDD VSS sg13g2f_FILL1
XFILLER_28_990 AVDD VSS sg13g2f_FILL8
XFILLER_28_998 AVDD VSS sg13g2f_FILL8
XFILLER_28_1006 AVDD VSS sg13g2f_FILL2
XFILLER_28_1015 AVDD VSS sg13g2f_FILL1
XFILLER_28_1059 AVDD VSS sg13g2f_FILL4
XFILLER_28_1063 AVDD VSS sg13g2f_FILL2
XFILLER_28_1081 AVDD VSS sg13g2f_FILL1
XFILLER_28_1118 AVDD VSS sg13g2f_FILL2
XFILLER_28_1127 AVDD VSS sg13g2f_FILL1
XFILLER_28_1182 AVDD VSS sg13g2f_FILL8
XFILLER_28_1190 AVDD VSS sg13g2f_FILL8
XFILLER_28_1198 AVDD VSS sg13g2f_FILL8
XFILLER_28_1206 AVDD VSS sg13g2f_FILL8
XFILLER_28_1214 AVDD VSS sg13g2f_FILL8
XFILLER_28_1222 AVDD VSS sg13g2f_FILL8
XFILLER_28_1230 AVDD VSS sg13g2f_FILL2
XFILLER_28_1239 AVDD VSS sg13g2f_FILL8
XFILLER_28_1247 AVDD VSS sg13g2f_FILL8
XFILLER_28_1255 AVDD VSS sg13g2f_FILL8
XFILLER_28_1263 AVDD VSS sg13g2f_FILL4
XFILLER_28_1267 AVDD VSS sg13g2f_FILL1
XFILLER_28_1390 VDD VSS sg13g2f_FILL8
XFILLER_28_1398 VDD VSS sg13g2f_FILL8
XFILLER_28_1406 VDD VSS sg13g2f_FILL8
XFILLER_28_1414 VDD VSS sg13g2f_FILL8
XFILLER_28_1422 VDD VSS sg13g2f_FILL8
XFILLER_28_1430 VDD VSS sg13g2f_FILL8
XFILLER_28_1438 VDD VSS sg13g2f_FILL8
XFILLER_28_1446 VDD VSS sg13g2f_FILL8
XFILLER_28_1454 VDD VSS sg13g2f_FILL8
XFILLER_28_1462 VDD VSS sg13g2f_FILL8
XFILLER_28_1470 VDD VSS sg13g2f_FILL8
XFILLER_28_1478 VDD VSS sg13g2f_FILL8
XFILLER_28_1486 VDD VSS sg13g2f_FILL1
XFILLER_28_1513 VDD VSS sg13g2f_FILL8
XFILLER_28_1521 VDD VSS sg13g2f_FILL8
XFILLER_28_1529 VDD VSS sg13g2f_FILL8
XFILLER_28_1537 VDD VSS sg13g2f_FILL8
XFILLER_28_1545 VDD VSS sg13g2f_FILL4
XFILLER_28_1549 VDD VSS sg13g2f_FILL2
XFILLER_29_7 AVDD VSS sg13g2f_FILL4
XFILLER_29_11 AVDD VSS sg13g2f_FILL1
XFILLER_29_76 AVDD VSS sg13g2f_FILL8
XFILLER_29_84 AVDD VSS sg13g2f_FILL8
XFILLER_29_92 AVDD VSS sg13g2f_FILL8
XFILLER_29_100 AVDD VSS sg13g2f_FILL8
XFILLER_29_108 AVDD VSS sg13g2f_FILL8
XFILLER_29_116 AVDD VSS sg13g2f_FILL8
XFILLER_29_124 AVDD VSS sg13g2f_FILL8
XFILLER_29_132 AVDD VSS sg13g2f_FILL4
XFILLER_29_152 AVDD VSS sg13g2f_FILL4
XFILLER_29_156 AVDD VSS sg13g2f_FILL1
XFILLER_29_168 AVDD VSS sg13g2f_FILL8
XFILLER_29_176 AVDD VSS sg13g2f_FILL8
XFILLER_29_184 AVDD VSS sg13g2f_FILL8
XFILLER_29_192 AVDD VSS sg13g2f_FILL8
XFILLER_29_200 AVDD VSS sg13g2f_FILL8
XFILLER_29_208 AVDD VSS sg13g2f_FILL8
XFILLER_29_216 AVDD VSS sg13g2f_FILL8
XFILLER_29_224 AVDD VSS sg13g2f_FILL4
XFILLER_29_228 AVDD VSS sg13g2f_FILL2
XFILLER_29_230 AVDD VSS sg13g2f_FILL1
XFILLER_29_238 AVDD VSS sg13g2f_FILL8
XFILLER_29_246 AVDD VSS sg13g2f_FILL8
XFILLER_29_254 AVDD VSS sg13g2f_FILL8
XFILLER_29_262 AVDD VSS sg13g2f_FILL8
XFILLER_29_270 AVDD VSS sg13g2f_FILL8
XFILLER_29_278 AVDD VSS sg13g2f_FILL8
XFILLER_29_286 AVDD VSS sg13g2f_FILL8
XFILLER_29_294 AVDD VSS sg13g2f_FILL8
XFILLER_29_302 AVDD VSS sg13g2f_FILL8
XFILLER_29_310 AVDD VSS sg13g2f_FILL8
XFILLER_29_318 AVDD VSS sg13g2f_FILL8
XFILLER_29_326 AVDD VSS sg13g2f_FILL8
XFILLER_29_334 AVDD VSS sg13g2f_FILL8
XFILLER_29_342 AVDD VSS sg13g2f_FILL8
XFILLER_29_350 AVDD VSS sg13g2f_FILL8
XFILLER_29_358 AVDD VSS sg13g2f_FILL1
XFILLER_29_364 AVDD VSS sg13g2f_FILL8
XFILLER_29_372 AVDD VSS sg13g2f_FILL8
XFILLER_29_380 AVDD VSS sg13g2f_FILL4
XFILLER_29_448 AVDD VSS sg13g2f_FILL2
XFILLER_29_450 AVDD VSS sg13g2f_FILL1
XFILLER_29_485 AVDD VSS sg13g2f_FILL8
XFILLER_29_493 AVDD VSS sg13g2f_FILL8
XFILLER_29_501 AVDD VSS sg13g2f_FILL8
XFILLER_29_509 AVDD VSS sg13g2f_FILL4
XFILLER_29_593 AVDD VSS sg13g2f_FILL4
XFILLER_29_613 AVDD VSS sg13g2f_FILL8
XFILLER_29_621 AVDD VSS sg13g2f_FILL8
XFILLER_29_629 AVDD VSS sg13g2f_FILL8
XFILLER_29_637 AVDD VSS sg13g2f_FILL8
XFILLER_29_645 AVDD VSS sg13g2f_FILL8
XFILLER_29_653 AVDD VSS sg13g2f_FILL8
XFILLER_29_661 AVDD VSS sg13g2f_FILL1
XFILLER_29_673 AVDD VSS sg13g2f_FILL4
XFILLER_29_741 AVDD VSS sg13g2f_FILL8
XFILLER_29_749 AVDD VSS sg13g2f_FILL8
XFILLER_29_757 AVDD VSS sg13g2f_FILL8
XFILLER_29_765 AVDD VSS sg13g2f_FILL8
XFILLER_29_773 AVDD VSS sg13g2f_FILL8
XFILLER_29_781 AVDD VSS sg13g2f_FILL8
XFILLER_29_789 AVDD VSS sg13g2f_FILL4
XFILLER_29_793 AVDD VSS sg13g2f_FILL2
XFILLER_29_827 AVDD VSS sg13g2f_FILL2
XFILLER_29_829 AVDD VSS sg13g2f_FILL1
XFILLER_29_855 AVDD VSS sg13g2f_FILL2
XFILLER_29_868 AVDD VSS sg13g2f_FILL8
XFILLER_29_876 AVDD VSS sg13g2f_FILL8
XFILLER_29_909 AVDD VSS sg13g2f_FILL4
XFILLER_29_931 AVDD VSS sg13g2f_FILL8
XFILLER_29_939 AVDD VSS sg13g2f_FILL8
XFILLER_29_947 AVDD VSS sg13g2f_FILL1
XFILLER_29_991 AVDD VSS sg13g2f_FILL8
XFILLER_29_999 AVDD VSS sg13g2f_FILL8
XFILLER_29_1007 AVDD VSS sg13g2f_FILL4
XFILLER_29_1011 AVDD VSS sg13g2f_FILL2
XFILLER_29_1013 AVDD VSS sg13g2f_FILL1
XFILLER_29_1047 AVDD VSS sg13g2f_FILL8
XFILLER_29_1055 AVDD VSS sg13g2f_FILL8
XFILLER_29_1063 AVDD VSS sg13g2f_FILL8
XFILLER_29_1071 AVDD VSS sg13g2f_FILL4
XFILLER_29_1118 AVDD VSS sg13g2f_FILL8
XFILLER_29_1126 AVDD VSS sg13g2f_FILL8
XFILLER_29_1134 AVDD VSS sg13g2f_FILL1
XFILLER_29_1151 AVDD VSS sg13g2f_FILL4
XFILLER_29_1173 AVDD VSS sg13g2f_FILL8
XFILLER_29_1181 AVDD VSS sg13g2f_FILL8
XFILLER_29_1189 AVDD VSS sg13g2f_FILL8
XFILLER_29_1197 AVDD VSS sg13g2f_FILL8
XFILLER_29_1205 AVDD VSS sg13g2f_FILL8
XFILLER_29_1213 AVDD VSS sg13g2f_FILL8
XFILLER_29_1221 AVDD VSS sg13g2f_FILL8
XFILLER_29_1229 AVDD VSS sg13g2f_FILL8
XFILLER_29_1237 AVDD VSS sg13g2f_FILL8
XFILLER_29_1245 AVDD VSS sg13g2f_FILL8
XFILLER_29_1253 AVDD VSS sg13g2f_FILL8
XFILLER_29_1261 AVDD VSS sg13g2f_FILL4
XFILLER_29_1265 AVDD VSS sg13g2f_FILL2
XFILLER_29_1267 AVDD VSS sg13g2f_FILL1
XFILLER_29_1390 VDD VSS sg13g2f_FILL8
XFILLER_29_1398 VDD VSS sg13g2f_FILL8
XFILLER_29_1406 VDD VSS sg13g2f_FILL8
XFILLER_29_1414 VDD VSS sg13g2f_FILL8
XFILLER_29_1422 VDD VSS sg13g2f_FILL8
XFILLER_29_1430 VDD VSS sg13g2f_FILL8
XFILLER_29_1438 VDD VSS sg13g2f_FILL8
XFILLER_29_1446 VDD VSS sg13g2f_FILL8
XFILLER_29_1454 VDD VSS sg13g2f_FILL8
XFILLER_29_1462 VDD VSS sg13g2f_FILL8
XFILLER_29_1470 VDD VSS sg13g2f_FILL4
XFILLER_29_1474 VDD VSS sg13g2f_FILL1
XFILLER_29_1528 VDD VSS sg13g2f_FILL8
XFILLER_29_1536 VDD VSS sg13g2f_FILL8
XFILLER_29_1544 VDD VSS sg13g2f_FILL4
XFILLER_29_1548 VDD VSS sg13g2f_FILL2
XFILLER_29_1550 VDD VSS sg13g2f_FILL1
XFILLER_30_7 AVDD VSS sg13g2f_FILL8
XFILLER_30_15 AVDD VSS sg13g2f_FILL8
XFILLER_30_23 AVDD VSS sg13g2f_FILL2
XFILLER_30_25 AVDD VSS sg13g2f_FILL1
XFILLER_30_47 AVDD VSS sg13g2f_FILL1
XFILLER_30_119 AVDD VSS sg13g2f_FILL8
XFILLER_30_127 AVDD VSS sg13g2f_FILL8
XFILLER_30_135 AVDD VSS sg13g2f_FILL8
XFILLER_30_143 AVDD VSS sg13g2f_FILL8
XFILLER_30_151 AVDD VSS sg13g2f_FILL8
XFILLER_30_159 AVDD VSS sg13g2f_FILL8
XFILLER_30_167 AVDD VSS sg13g2f_FILL8
XFILLER_30_175 AVDD VSS sg13g2f_FILL8
XFILLER_30_183 AVDD VSS sg13g2f_FILL8
XFILLER_30_191 AVDD VSS sg13g2f_FILL8
XFILLER_30_199 AVDD VSS sg13g2f_FILL8
XFILLER_30_207 AVDD VSS sg13g2f_FILL8
XFILLER_30_215 AVDD VSS sg13g2f_FILL8
XFILLER_30_223 AVDD VSS sg13g2f_FILL1
XFILLER_30_231 AVDD VSS sg13g2f_FILL8
XFILLER_30_239 AVDD VSS sg13g2f_FILL8
XFILLER_30_247 AVDD VSS sg13g2f_FILL8
XFILLER_30_255 AVDD VSS sg13g2f_FILL8
XFILLER_30_263 AVDD VSS sg13g2f_FILL8
XFILLER_30_271 AVDD VSS sg13g2f_FILL8
XFILLER_30_279 AVDD VSS sg13g2f_FILL8
XFILLER_30_287 AVDD VSS sg13g2f_FILL8
XFILLER_30_295 AVDD VSS sg13g2f_FILL8
XFILLER_30_303 AVDD VSS sg13g2f_FILL8
XFILLER_30_311 AVDD VSS sg13g2f_FILL8
XFILLER_30_319 AVDD VSS sg13g2f_FILL8
XFILLER_30_327 AVDD VSS sg13g2f_FILL8
XFILLER_30_335 AVDD VSS sg13g2f_FILL1
XFILLER_30_343 AVDD VSS sg13g2f_FILL8
XFILLER_30_351 AVDD VSS sg13g2f_FILL8
XFILLER_30_359 AVDD VSS sg13g2f_FILL8
XFILLER_30_367 AVDD VSS sg13g2f_FILL8
XFILLER_30_375 AVDD VSS sg13g2f_FILL8
XFILLER_30_383 AVDD VSS sg13g2f_FILL1
XFILLER_30_455 AVDD VSS sg13g2f_FILL1
XFILLER_30_467 AVDD VSS sg13g2f_FILL8
XFILLER_30_475 AVDD VSS sg13g2f_FILL8
XFILLER_30_483 AVDD VSS sg13g2f_FILL8
XFILLER_30_491 AVDD VSS sg13g2f_FILL8
XFILLER_30_499 AVDD VSS sg13g2f_FILL8
XFILLER_30_507 AVDD VSS sg13g2f_FILL8
XFILLER_30_515 AVDD VSS sg13g2f_FILL8
XFILLER_30_523 AVDD VSS sg13g2f_FILL8
XFILLER_30_531 AVDD VSS sg13g2f_FILL8
XFILLER_30_539 AVDD VSS sg13g2f_FILL8
XFILLER_30_547 AVDD VSS sg13g2f_FILL8
XFILLER_30_555 AVDD VSS sg13g2f_FILL4
XFILLER_30_559 AVDD VSS sg13g2f_FILL1
XFILLER_30_567 AVDD VSS sg13g2f_FILL8
XFILLER_30_575 AVDD VSS sg13g2f_FILL8
XFILLER_30_583 AVDD VSS sg13g2f_FILL8
XFILLER_30_591 AVDD VSS sg13g2f_FILL8
XFILLER_30_599 AVDD VSS sg13g2f_FILL8
XFILLER_30_607 AVDD VSS sg13g2f_FILL8
XFILLER_30_615 AVDD VSS sg13g2f_FILL8
XFILLER_30_623 AVDD VSS sg13g2f_FILL8
XFILLER_30_631 AVDD VSS sg13g2f_FILL8
XFILLER_30_639 AVDD VSS sg13g2f_FILL8
XFILLER_30_647 AVDD VSS sg13g2f_FILL8
XFILLER_30_655 AVDD VSS sg13g2f_FILL8
XFILLER_30_663 AVDD VSS sg13g2f_FILL8
XFILLER_30_671 AVDD VSS sg13g2f_FILL1
XFILLER_30_679 AVDD VSS sg13g2f_FILL8
XFILLER_30_687 AVDD VSS sg13g2f_FILL8
XFILLER_30_695 AVDD VSS sg13g2f_FILL8
XFILLER_30_714 AVDD VSS sg13g2f_FILL8
XFILLER_30_722 AVDD VSS sg13g2f_FILL8
XFILLER_30_730 AVDD VSS sg13g2f_FILL8
XFILLER_30_738 AVDD VSS sg13g2f_FILL8
XFILLER_30_746 AVDD VSS sg13g2f_FILL8
XFILLER_30_754 AVDD VSS sg13g2f_FILL8
XFILLER_30_762 AVDD VSS sg13g2f_FILL8
XFILLER_30_770 AVDD VSS sg13g2f_FILL8
XFILLER_30_778 AVDD VSS sg13g2f_FILL4
XFILLER_30_782 AVDD VSS sg13g2f_FILL2
XFILLER_30_791 AVDD VSS sg13g2f_FILL8
XFILLER_30_799 AVDD VSS sg13g2f_FILL8
XFILLER_30_807 AVDD VSS sg13g2f_FILL8
XFILLER_30_815 AVDD VSS sg13g2f_FILL8
XFILLER_30_823 AVDD VSS sg13g2f_FILL8
XFILLER_30_831 AVDD VSS sg13g2f_FILL8
XFILLER_30_839 AVDD VSS sg13g2f_FILL8
XFILLER_30_847 AVDD VSS sg13g2f_FILL8
XFILLER_30_855 AVDD VSS sg13g2f_FILL8
XFILLER_30_863 AVDD VSS sg13g2f_FILL8
XFILLER_30_871 AVDD VSS sg13g2f_FILL8
XFILLER_30_879 AVDD VSS sg13g2f_FILL8
XFILLER_30_887 AVDD VSS sg13g2f_FILL8
XFILLER_30_895 AVDD VSS sg13g2f_FILL1
XFILLER_30_903 AVDD VSS sg13g2f_FILL8
XFILLER_30_911 AVDD VSS sg13g2f_FILL8
XFILLER_30_919 AVDD VSS sg13g2f_FILL8
XFILLER_30_927 AVDD VSS sg13g2f_FILL8
XFILLER_30_935 AVDD VSS sg13g2f_FILL8
XFILLER_30_943 AVDD VSS sg13g2f_FILL8
XFILLER_30_951 AVDD VSS sg13g2f_FILL8
XFILLER_30_959 AVDD VSS sg13g2f_FILL8
XFILLER_30_967 AVDD VSS sg13g2f_FILL1
XFILLER_30_979 AVDD VSS sg13g2f_FILL8
XFILLER_30_987 AVDD VSS sg13g2f_FILL8
XFILLER_30_995 AVDD VSS sg13g2f_FILL8
XFILLER_30_1003 AVDD VSS sg13g2f_FILL4
XFILLER_30_1007 AVDD VSS sg13g2f_FILL1
XFILLER_30_1015 AVDD VSS sg13g2f_FILL8
XFILLER_30_1023 AVDD VSS sg13g2f_FILL8
XFILLER_30_1031 AVDD VSS sg13g2f_FILL8
XFILLER_30_1039 AVDD VSS sg13g2f_FILL8
XFILLER_30_1047 AVDD VSS sg13g2f_FILL8
XFILLER_30_1055 AVDD VSS sg13g2f_FILL8
XFILLER_30_1063 AVDD VSS sg13g2f_FILL8
XFILLER_30_1071 AVDD VSS sg13g2f_FILL8
XFILLER_30_1079 AVDD VSS sg13g2f_FILL8
XFILLER_30_1087 AVDD VSS sg13g2f_FILL8
XFILLER_30_1095 AVDD VSS sg13g2f_FILL8
XFILLER_30_1103 AVDD VSS sg13g2f_FILL8
XFILLER_30_1111 AVDD VSS sg13g2f_FILL8
XFILLER_30_1119 AVDD VSS sg13g2f_FILL1
XFILLER_30_1127 AVDD VSS sg13g2f_FILL8
XFILLER_30_1135 AVDD VSS sg13g2f_FILL8
XFILLER_30_1143 AVDD VSS sg13g2f_FILL8
XFILLER_30_1151 AVDD VSS sg13g2f_FILL8
XFILLER_30_1159 AVDD VSS sg13g2f_FILL8
XFILLER_30_1167 AVDD VSS sg13g2f_FILL8
XFILLER_30_1175 AVDD VSS sg13g2f_FILL8
XFILLER_30_1183 AVDD VSS sg13g2f_FILL8
XFILLER_30_1191 AVDD VSS sg13g2f_FILL8
XFILLER_30_1199 AVDD VSS sg13g2f_FILL8
XFILLER_30_1207 AVDD VSS sg13g2f_FILL8
XFILLER_30_1215 AVDD VSS sg13g2f_FILL8
XFILLER_30_1223 AVDD VSS sg13g2f_FILL8
XFILLER_30_1231 AVDD VSS sg13g2f_FILL1
XFILLER_30_1239 AVDD VSS sg13g2f_FILL8
XFILLER_30_1247 AVDD VSS sg13g2f_FILL8
XFILLER_30_1255 AVDD VSS sg13g2f_FILL8
XFILLER_30_1263 AVDD VSS sg13g2f_FILL4
XFILLER_30_1267 AVDD VSS sg13g2f_FILL1
XFILLER_30_1390 VDD VSS sg13g2f_FILL8
XFILLER_30_1398 VDD VSS sg13g2f_FILL8
XFILLER_30_1406 VDD VSS sg13g2f_FILL8
XFILLER_30_1414 VDD VSS sg13g2f_FILL8
XFILLER_30_1422 VDD VSS sg13g2f_FILL8
XFILLER_30_1430 VDD VSS sg13g2f_FILL8
XFILLER_30_1438 VDD VSS sg13g2f_FILL8
XFILLER_30_1446 VDD VSS sg13g2f_FILL8
XFILLER_30_1454 VDD VSS sg13g2f_FILL2
XFILLER_30_1547 VDD VSS sg13g2f_FILL4
XFILLER_31_1390 VDD VSS sg13g2f_FILL8
XFILLER_31_1398 VDD VSS sg13g2f_FILL8
XFILLER_31_1406 VDD VSS sg13g2f_FILL8
XFILLER_31_1414 VDD VSS sg13g2f_FILL8
XFILLER_31_1422 VDD VSS sg13g2f_FILL8
XFILLER_31_1430 VDD VSS sg13g2f_FILL8
XFILLER_31_1438 VDD VSS sg13g2f_FILL8
XFILLER_31_1446 VDD VSS sg13g2f_FILL8
XFILLER_31_1454 VDD VSS sg13g2f_FILL8
XFILLER_31_1462 VDD VSS sg13g2f_FILL8
XFILLER_31_1470 VDD VSS sg13g2f_FILL8
XFILLER_31_1478 VDD VSS sg13g2f_FILL8
XFILLER_31_1486 VDD VSS sg13g2f_FILL8
XFILLER_31_1494 VDD VSS sg13g2f_FILL8
XFILLER_31_1502 VDD VSS sg13g2f_FILL4
XFILLER_31_1517 VDD VSS sg13g2f_FILL8
XFILLER_31_1525 VDD VSS sg13g2f_FILL8
XFILLER_31_1533 VDD VSS sg13g2f_FILL8
XFILLER_31_1541 VDD VSS sg13g2f_FILL8
XFILLER_31_1549 VDD VSS sg13g2f_FILL2
XFILLER_32_1390 VDD VSS sg13g2f_FILL8
XFILLER_32_1398 VDD VSS sg13g2f_FILL8
XFILLER_32_1406 VDD VSS sg13g2f_FILL8
XFILLER_32_1414 VDD VSS sg13g2f_FILL8
XFILLER_32_1422 VDD VSS sg13g2f_FILL8
XFILLER_32_1430 VDD VSS sg13g2f_FILL8
XFILLER_32_1438 VDD VSS sg13g2f_FILL8
XFILLER_32_1446 VDD VSS sg13g2f_FILL8
XFILLER_32_1454 VDD VSS sg13g2f_FILL8
XFILLER_32_1462 VDD VSS sg13g2f_FILL8
XFILLER_32_1470 VDD VSS sg13g2f_FILL8
XFILLER_32_1478 VDD VSS sg13g2f_FILL8
XFILLER_32_1486 VDD VSS sg13g2f_FILL8
XFILLER_32_1494 VDD VSS sg13g2f_FILL4
XFILLER_32_1516 VDD VSS sg13g2f_FILL8
XFILLER_32_1524 VDD VSS sg13g2f_FILL8
XFILLER_32_1532 VDD VSS sg13g2f_FILL8
XFILLER_32_1540 VDD VSS sg13g2f_FILL8
XFILLER_32_1548 VDD VSS sg13g2f_FILL2
XFILLER_32_1550 VDD VSS sg13g2f_FILL1
XFILLER_33_1390 VDD VSS sg13g2f_FILL8
XFILLER_33_1398 VDD VSS sg13g2f_FILL8
XFILLER_33_1406 VDD VSS sg13g2f_FILL8
XFILLER_33_1414 VDD VSS sg13g2f_FILL8
XFILLER_33_1422 VDD VSS sg13g2f_FILL8
XFILLER_33_1430 VDD VSS sg13g2f_FILL8
XFILLER_33_1438 VDD VSS sg13g2f_FILL8
XFILLER_33_1446 VDD VSS sg13g2f_FILL8
XFILLER_33_1454 VDD VSS sg13g2f_FILL8
XFILLER_33_1462 VDD VSS sg13g2f_FILL8
XFILLER_33_1470 VDD VSS sg13g2f_FILL4
XFILLER_33_1474 VDD VSS sg13g2f_FILL1
XFILLER_33_1531 VDD VSS sg13g2f_FILL8
XFILLER_33_1539 VDD VSS sg13g2f_FILL8
XFILLER_33_1547 VDD VSS sg13g2f_FILL4
XFILLER_34_1390 VDD VSS sg13g2f_FILL8
XFILLER_34_1398 VDD VSS sg13g2f_FILL8
XFILLER_34_1406 VDD VSS sg13g2f_FILL8
XFILLER_34_1414 VDD VSS sg13g2f_FILL8
XFILLER_34_1422 VDD VSS sg13g2f_FILL8
XFILLER_34_1430 VDD VSS sg13g2f_FILL8
XFILLER_34_1438 VDD VSS sg13g2f_FILL8
XFILLER_34_1446 VDD VSS sg13g2f_FILL8
XFILLER_34_1454 VDD VSS sg13g2f_FILL8
XFILLER_34_1462 VDD VSS sg13g2f_FILL8
XFILLER_34_1470 VDD VSS sg13g2f_FILL8
XFILLER_34_1478 VDD VSS sg13g2f_FILL8
XFILLER_34_1486 VDD VSS sg13g2f_FILL8
XFILLER_34_1494 VDD VSS sg13g2f_FILL4
XFILLER_34_1505 VDD VSS sg13g2f_FILL4
XFILLER_34_1520 VDD VSS sg13g2f_FILL8
XFILLER_34_1528 VDD VSS sg13g2f_FILL8
XFILLER_34_1536 VDD VSS sg13g2f_FILL8
XFILLER_34_1544 VDD VSS sg13g2f_FILL4
XFILLER_34_1548 VDD VSS sg13g2f_FILL2
XFILLER_34_1550 VDD VSS sg13g2f_FILL1
XFILLER_35_1390 VDD VSS sg13g2f_FILL8
XFILLER_35_1398 VDD VSS sg13g2f_FILL8
XFILLER_35_1406 VDD VSS sg13g2f_FILL8
XFILLER_35_1414 VDD VSS sg13g2f_FILL8
XFILLER_35_1422 VDD VSS sg13g2f_FILL8
XFILLER_35_1430 VDD VSS sg13g2f_FILL8
XFILLER_35_1438 VDD VSS sg13g2f_FILL8
XFILLER_35_1446 VDD VSS sg13g2f_FILL8
XFILLER_35_1454 VDD VSS sg13g2f_FILL8
XFILLER_35_1462 VDD VSS sg13g2f_FILL8
XFILLER_35_1470 VDD VSS sg13g2f_FILL8
XFILLER_35_1478 VDD VSS sg13g2f_FILL8
XFILLER_35_1486 VDD VSS sg13g2f_FILL8
XFILLER_35_1536 VDD VSS sg13g2f_FILL8
XFILLER_35_1544 VDD VSS sg13g2f_FILL4
XFILLER_35_1548 VDD VSS sg13g2f_FILL2
XFILLER_35_1550 VDD VSS sg13g2f_FILL1
XFILLER_36_1390 VDD VSS sg13g2f_FILL8
XFILLER_36_1398 VDD VSS sg13g2f_FILL8
XFILLER_36_1406 VDD VSS sg13g2f_FILL8
XFILLER_36_1414 VDD VSS sg13g2f_FILL8
XFILLER_36_1422 VDD VSS sg13g2f_FILL8
XFILLER_36_1430 VDD VSS sg13g2f_FILL8
XFILLER_36_1438 VDD VSS sg13g2f_FILL8
XFILLER_36_1446 VDD VSS sg13g2f_FILL8
XFILLER_36_1454 VDD VSS sg13g2f_FILL8
XFILLER_36_1462 VDD VSS sg13g2f_FILL8
XFILLER_36_1470 VDD VSS sg13g2f_FILL8
XFILLER_36_1478 VDD VSS sg13g2f_FILL8
XFILLER_36_1486 VDD VSS sg13g2f_FILL8
XFILLER_36_1494 VDD VSS sg13g2f_FILL4
XFILLER_36_1505 VDD VSS sg13g2f_FILL4
XFILLER_36_1509 VDD VSS sg13g2f_FILL2
XFILLER_36_1511 VDD VSS sg13g2f_FILL1
XFILLER_36_1545 VDD VSS sg13g2f_FILL4
XFILLER_36_1549 VDD VSS sg13g2f_FILL2
XFILLER_37_1390 VDD VSS sg13g2f_FILL8
XFILLER_37_1398 VDD VSS sg13g2f_FILL8
XFILLER_37_1406 VDD VSS sg13g2f_FILL8
XFILLER_37_1414 VDD VSS sg13g2f_FILL8
XFILLER_37_1422 VDD VSS sg13g2f_FILL8
XFILLER_37_1430 VDD VSS sg13g2f_FILL8
XFILLER_37_1438 VDD VSS sg13g2f_FILL8
XFILLER_37_1446 VDD VSS sg13g2f_FILL8
XFILLER_37_1454 VDD VSS sg13g2f_FILL8
XFILLER_37_1462 VDD VSS sg13g2f_FILL8
XFILLER_37_1470 VDD VSS sg13g2f_FILL8
XFILLER_37_1478 VDD VSS sg13g2f_FILL8
XFILLER_37_1486 VDD VSS sg13g2f_FILL8
XFILLER_37_1494 VDD VSS sg13g2f_FILL8
XFILLER_37_1502 VDD VSS sg13g2f_FILL8
XFILLER_37_1510 VDD VSS sg13g2f_FILL4
XFILLER_37_1525 VDD VSS sg13g2f_FILL8
XFILLER_37_1533 VDD VSS sg13g2f_FILL8
XFILLER_37_1541 VDD VSS sg13g2f_FILL8
XFILLER_37_1549 VDD VSS sg13g2f_FILL2
XFILLER_38_1390 VDD VSS sg13g2f_FILL8
XFILLER_38_1398 VDD VSS sg13g2f_FILL8
XFILLER_38_1406 VDD VSS sg13g2f_FILL8
XFILLER_38_1414 VDD VSS sg13g2f_FILL8
XFILLER_38_1422 VDD VSS sg13g2f_FILL8
XFILLER_38_1430 VDD VSS sg13g2f_FILL8
XFILLER_38_1438 VDD VSS sg13g2f_FILL8
XFILLER_38_1446 VDD VSS sg13g2f_FILL8
XFILLER_38_1454 VDD VSS sg13g2f_FILL8
XFILLER_38_1462 VDD VSS sg13g2f_FILL8
XFILLER_38_1470 VDD VSS sg13g2f_FILL8
XFILLER_38_1478 VDD VSS sg13g2f_FILL8
XFILLER_38_1486 VDD VSS sg13g2f_FILL8
XFILLER_38_1494 VDD VSS sg13g2f_FILL4
XFILLER_38_1505 VDD VSS sg13g2f_FILL8
XFILLER_38_1513 VDD VSS sg13g2f_FILL1
XFILLER_38_1528 VDD VSS sg13g2f_FILL8
XFILLER_38_1536 VDD VSS sg13g2f_FILL8
XFILLER_38_1544 VDD VSS sg13g2f_FILL4
XFILLER_38_1548 VDD VSS sg13g2f_FILL2
XFILLER_38_1550 VDD VSS sg13g2f_FILL1
XFILLER_39_1390 VDD VSS sg13g2f_FILL8
XFILLER_39_1398 VDD VSS sg13g2f_FILL8
XFILLER_39_1406 VDD VSS sg13g2f_FILL8
XFILLER_39_1414 VDD VSS sg13g2f_FILL8
XFILLER_39_1422 VDD VSS sg13g2f_FILL8
XFILLER_39_1430 VDD VSS sg13g2f_FILL8
XFILLER_39_1438 VDD VSS sg13g2f_FILL8
XFILLER_39_1446 VDD VSS sg13g2f_FILL8
XFILLER_39_1454 VDD VSS sg13g2f_FILL8
XFILLER_39_1462 VDD VSS sg13g2f_FILL8
XFILLER_39_1470 VDD VSS sg13g2f_FILL8
XFILLER_39_1478 VDD VSS sg13g2f_FILL8
XFILLER_39_1486 VDD VSS sg13g2f_FILL8
XFILLER_39_1494 VDD VSS sg13g2f_FILL8
XFILLER_39_1502 VDD VSS sg13g2f_FILL8
XFILLER_39_1510 VDD VSS sg13g2f_FILL4
XFILLER_39_1514 VDD VSS sg13g2f_FILL1
XFILLER_39_1526 VDD VSS sg13g2f_FILL8
XFILLER_39_1534 VDD VSS sg13g2f_FILL8
XFILLER_39_1542 VDD VSS sg13g2f_FILL8
XFILLER_39_1550 VDD VSS sg13g2f_FILL1
XFILLER_40_1390 VDD VSS sg13g2f_FILL8
XFILLER_40_1398 VDD VSS sg13g2f_FILL8
XFILLER_40_1406 VDD VSS sg13g2f_FILL8
XFILLER_40_1414 VDD VSS sg13g2f_FILL8
XFILLER_40_1422 VDD VSS sg13g2f_FILL8
XFILLER_40_1430 VDD VSS sg13g2f_FILL8
XFILLER_40_1438 VDD VSS sg13g2f_FILL8
XFILLER_40_1446 VDD VSS sg13g2f_FILL8
XFILLER_40_1454 VDD VSS sg13g2f_FILL8
XFILLER_40_1462 VDD VSS sg13g2f_FILL8
XFILLER_40_1470 VDD VSS sg13g2f_FILL8
XFILLER_40_1478 VDD VSS sg13g2f_FILL8
XFILLER_40_1486 VDD VSS sg13g2f_FILL8
XFILLER_40_1494 VDD VSS sg13g2f_FILL4
XFILLER_40_1505 VDD VSS sg13g2f_FILL8
XFILLER_40_1513 VDD VSS sg13g2f_FILL4
XFILLER_40_1517 VDD VSS sg13g2f_FILL1
XFILLER_40_1529 VDD VSS sg13g2f_FILL8
XFILLER_40_1537 VDD VSS sg13g2f_FILL8
XFILLER_40_1545 VDD VSS sg13g2f_FILL4
XFILLER_40_1549 VDD VSS sg13g2f_FILL2
XFILLER_41_1390 VDD VSS sg13g2f_FILL8
XFILLER_41_1398 VDD VSS sg13g2f_FILL8
XFILLER_41_1406 VDD VSS sg13g2f_FILL8
XFILLER_41_1414 VDD VSS sg13g2f_FILL8
XFILLER_41_1422 VDD VSS sg13g2f_FILL8
XFILLER_41_1430 VDD VSS sg13g2f_FILL8
XFILLER_41_1438 VDD VSS sg13g2f_FILL8
XFILLER_41_1446 VDD VSS sg13g2f_FILL8
XFILLER_41_1454 VDD VSS sg13g2f_FILL8
XFILLER_41_1462 VDD VSS sg13g2f_FILL8
XFILLER_41_1470 VDD VSS sg13g2f_FILL8
XFILLER_41_1478 VDD VSS sg13g2f_FILL8
XFILLER_41_1486 VDD VSS sg13g2f_FILL8
XFILLER_41_1494 VDD VSS sg13g2f_FILL8
XFILLER_41_1502 VDD VSS sg13g2f_FILL8
XFILLER_41_1510 VDD VSS sg13g2f_FILL2
XFILLER_41_1512 VDD VSS sg13g2f_FILL1
XFILLER_41_1534 VDD VSS sg13g2f_FILL8
XFILLER_41_1542 VDD VSS sg13g2f_FILL8
XFILLER_41_1550 VDD VSS sg13g2f_FILL1
XFILLER_42_1390 VDD VSS sg13g2f_FILL8
XFILLER_42_1398 VDD VSS sg13g2f_FILL8
XFILLER_42_1406 VDD VSS sg13g2f_FILL8
XFILLER_42_1414 VDD VSS sg13g2f_FILL8
XFILLER_42_1422 VDD VSS sg13g2f_FILL8
XFILLER_42_1430 VDD VSS sg13g2f_FILL8
XFILLER_42_1438 VDD VSS sg13g2f_FILL8
XFILLER_42_1446 VDD VSS sg13g2f_FILL8
XFILLER_42_1454 VDD VSS sg13g2f_FILL8
XFILLER_42_1462 VDD VSS sg13g2f_FILL8
XFILLER_42_1470 VDD VSS sg13g2f_FILL8
XFILLER_42_1478 VDD VSS sg13g2f_FILL8
XFILLER_42_1486 VDD VSS sg13g2f_FILL8
XFILLER_42_1494 VDD VSS sg13g2f_FILL4
XFILLER_42_1505 VDD VSS sg13g2f_FILL8
XFILLER_42_1513 VDD VSS sg13g2f_FILL4
XFILLER_42_1531 VDD VSS sg13g2f_FILL8
XFILLER_42_1539 VDD VSS sg13g2f_FILL8
XFILLER_42_1547 VDD VSS sg13g2f_FILL4
XFILLER_43_1390 VDD VSS sg13g2f_FILL8
XFILLER_43_1398 VDD VSS sg13g2f_FILL8
XFILLER_43_1406 VDD VSS sg13g2f_FILL8
XFILLER_43_1414 VDD VSS sg13g2f_FILL8
XFILLER_43_1422 VDD VSS sg13g2f_FILL8
XFILLER_43_1430 VDD VSS sg13g2f_FILL8
XFILLER_43_1438 VDD VSS sg13g2f_FILL8
XFILLER_43_1446 VDD VSS sg13g2f_FILL8
XFILLER_43_1454 VDD VSS sg13g2f_FILL8
XFILLER_43_1462 VDD VSS sg13g2f_FILL8
XFILLER_43_1470 VDD VSS sg13g2f_FILL8
XFILLER_43_1478 VDD VSS sg13g2f_FILL8
XFILLER_43_1486 VDD VSS sg13g2f_FILL8
XFILLER_43_1494 VDD VSS sg13g2f_FILL8
XFILLER_43_1502 VDD VSS sg13g2f_FILL8
XFILLER_43_1510 VDD VSS sg13g2f_FILL8
XFILLER_43_1529 VDD VSS sg13g2f_FILL8
XFILLER_43_1537 VDD VSS sg13g2f_FILL8
XFILLER_43_1545 VDD VSS sg13g2f_FILL4
XFILLER_43_1549 VDD VSS sg13g2f_FILL2
XFILLER_44_1390 VDD VSS sg13g2f_FILL8
XFILLER_44_1398 VDD VSS sg13g2f_FILL8
XFILLER_44_1406 VDD VSS sg13g2f_FILL8
XFILLER_44_1414 VDD VSS sg13g2f_FILL8
XFILLER_44_1422 VDD VSS sg13g2f_FILL8
XFILLER_44_1430 VDD VSS sg13g2f_FILL8
XFILLER_44_1438 VDD VSS sg13g2f_FILL8
XFILLER_44_1446 VDD VSS sg13g2f_FILL8
XFILLER_44_1454 VDD VSS sg13g2f_FILL8
XFILLER_44_1462 VDD VSS sg13g2f_FILL8
XFILLER_44_1470 VDD VSS sg13g2f_FILL8
XFILLER_44_1478 VDD VSS sg13g2f_FILL8
XFILLER_44_1486 VDD VSS sg13g2f_FILL8
XFILLER_44_1494 VDD VSS sg13g2f_FILL4
XFILLER_44_1547 VDD VSS sg13g2f_FILL4
XFILLER_45_1390 VDD VSS sg13g2f_FILL8
XFILLER_45_1398 VDD VSS sg13g2f_FILL8
XFILLER_45_1406 VDD VSS sg13g2f_FILL8
XFILLER_45_1414 VDD VSS sg13g2f_FILL8
XFILLER_45_1422 VDD VSS sg13g2f_FILL8
XFILLER_45_1430 VDD VSS sg13g2f_FILL8
XFILLER_45_1438 VDD VSS sg13g2f_FILL8
XFILLER_45_1446 VDD VSS sg13g2f_FILL8
XFILLER_45_1454 VDD VSS sg13g2f_FILL8
XFILLER_45_1462 VDD VSS sg13g2f_FILL8
XFILLER_45_1470 VDD VSS sg13g2f_FILL8
XFILLER_45_1478 VDD VSS sg13g2f_FILL8
XFILLER_45_1486 VDD VSS sg13g2f_FILL8
XFILLER_45_1494 VDD VSS sg13g2f_FILL8
XFILLER_45_1502 VDD VSS sg13g2f_FILL8
XFILLER_45_1510 VDD VSS sg13g2f_FILL8
XFILLER_45_1529 VDD VSS sg13g2f_FILL8
XFILLER_45_1537 VDD VSS sg13g2f_FILL8
XFILLER_45_1545 VDD VSS sg13g2f_FILL4
XFILLER_45_1549 VDD VSS sg13g2f_FILL2
XFILLER_46_1390 VDD VSS sg13g2f_FILL8
XFILLER_46_1398 VDD VSS sg13g2f_FILL8
XFILLER_46_1406 VDD VSS sg13g2f_FILL8
XFILLER_46_1414 VDD VSS sg13g2f_FILL8
XFILLER_46_1422 VDD VSS sg13g2f_FILL8
XFILLER_46_1430 VDD VSS sg13g2f_FILL8
XFILLER_46_1438 VDD VSS sg13g2f_FILL8
XFILLER_46_1446 VDD VSS sg13g2f_FILL8
XFILLER_46_1454 VDD VSS sg13g2f_FILL8
XFILLER_46_1462 VDD VSS sg13g2f_FILL8
XFILLER_46_1470 VDD VSS sg13g2f_FILL8
XFILLER_46_1478 VDD VSS sg13g2f_FILL8
XFILLER_46_1486 VDD VSS sg13g2f_FILL8
XFILLER_46_1494 VDD VSS sg13g2f_FILL4
XFILLER_46_1505 VDD VSS sg13g2f_FILL8
XFILLER_46_1513 VDD VSS sg13g2f_FILL4
XFILLER_46_1517 VDD VSS sg13g2f_FILL1
XFILLER_46_1537 VDD VSS sg13g2f_FILL8
XFILLER_46_1545 VDD VSS sg13g2f_FILL4
XFILLER_46_1549 VDD VSS sg13g2f_FILL2
XFILLER_47_1390 VDD VSS sg13g2f_FILL8
XFILLER_47_1398 VDD VSS sg13g2f_FILL8
XFILLER_47_1406 VDD VSS sg13g2f_FILL8
XFILLER_47_1414 VDD VSS sg13g2f_FILL8
XFILLER_47_1422 VDD VSS sg13g2f_FILL8
XFILLER_47_1430 VDD VSS sg13g2f_FILL8
XFILLER_47_1438 VDD VSS sg13g2f_FILL8
XFILLER_47_1446 VDD VSS sg13g2f_FILL8
XFILLER_47_1454 VDD VSS sg13g2f_FILL8
XFILLER_47_1462 VDD VSS sg13g2f_FILL8
XFILLER_47_1470 VDD VSS sg13g2f_FILL8
XFILLER_47_1478 VDD VSS sg13g2f_FILL8
XFILLER_47_1486 VDD VSS sg13g2f_FILL8
XFILLER_47_1494 VDD VSS sg13g2f_FILL8
XFILLER_47_1502 VDD VSS sg13g2f_FILL4
XFILLER_47_1506 VDD VSS sg13g2f_FILL1
XFILLER_47_1534 VDD VSS sg13g2f_FILL8
XFILLER_47_1542 VDD VSS sg13g2f_FILL8
XFILLER_47_1550 VDD VSS sg13g2f_FILL1
XFILLER_48_1390 VDD VSS sg13g2f_FILL8
XFILLER_48_1398 VDD VSS sg13g2f_FILL8
XFILLER_48_1406 VDD VSS sg13g2f_FILL8
XFILLER_48_1414 VDD VSS sg13g2f_FILL8
XFILLER_48_1422 VDD VSS sg13g2f_FILL8
XFILLER_48_1430 VDD VSS sg13g2f_FILL8
XFILLER_48_1438 VDD VSS sg13g2f_FILL8
XFILLER_48_1446 VDD VSS sg13g2f_FILL8
XFILLER_48_1454 VDD VSS sg13g2f_FILL8
XFILLER_48_1462 VDD VSS sg13g2f_FILL8
XFILLER_48_1470 VDD VSS sg13g2f_FILL8
XFILLER_48_1478 VDD VSS sg13g2f_FILL8
XFILLER_48_1486 VDD VSS sg13g2f_FILL8
XFILLER_48_1494 VDD VSS sg13g2f_FILL4
XFILLER_48_1505 VDD VSS sg13g2f_FILL8
XFILLER_48_1513 VDD VSS sg13g2f_FILL4
XFILLER_48_1517 VDD VSS sg13g2f_FILL1
XFILLER_48_1529 VDD VSS sg13g2f_FILL8
XFILLER_48_1537 VDD VSS sg13g2f_FILL8
XFILLER_48_1545 VDD VSS sg13g2f_FILL4
XFILLER_48_1549 VDD VSS sg13g2f_FILL2
XFILLER_49_1390 VDD VSS sg13g2f_FILL8
XFILLER_49_1398 VDD VSS sg13g2f_FILL8
XFILLER_49_1406 VDD VSS sg13g2f_FILL8
XFILLER_49_1414 VDD VSS sg13g2f_FILL8
XFILLER_49_1422 VDD VSS sg13g2f_FILL8
XFILLER_49_1430 VDD VSS sg13g2f_FILL8
XFILLER_49_1438 VDD VSS sg13g2f_FILL8
XFILLER_49_1446 VDD VSS sg13g2f_FILL8
XFILLER_49_1454 VDD VSS sg13g2f_FILL8
XFILLER_49_1462 VDD VSS sg13g2f_FILL8
XFILLER_49_1470 VDD VSS sg13g2f_FILL8
XFILLER_49_1478 VDD VSS sg13g2f_FILL8
XFILLER_49_1486 VDD VSS sg13g2f_FILL8
XFILLER_49_1494 VDD VSS sg13g2f_FILL8
XFILLER_49_1502 VDD VSS sg13g2f_FILL8
XFILLER_49_1510 VDD VSS sg13g2f_FILL8
XFILLER_49_1518 VDD VSS sg13g2f_FILL8
XFILLER_49_1526 VDD VSS sg13g2f_FILL8
XFILLER_49_1534 VDD VSS sg13g2f_FILL8
XFILLER_49_1542 VDD VSS sg13g2f_FILL8
XFILLER_49_1550 VDD VSS sg13g2f_FILL1
XFILLER_50_1390 VDD VSS sg13g2f_FILL8
XFILLER_50_1398 VDD VSS sg13g2f_FILL8
XFILLER_50_1406 VDD VSS sg13g2f_FILL8
XFILLER_50_1414 VDD VSS sg13g2f_FILL8
XFILLER_50_1422 VDD VSS sg13g2f_FILL8
XFILLER_50_1430 VDD VSS sg13g2f_FILL8
XFILLER_50_1438 VDD VSS sg13g2f_FILL8
XFILLER_50_1446 VDD VSS sg13g2f_FILL8
XFILLER_50_1454 VDD VSS sg13g2f_FILL8
XFILLER_50_1462 VDD VSS sg13g2f_FILL8
XFILLER_50_1470 VDD VSS sg13g2f_FILL8
XFILLER_50_1478 VDD VSS sg13g2f_FILL8
XFILLER_50_1486 VDD VSS sg13g2f_FILL8
XFILLER_50_1494 VDD VSS sg13g2f_FILL4
XFILLER_50_1505 VDD VSS sg13g2f_FILL8
XFILLER_50_1513 VDD VSS sg13g2f_FILL8
XFILLER_50_1521 VDD VSS sg13g2f_FILL8
XFILLER_50_1529 VDD VSS sg13g2f_FILL8
XFILLER_50_1537 VDD VSS sg13g2f_FILL8
XFILLER_50_1545 VDD VSS sg13g2f_FILL4
XFILLER_50_1549 VDD VSS sg13g2f_FILL2
XFILLER_51_1390 VDD VSS sg13g2f_FILL8
XFILLER_51_1398 VDD VSS sg13g2f_FILL8
XFILLER_51_1406 VDD VSS sg13g2f_FILL8
XFILLER_51_1414 VDD VSS sg13g2f_FILL8
XFILLER_51_1422 VDD VSS sg13g2f_FILL8
XFILLER_51_1430 VDD VSS sg13g2f_FILL8
XFILLER_51_1438 VDD VSS sg13g2f_FILL8
XFILLER_51_1446 VDD VSS sg13g2f_FILL8
XFILLER_51_1454 VDD VSS sg13g2f_FILL8
XFILLER_51_1462 VDD VSS sg13g2f_FILL8
XFILLER_51_1470 VDD VSS sg13g2f_FILL8
XFILLER_51_1478 VDD VSS sg13g2f_FILL8
XFILLER_51_1486 VDD VSS sg13g2f_FILL8
XFILLER_51_1494 VDD VSS sg13g2f_FILL8
XFILLER_51_1502 VDD VSS sg13g2f_FILL8
XFILLER_51_1533 VDD VSS sg13g2f_FILL8
XFILLER_51_1541 VDD VSS sg13g2f_FILL8
XFILLER_51_1549 VDD VSS sg13g2f_FILL2
XFILLER_52_1390 VDD VSS sg13g2f_FILL8
XFILLER_52_1398 VDD VSS sg13g2f_FILL8
XFILLER_52_1406 VDD VSS sg13g2f_FILL8
XFILLER_52_1414 VDD VSS sg13g2f_FILL8
XFILLER_52_1422 VDD VSS sg13g2f_FILL8
XFILLER_52_1430 VDD VSS sg13g2f_FILL8
XFILLER_52_1438 VDD VSS sg13g2f_FILL8
XFILLER_52_1446 VDD VSS sg13g2f_FILL8
XFILLER_52_1454 VDD VSS sg13g2f_FILL8
XFILLER_52_1462 VDD VSS sg13g2f_FILL8
XFILLER_52_1470 VDD VSS sg13g2f_FILL8
XFILLER_52_1478 VDD VSS sg13g2f_FILL8
XFILLER_52_1486 VDD VSS sg13g2f_FILL8
XFILLER_52_1494 VDD VSS sg13g2f_FILL1
XFILLER_52_1502 VDD VSS sg13g2f_FILL8
XFILLER_52_1510 VDD VSS sg13g2f_FILL8
XFILLER_52_1518 VDD VSS sg13g2f_FILL8
XFILLER_52_1526 VDD VSS sg13g2f_FILL8
XFILLER_52_1534 VDD VSS sg13g2f_FILL8
XFILLER_52_1542 VDD VSS sg13g2f_FILL8
XFILLER_52_1550 VDD VSS sg13g2f_FILL1
.ENDS SARADC
* CDL Netlist generated by OpenROAD

*.BUSDELIMITER [

.SUBCKT SPI CEB CLK DATA DOUT_DAT DOUT_EN RD[0] RD[10] RD[11]
+ RD[12] RD[13] RD[14] RD[15] RD[16] RD[17] RD[18] RD[19] RD[1]
+ RD[20] RD[21] RD[22] RD[23] RD[24] RD[25] RD[26] RD[27] RD[28]
+ RD[29] RD[2] RD[30] RD[31] RD[32] RD[33] RD[34] RD[35] RD[36]
+ RD[37] RD[38] RD[39] RD[3] RD[40] RD[41] RD[42] RD[43] RD[44]
+ RD[45] RD[46] RD[47] RD[4] RD[5] RD[6] RD[7] RD[8] RD[9] RST
+ R[0] R[10] R[11] R[12] R[13] R[14] R[15] R[16] R[17] R[18]
+ R[19] R[1] R[20] R[21] R[22] R[23] R[24] R[25] R[26] R[27]
+ R[28] R[29] R[2] R[30] R[31] R[32] R[33] R[34] R[35] R[36]
+ R[37] R[38] R[39] R[3] R[40] R[41] R[42] R[43] R[44] R[45]
+ R[46] R[47] R[48] R[49] R[4] R[50] R[51] R[52] R[53] R[54]
+ R[55] R[56] R[57] R[58] R[59] R[5] R[60] R[61] R[62] R[63]
+ R[6] R[7] R[8] R[9] VSS VDD
Xins_223_ R[42] raddr\[2\] ins_124_ VDD VSS ins_036_ sg13g2_MUX2D1
Xins_224_ R[43] sft_reg\[3\] ins_124_ VDD VSS ins_037_ sg13g2_MUX2D1
Xins_225_ R[44] sft_reg\[4\] ins_124_ VDD VSS ins_038_ sg13g2_MUX2D1
Xins_226_ R[45] sft_reg\[5\] ins_124_ VDD VSS ins_039_ sg13g2_MUX2D1
Xins_227_ R[46] sft_reg\[6\] ins_124_ VDD VSS ins_040_ sg13g2_MUX2D1
Xins_228_ R[47] sft_reg\[7\] ins_124_ VDD VSS ins_041_ sg13g2_MUX2D1
Xins_229_ addr\[0\] addr\[1\] VDD VSS ins_125_ sg13g2_NR2D1
Xins_230_ ins_110_ ins_125_ VDD VSS ins_126_ sg13g2_AN2D1
Xins_231_ ins_121_ ins_126_ VDD VSS ins_127_ sg13g2_AN2D1
Xins_232_ R[0] raddr\[0\] ins_127_ VDD VSS ins_042_ sg13g2_MUX2D1
Xins_233_ R[1] raddr\[1\] ins_127_ VDD VSS ins_043_ sg13g2_MUX2D1
Xins_234_ R[2] raddr\[2\] ins_127_ VDD VSS ins_044_ sg13g2_MUX2D1
Xins_235_ R[3] sft_reg\[3\] ins_127_ VDD VSS ins_045_ sg13g2_MUX2D1
Xins_236_ R[4] sft_reg\[4\] ins_127_ VDD VSS ins_046_ sg13g2_MUX2D1
Xins_237_ R[5] sft_reg\[5\] ins_127_ VDD VSS ins_047_ sg13g2_MUX2D1
Xins_238_ R[6] sft_reg\[6\] ins_127_ VDD VSS ins_048_ sg13g2_MUX2D1
Xins_239_ R[7] sft_reg\[7\] ins_127_ VDD VSS ins_049_ sg13g2_MUX2D1
Xins_240_ ins_108_ addr\[1\] ins_110_ VDD VSS ins_128_ sg13g2_ND3D1
Xins_241_ ins_122_ ins_128_ VDD VSS ins_129_ sg13g2_NR2D1
Xins_242_ R[16] raddr\[0\] ins_129_ VDD VSS ins_050_ sg13g2_MUX2D1
Xins_243_ R[17] raddr\[1\] ins_129_ VDD VSS ins_051_ sg13g2_MUX2D1
Xins_244_ R[18] raddr\[2\] ins_129_ VDD VSS ins_052_ sg13g2_MUX2D1
Xins_245_ R[19] sft_reg\[3\] ins_129_ VDD VSS ins_053_ sg13g2_MUX2D1
Xins_246_ R[20] sft_reg\[4\] ins_129_ VDD VSS ins_054_ sg13g2_MUX2D1
Xins_247_ R[21] sft_reg\[5\] ins_129_ VDD VSS ins_055_ sg13g2_MUX2D1
Xins_248_ R[22] sft_reg\[6\] ins_129_ VDD VSS ins_056_ sg13g2_MUX2D1
Xins_249_ R[23] sft_reg\[7\] ins_129_ VDD VSS ins_057_ sg13g2_MUX2D1
Xins_250_ addr\[0\] addr\[1\] VDD VSS ins_130_ sg13g2_AN2D1
Xins_251_ addr\[2\] ins_121_ ins_130_ VDD VSS ins_131_ sg13g2_ND3D1
Xins_252_ raddr\[0\] R[56] ins_131_ VDD VSS ins_058_ sg13g2_MUX2D1
Xins_253_ raddr\[1\] R[57] ins_131_ VDD VSS ins_059_ sg13g2_MUX2D1
Xins_254_ raddr\[2\] R[58] ins_131_ VDD VSS ins_060_ sg13g2_MUX2D1
Xins_255_ sft_reg\[3\] R[59] ins_131_ VDD VSS ins_061_ sg13g2_MUX2D1
Xins_256_ sft_reg\[4\] R[60] ins_131_ VDD VSS ins_062_ sg13g2_MUX2D1
Xins_257_ sft_reg\[5\] R[61] ins_131_ VDD VSS ins_063_ sg13g2_MUX2D1
Xins_258_ sft_reg\[6\] R[62] ins_131_ VDD VSS ins_064_ sg13g2_MUX2D1
Xins_259_ sft_reg\[7\] R[63] ins_131_ VDD VSS ins_065_ sg13g2_MUX2D1
Xins_260_ genblk1.counter\[18\] genblk1.counter\[19\] VDD
+ VSS ins_132_ sg13g2_NR2D1
Xins_261_ genblk1.counter\[17\] genblk1.counter\[20\] VDD
+ VSS ins_133_ sg13g2_NR2D1
Xins_262_ genblk1.counter\[14\] genblk1.counter\[15\] VDD
+ VSS ins_134_ sg13g2_NR2D1
Xins_263_ genblk1.counter\[13\] genblk1.counter\[16\] VDD
+ VSS ins_135_ sg13g2_NR2D1
Xins_264_ ins_132_ ins_133_ ins_134_ ins_135_ VDD VSS ins_136_
+ sg13g2_ND4D1
Xins_265_ re ins_136_ VDD VSS ins_137_ sg13g2_ND2D1
Xins_266_ ins_137_ eno VSS VDD sg13g2_INVD1
Xins_267_ addr\[0\] ins_109_ ins_110_ VDD VSS ins_138_ sg13g2_ND3D1
Xins_268_ addr\[0\] ins_109_ ins_110_ RD[8] VDD VSS ins_139_
+ sg13g2_ND4D1
Xins_269_ ins_110_ RD[0] ins_125_ VDD VSS ins_140_ sg13g2_ND3D1
Xins_270_ addr\[2\] RD[32] ins_125_ VDD VSS ins_141_ sg13g2_ND3D1
Xins_271_ addr\[0\] ins_109_ addr\[2\] RD[40] VDD VSS ins_142_
+ sg13g2_ND4D1
Xins_272_ ins_108_ addr\[1\] ins_110_ RD[16] VDD VSS ins_143_
+ sg13g2_ND4D1
Xins_273_ ins_110_ ins_130_ VDD VSS ins_144_ sg13g2_AN2D1
Xins_274_ ins_110_ RD[24] ins_130_ VDD VSS ins_145_ sg13g2_ND3D1
Xins_275_ ins_139_ ins_140_ ins_143_ ins_145_ VDD VSS ins_146_
+ sg13g2_ND4D1
Xins_276_ encap ins_141_ ins_142_ VDD VSS ins_147_ sg13g2_ND3D1
Xins_277_ bus_cap\[0\] ins_137_ encap VDD VSS ins_148_ sg13g2_AO21D1
Xins_278_ ins_146_ ins_147_ ins_148_ VDD VSS ins_066_ sg13g2_OA21D1
Xins_279_ bus_cap\[0\] bus_cap\[1\] ins_137_ VDD VSS ins_149_
+ sg13g2_MUX2D1
Xins_280_ ins_108_ addr\[1\] ins_110_ RD[17] VDD VSS ins_150_
+ sg13g2_ND4D1
Xins_281_ ins_110_ RD[1] ins_125_ VDD VSS ins_151_ sg13g2_ND3D1
Xins_282_ ins_150_ ins_151_ VDD VSS ins_152_ sg13g2_AN2D1
Xins_283_ addr\[2\] RD[33] ins_125_ VDD VSS ins_153_ sg13g2_ND3D1
Xins_284_ addr\[0\] ins_109_ ins_110_ RD[9] VDD VSS ins_154_
+ sg13g2_ND4D1
Xins_285_ ins_153_ ins_154_ VDD VSS ins_155_ sg13g2_AN2D1
Xins_286_ addr\[0\] ins_109_ addr\[2\] RD[41] VDD VSS ins_156_
+ sg13g2_ND4D1
Xins_287_ ins_110_ RD[25] ins_130_ VDD VSS ins_157_ sg13g2_ND3D1
Xins_288_ ins_152_ ins_155_ ins_156_ ins_157_ VDD VSS ins_158_
+ sg13g2_ND4D1
Xins_289_ ins_149_ ins_158_ encap VDD VSS ins_067_ sg13g2_MUX2D1
Xins_290_ bus_cap\[1\] bus_cap\[2\] ins_137_ VDD VSS ins_159_
+ sg13g2_MUX2D1
Xins_291_ addr\[2\] RD[34] ins_125_ VDD VSS ins_160_ sg13g2_ND3D1
Xins_292_ addr\[0\] ins_109_ ins_110_ RD[10] VDD VSS ins_161_
+ sg13g2_ND4D1
Xins_293_ ins_160_ ins_161_ VDD VSS ins_162_ sg13g2_ND2D1
Xins_294_ ins_110_ RD[26] ins_130_ VDD VSS ins_163_ sg13g2_ND3D1
Xins_295_ ins_108_ addr\[1\] ins_110_ RD[18] VDD VSS ins_164_
+ sg13g2_ND4D1
Xins_296_ ins_110_ RD[2] ins_125_ VDD VSS ins_165_ sg13g2_ND3D1
Xins_297_ addr\[0\] ins_109_ addr\[2\] RD[42] VDD VSS ins_166_
+ sg13g2_ND4D1
Xins_298_ ins_163_ ins_164_ ins_165_ ins_166_ VDD VSS ins_167_
+ sg13g2_ND4D1
Xins_299_ ins_162_ ins_167_ VDD VSS ins_168_ sg13g2_OR2D1
Xins_300_ ins_159_ ins_168_ encap VDD VSS ins_068_ sg13g2_MUX2D1
Xins_301_ bus_cap\[2\] bus_cap\[3\] ins_137_ VDD VSS ins_169_
+ sg13g2_MUX2D1
Xins_302_ addr\[0\] ins_109_ ins_110_ RD[11] VDD VSS ins_170_
+ sg13g2_ND4D1
Xins_303_ ins_110_ RD[27] ins_130_ VDD VSS ins_171_ sg13g2_ND3D1
Xins_304_ ins_170_ ins_171_ VDD VSS ins_172_ sg13g2_ND2D1
Xins_305_ ins_110_ RD[3] ins_125_ VDD VSS ins_173_ sg13g2_ND3D1
Xins_306_ ins_108_ addr\[1\] ins_110_ RD[19] VDD VSS ins_174_
+ sg13g2_ND4D1
Xins_307_ addr\[2\] RD[35] ins_125_ VDD VSS ins_175_ sg13g2_ND3D1
Xins_308_ addr\[0\] ins_109_ addr\[2\] RD[43] VDD VSS ins_176_
+ sg13g2_ND4D1
Xins_309_ ins_173_ ins_174_ ins_175_ ins_176_ VDD VSS ins_177_
+ sg13g2_ND4D1
Xins_310_ ins_172_ ins_177_ VDD VSS ins_178_ sg13g2_OR2D1
Xins_311_ ins_169_ ins_178_ encap VDD VSS ins_069_ sg13g2_MUX2D1
Xins_312_ bus_cap\[3\] bus_cap\[4\] ins_137_ VDD VSS ins_179_
+ sg13g2_MUX2D1
Xins_313_ addr\[0\] ins_109_ ins_110_ RD[12] VDD VSS ins_180_
+ sg13g2_ND4D1
Xins_314_ ins_108_ addr\[1\] ins_110_ RD[20] VDD VSS ins_181_
+ sg13g2_ND4D1
Xins_315_ ins_180_ ins_181_ VDD VSS ins_182_ sg13g2_ND2D1
Xins_316_ ins_110_ RD[4] ins_125_ VDD VSS ins_183_ sg13g2_ND3D1
Xins_317_ ins_110_ RD[28] ins_130_ VDD VSS ins_184_ sg13g2_ND3D1
Xins_318_ addr\[2\] RD[36] ins_125_ VDD VSS ins_185_ sg13g2_ND3D1
Xins_319_ addr\[0\] ins_109_ addr\[2\] RD[44] VDD VSS ins_186_
+ sg13g2_ND4D1
Xins_320_ ins_183_ ins_184_ ins_185_ ins_186_ VDD VSS ins_187_
+ sg13g2_ND4D1
Xins_321_ ins_182_ ins_187_ VDD VSS ins_188_ sg13g2_OR2D1
Xins_322_ ins_179_ ins_188_ encap VDD VSS ins_070_ sg13g2_MUX2D1
Xins_323_ bus_cap\[4\] bus_cap\[5\] ins_137_ VDD VSS ins_189_
+ sg13g2_MUX2D1
Xins_324_ addr\[0\] ins_109_ ins_110_ RD[13] VDD VSS ins_190_
+ sg13g2_ND4D1
Xins_325_ ins_110_ RD[29] ins_130_ VDD VSS ins_191_ sg13g2_ND3D1
Xins_326_ ins_190_ ins_191_ VDD VSS ins_192_ sg13g2_ND2D1
Xins_327_ ins_110_ RD[5] ins_125_ VDD VSS ins_193_ sg13g2_ND3D1
Xins_328_ ins_108_ addr\[1\] ins_110_ RD[21] VDD VSS ins_194_
+ sg13g2_ND4D1
Xins_329_ addr\[2\] RD[37] ins_125_ VDD VSS ins_195_ sg13g2_ND3D1
Xins_330_ addr\[0\] ins_109_ addr\[2\] RD[45] VDD VSS ins_196_
+ sg13g2_ND4D1
Xins_331_ ins_193_ ins_194_ ins_195_ ins_196_ VDD VSS ins_197_
+ sg13g2_ND4D1
Xins_332_ ins_192_ ins_197_ VDD VSS ins_198_ sg13g2_OR2D1
Xins_333_ ins_189_ ins_198_ encap VDD VSS ins_071_ sg13g2_MUX2D1
Xins_334_ bus_cap\[5\] bus_cap\[6\] ins_137_ VDD VSS ins_199_
+ sg13g2_MUX2D1
Xins_335_ ins_110_ RD[6] ins_125_ VDD VSS ins_200_ sg13g2_ND3D1
Xins_336_ ins_108_ addr\[1\] ins_110_ RD[22] VDD VSS ins_201_
+ sg13g2_ND4D1
Xins_337_ ins_200_ ins_201_ VDD VSS ins_202_ sg13g2_AN2D1
Xins_338_ addr\[0\] ins_109_ addr\[2\] RD[46] VDD VSS ins_203_
+ sg13g2_ND4D1
Xins_339_ ins_110_ RD[30] ins_130_ VDD VSS ins_204_ sg13g2_ND3D1
Xins_340_ addr\[2\] RD[38] ins_125_ VDD VSS ins_205_ sg13g2_ND3D1
Xins_341_ addr\[0\] ins_109_ ins_110_ RD[14] VDD VSS ins_206_
+ sg13g2_ND4D1
Xins_342_ ins_205_ ins_206_ VDD VSS ins_207_ sg13g2_AN2D1
Xins_343_ ins_202_ ins_203_ ins_204_ ins_207_ VDD VSS ins_208_
+ sg13g2_ND4D1
Xins_344_ ins_199_ ins_208_ encap VDD VSS ins_072_ sg13g2_MUX2D1
Xins_345_ bus_cap\[6\] bus_cap\[7\] ins_137_ VDD VSS ins_209_
+ sg13g2_MUX2D1
Xins_346_ addr\[2\] RD[39] ins_125_ VDD VSS ins_210_ sg13g2_ND3D1
Xins_347_ addr\[0\] ins_109_ ins_110_ RD[15] VDD VSS ins_211_
+ sg13g2_ND4D1
Xins_348_ ins_108_ addr\[1\] ins_110_ RD[23] VDD VSS ins_212_
+ sg13g2_ND4D1
Xins_349_ ins_110_ RD[7] ins_125_ VDD VSS ins_213_ sg13g2_ND3D1
Xins_350_ ins_212_ ins_213_ VDD VSS ins_214_ sg13g2_AN2D1
Xins_351_ ins_110_ RD[31] ins_130_ VDD VSS ins_215_ sg13g2_ND3D1
Xins_352_ addr\[0\] ins_109_ addr\[2\] RD[47] VDD VSS ins_216_
+ sg13g2_ND4D1
Xins_353_ ins_211_ ins_216_ VDD VSS ins_217_ sg13g2_AN2D1
Xins_354_ ins_210_ ins_214_ ins_215_ ins_217_ VDD VSS ins_218_
+ sg13g2_ND4D1
Xins_355_ ins_209_ ins_218_ encap VDD VSS ins_073_ sg13g2_MUX2D1
Xins_356_ ins_108_ addr\[1\] addr\[2\] ins_121_ VDD VSS ins_219_
+ sg13g2_ND4D1
Xins_357_ raddr\[0\] R[48] ins_219_ VDD VSS ins_074_ sg13g2_MUX2D1
Xins_358_ raddr\[1\] R[49] ins_219_ VDD VSS ins_075_ sg13g2_MUX2D1
Xins_359_ raddr\[2\] R[50] ins_219_ VDD VSS ins_076_ sg13g2_MUX2D1
Xins_360_ sft_reg\[3\] R[51] ins_219_ VDD VSS ins_077_ sg13g2_MUX2D1
Xins_361_ sft_reg\[4\] R[52] ins_219_ VDD VSS ins_078_ sg13g2_MUX2D1
Xins_362_ sft_reg\[5\] R[53] ins_219_ VDD VSS ins_079_ sg13g2_MUX2D1
Xins_363_ sft_reg\[6\] R[54] ins_219_ VDD VSS ins_080_ sg13g2_MUX2D1
Xins_364_ sft_reg\[7\] R[55] ins_219_ VDD VSS ins_081_ sg13g2_MUX2D1
Xins_365_ CEB ins_021_ VDD VSS ins_011_ sg13g2_NR2D1
Xins_366_ we DATA ins_011_ VDD VSS ins_082_ sg13g2_MUX2D1
Xins_367_ addr\[2\] ins_121_ ins_125_ VDD VSS ins_220_ sg13g2_ND3D1
Xins_368_ raddr\[0\] R[32] ins_220_ VDD VSS ins_083_ sg13g2_MUX2D1
Xins_369_ raddr\[1\] R[33] ins_220_ VDD VSS ins_084_ sg13g2_MUX2D1
Xins_370_ raddr\[2\] R[34] ins_220_ VDD VSS ins_085_ sg13g2_MUX2D1
Xins_371_ sft_reg\[3\] R[35] ins_220_ VDD VSS ins_086_ sg13g2_MUX2D1
Xins_372_ sft_reg\[4\] R[36] ins_220_ VDD VSS ins_087_ sg13g2_MUX2D1
Xins_373_ sft_reg\[5\] R[37] ins_220_ VDD VSS ins_088_ sg13g2_MUX2D1
Xins_374_ sft_reg\[6\] R[38] ins_220_ VDD VSS ins_089_ sg13g2_MUX2D1
Xins_375_ sft_reg\[7\] R[39] ins_220_ VDD VSS ins_090_ sg13g2_MUX2D1
Xins_376_ ins_121_ ins_144_ VDD VSS ins_221_ sg13g2_AN2D1
Xins_377_ R[24] raddr\[0\] ins_221_ VDD VSS ins_091_ sg13g2_MUX2D1
Xins_378_ R[25] raddr\[1\] ins_221_ VDD VSS ins_092_ sg13g2_MUX2D1
Xins_379_ R[26] raddr\[2\] ins_221_ VDD VSS ins_093_ sg13g2_MUX2D1
Xins_380_ R[27] sft_reg\[3\] ins_221_ VDD VSS ins_094_ sg13g2_MUX2D1
Xins_381_ R[28] sft_reg\[4\] ins_221_ VDD VSS ins_095_ sg13g2_MUX2D1
Xins_382_ R[29] sft_reg\[5\] ins_221_ VDD VSS ins_096_ sg13g2_MUX2D1
Xins_383_ R[30] sft_reg\[6\] ins_221_ VDD VSS ins_097_ sg13g2_MUX2D1
Xins_384_ R[31] sft_reg\[7\] ins_221_ VDD VSS ins_098_ sg13g2_MUX2D1
Xins_385_ ins_122_ ins_138_ VDD VSS ins_222_ sg13g2_NR2D1
Xins_386_ R[8] raddr\[0\] ins_222_ VDD VSS ins_099_ sg13g2_MUX2D1
Xins_387_ R[9] raddr\[1\] ins_222_ VDD VSS ins_100_ sg13g2_MUX2D1
Xins_388_ R[10] raddr\[2\] ins_222_ VDD VSS ins_101_ sg13g2_MUX2D1
Xins_389_ R[11] sft_reg\[3\] ins_222_ VDD VSS ins_102_ sg13g2_MUX2D1
Xins_390_ R[12] sft_reg\[4\] ins_222_ VDD VSS ins_103_ sg13g2_MUX2D1
Xins_391_ R[13] sft_reg\[5\] ins_222_ VDD VSS ins_104_ sg13g2_MUX2D1
Xins_392_ R[14] sft_reg\[6\] ins_222_ VDD VSS ins_105_ sg13g2_MUX2D1
Xins_393_ R[15] sft_reg\[7\] ins_222_ VDD VSS ins_106_ sg13g2_MUX2D1
Xins_394_ ins_022_ genblk1.counter\[1\] VDD VSS ins_013_ sg13g2_AN2D1
Xins_395_ re DATA ins_013_ VDD VSS ins_107_ sg13g2_MUX2D1
Xins_396_ ins_022_ genblk1.counter\[2\] VDD VSS ins_014_ sg13g2_AN2D1
Xins_397_ ins_022_ genblk1.counter\[3\] VDD VSS ins_015_ sg13g2_AN2D1
Xins_398_ ins_022_ genblk1.counter\[4\] VDD VSS ins_016_ sg13g2_AN2D1
Xins_399_ ins_022_ encap VDD VSS ins_017_ sg13g2_AN2D1
Xins_400_ ins_022_ genblk1.counter\[6\] VDD VSS ins_018_ sg13g2_AN2D1
Xins_401_ ins_022_ genblk1.counter\[7\] VDD VSS ins_019_ sg13g2_AN2D1
Xins_402_ ins_022_ genblk1.counter\[8\] VDD VSS ins_020_ sg13g2_AN2D1
Xins_403_ ins_022_ genblk1.counter\[9\] VDD VSS ins_001_ sg13g2_AN2D1
Xins_404_ ins_022_ genblk1.counter\[10\] VDD VSS ins_002_
+ sg13g2_AN2D1
Xins_405_ ins_022_ genblk1.counter\[11\] VDD VSS ins_003_
+ sg13g2_AN2D1
Xins_406_ ins_022_ genblk1.counter\[12\] VDD VSS ins_004_
+ sg13g2_AN2D1
Xins_407_ ins_022_ genblk1.counter\[13\] VDD VSS ins_005_
+ sg13g2_AN2D1
Xins_408_ ins_022_ genblk1.counter\[14\] VDD VSS ins_006_
+ sg13g2_AN2D1
Xins_409_ ins_022_ genblk1.counter\[15\] VDD VSS ins_007_
+ sg13g2_AN2D1
Xins_410_ ins_022_ genblk1.counter\[16\] VDD VSS ins_008_
+ sg13g2_AN2D1
Xins_411_ ins_022_ genblk1.counter\[17\] VDD VSS ins_009_
+ sg13g2_AN2D1
Xins_412_ ins_022_ genblk1.counter\[18\] VDD VSS ins_010_
+ sg13g2_AN2D1
Xins_413_ ins_022_ genblk1.counter\[19\] VDD VSS ins_012_
+ sg13g2_AN2D1
Xins_414_ bus_cap\[7\] eno VDD VSS ins_000_ sg13g2_AN2D1
Xins_415_ ins_022_ enoz VDD VSS DOUT_EN sg13g2_AN2D1
Xins_416_ CEB ins_022_ VSS VDD sg13g2_INVD1
Xins_417_ addr\[0\] ins_108_ VSS VDD sg13g2_INVD1
Xins_418_ addr\[1\] ins_109_ VSS VDD sg13g2_INVD1
Xins_419_ addr\[2\] ins_110_ VSS VDD sg13g2_INVD1
Xins_420_ genblk1.counter\[1\] ins_111_ VSS VDD sg13g2_INVD1
Xins_421_ genblk1.counter\[12\] ins_112_ VSS VDD sg13g2_INVD1
Xins_422_ genblk1.counter\[2\] genblk1.counter\[3\] VDD VSS
+ ins_113_ sg13g2_NR2D1
Xins_423_ genblk1.counter\[4\] encap VDD VSS ins_114_ sg13g2_NR2D1
Xins_424_ ins_021_ ins_111_ ins_113_ ins_114_ VDD VSS ins_115_
+ sg13g2_ND4D1
Xins_425_ genblk1.counter\[10\] genblk1.counter\[11\] VDD
+ VSS ins_116_ sg13g2_NR2D1
Xins_426_ genblk1.counter\[6\] genblk1.counter\[7\] VDD VSS
+ ins_117_ sg13g2_NR2D1
Xins_427_ genblk1.counter\[8\] genblk1.counter\[9\] VDD VSS
+ ins_118_ sg13g2_NR2D1
Xins_428_ ins_112_ ins_116_ ins_117_ ins_118_ VDD VSS ins_119_
+ sg13g2_ND4D1
Xins_429_ ins_115_ ins_119_ ins_022_ VDD VSS ins_120_ sg13g2_OAI21D1
Xins_430_ DATA raddr\[0\] ins_120_ VDD VSS ins_023_ sg13g2_MUX2D1
Xins_431_ raddr\[0\] raddr\[1\] ins_120_ VDD VSS ins_024_
+ sg13g2_MUX2D1
Xins_432_ raddr\[1\] raddr\[2\] ins_120_ VDD VSS ins_025_
+ sg13g2_MUX2D1
Xins_433_ raddr\[2\] sft_reg\[3\] ins_120_ VDD VSS ins_026_
+ sg13g2_MUX2D1
Xins_434_ sft_reg\[3\] sft_reg\[4\] ins_120_ VDD VSS ins_027_
+ sg13g2_MUX2D1
Xins_435_ sft_reg\[4\] sft_reg\[5\] ins_120_ VDD VSS ins_028_
+ sg13g2_MUX2D1
Xins_436_ sft_reg\[5\] sft_reg\[6\] ins_120_ VDD VSS ins_029_
+ sg13g2_MUX2D1
Xins_437_ sft_reg\[6\] sft_reg\[7\] ins_120_ VDD VSS ins_030_
+ sg13g2_MUX2D1
Xins_438_ sft_reg\[7\] addr\[0\] ins_120_ VDD VSS ins_031_
+ sg13g2_MUX2D1
Xins_439_ addr\[0\] addr\[1\] ins_120_ VDD VSS ins_032_ sg13g2_MUX2D1
Xins_440_ addr\[1\] addr\[2\] ins_120_ VDD VSS ins_033_ sg13g2_MUX2D1
Xins_441_ we genblk1.counter\[13\] VDD VSS ins_121_ sg13g2_AN2D1
Xins_442_ we genblk1.counter\[13\] VDD VSS ins_122_ sg13g2_ND2D1
Xins_443_ addr\[0\] ins_109_ addr\[2\] VDD VSS ins_123_ sg13g2_ND3D1
Xins_444_ ins_122_ ins_123_ VDD VSS ins_124_ sg13g2_NR2D1
Xins_445_ R[40] raddr\[0\] ins_124_ VDD VSS ins_034_ sg13g2_MUX2D1
Xins_446_ R[41] raddr\[1\] ins_124_ VDD VSS ins_035_ sg13g2_MUX2D1
Xins_447_ RST clknet_3_1__leaf_CLK ins_023_ raddr\[0\] VDD
+ VSS sg13g2_DFCNQD1
Xins_448_ RST clknet_3_5__leaf_CLK ins_024_ raddr\[1\] VDD
+ VSS sg13g2_DFCNQD1
Xins_449_ RST clknet_3_5__leaf_CLK ins_025_ raddr\[2\] VDD
+ VSS sg13g2_DFCNQD1
Xins_450_ RST clknet_3_5__leaf_CLK ins_026_ sft_reg\[3\] VDD
+ VSS sg13g2_DFCNQD1
Xins_451_ RST clknet_3_5__leaf_CLK ins_027_ sft_reg\[4\] VDD
+ VSS sg13g2_DFCNQD1
Xins_452_ RST clknet_3_5__leaf_CLK ins_028_ sft_reg\[5\] VDD
+ VSS sg13g2_DFCNQD1
Xins_453_ RST clknet_3_5__leaf_CLK ins_029_ sft_reg\[6\] VDD
+ VSS sg13g2_DFCNQD1
Xins_454_ RST clknet_3_7__leaf_CLK ins_030_ sft_reg\[7\] VDD
+ VSS sg13g2_DFCNQD1
Xins_455_ RST clknet_3_1__leaf_CLK ins_031_ addr\[0\] VDD
+ VSS sg13g2_DFCNQD1
Xins_456_ RST clknet_3_1__leaf_CLK ins_032_ addr\[1\] VDD
+ VSS sg13g2_DFCNQD1
Xins_457_ RST clknet_3_1__leaf_CLK ins_033_ addr\[2\] VDD
+ VSS sg13g2_DFCNQD1
Xins_458_ RST clknet_3_7__leaf_CLK ins_034_ R[40] VDD VSS
+ sg13g2_DFCNQD1
Xins_459_ RST clknet_3_6__leaf_CLK ins_035_ R[41] VDD VSS
+ sg13g2_DFCNQD1
Xins_460_ RST clknet_3_7__leaf_CLK ins_036_ R[42] VDD VSS
+ sg13g2_DFCNQD1
Xins_461_ RST clknet_3_3__leaf_CLK ins_037_ R[43] VDD VSS
+ sg13g2_DFCNQD1
Xins_462_ RST clknet_3_7__leaf_CLK ins_038_ R[44] VDD VSS
+ sg13g2_DFCNQD1
Xins_463_ RST clknet_3_7__leaf_CLK ins_039_ R[45] VDD VSS
+ sg13g2_DFCNQD1
Xins_464_ RST clknet_3_6__leaf_CLK ins_040_ R[46] VDD VSS
+ sg13g2_DFCNQD1
Xins_465_ RST clknet_3_3__leaf_CLK ins_041_ R[47] VDD VSS
+ sg13g2_DFCNQD1
Xins_466_ RST clknet_3_6__leaf_CLK ins_042_ R[0] VDD VSS sg13g2_DFCNQD1
Xins_467_ RST clknet_3_6__leaf_CLK ins_043_ R[1] VDD VSS sg13g2_DFCNQD1
Xins_468_ RST clknet_3_6__leaf_CLK ins_044_ R[2] VDD VSS sg13g2_DFCNQD1
Xins_469_ RST clknet_3_3__leaf_CLK ins_045_ R[3] VDD VSS sg13g2_DFCNQD1
Xins_470_ RST clknet_3_6__leaf_CLK ins_046_ R[4] VDD VSS sg13g2_DFCNQD1
Xins_471_ RST clknet_3_2__leaf_CLK ins_047_ R[5] VDD VSS sg13g2_DFCNQD1
Xins_472_ RST clknet_3_6__leaf_CLK ins_048_ R[6] VDD VSS sg13g2_DFCNQD1
Xins_473_ RST clknet_3_3__leaf_CLK ins_049_ R[7] VDD VSS sg13g2_DFCNQD1
Xins_474_ RST clknet_3_6__leaf_CLK ins_050_ R[16] VDD VSS
+ sg13g2_DFCNQD1
Xins_475_ RST clknet_3_4__leaf_CLK ins_051_ R[17] VDD VSS
+ sg13g2_DFCNQD1
Xins_476_ RST clknet_3_1__leaf_CLK ins_052_ R[18] VDD VSS
+ sg13g2_DFCNQD1
Xins_477_ RST clknet_3_4__leaf_CLK ins_053_ R[19] VDD VSS
+ sg13g2_DFCNQD1
Xins_478_ RST clknet_3_5__leaf_CLK ins_054_ R[20] VDD VSS
+ sg13g2_DFCNQD1
Xins_479_ RST clknet_3_1__leaf_CLK ins_055_ R[21] VDD VSS
+ sg13g2_DFCNQD1
Xins_480_ RST clknet_3_5__leaf_CLK ins_056_ R[22] VDD VSS
+ sg13g2_DFCNQD1
Xins_481_ RST clknet_3_4__leaf_CLK ins_057_ R[23] VDD VSS
+ sg13g2_DFCNQD1
Xins_482_ RST clknet_3_7__leaf_CLK ins_058_ R[56] VDD VSS
+ sg13g2_DFCNQD1
Xins_483_ RST clknet_3_7__leaf_CLK ins_059_ R[57] VDD VSS
+ sg13g2_DFCNQD1
Xins_484_ RST clknet_3_3__leaf_CLK ins_060_ R[58] VDD VSS
+ sg13g2_DFCNQD1
Xins_485_ RST clknet_3_7__leaf_CLK ins_061_ R[59] VDD VSS
+ sg13g2_DFCNQD1
Xins_486_ RST clknet_3_7__leaf_CLK ins_062_ R[60] VDD VSS
+ sg13g2_DFCNQD1
Xins_487_ RST clknet_3_2__leaf_CLK ins_063_ R[61] VDD VSS
+ sg13g2_DFCNQD1
Xins_488_ RST clknet_3_7__leaf_CLK ins_064_ R[62] VDD VSS
+ sg13g2_DFCNQD1
Xins_489_ RST clknet_3_7__leaf_CLK ins_065_ R[63] VDD VSS
+ sg13g2_DFCNQD1
Xins_490_ RST clknet_3_2__leaf_CLK ins_066_ bus_cap\[0\] VDD
+ VSS sg13g2_DFCNQD1
Xins_491_ RST clknet_3_3__leaf_CLK ins_067_ bus_cap\[1\] VDD
+ VSS sg13g2_DFCNQD1
Xins_492_ RST clknet_3_2__leaf_CLK ins_068_ bus_cap\[2\] VDD
+ VSS sg13g2_DFCNQD1
Xins_493_ RST clknet_3_2__leaf_CLK ins_069_ bus_cap\[3\] VDD
+ VSS sg13g2_DFCNQD1
Xins_494_ RST clknet_3_2__leaf_CLK ins_070_ bus_cap\[4\] VDD
+ VSS sg13g2_DFCNQD1
Xins_495_ RST clknet_3_2__leaf_CLK ins_071_ bus_cap\[5\] VDD
+ VSS sg13g2_DFCNQD1
Xins_496_ RST clknet_3_2__leaf_CLK ins_072_ bus_cap\[6\] VDD
+ VSS sg13g2_DFCNQD1
Xins_497_ RST clknet_3_2__leaf_CLK ins_073_ bus_cap\[7\] VDD
+ VSS sg13g2_DFCNQD1
Xins_498_ RST clknet_3_7__leaf_CLK ins_074_ R[48] VDD VSS
+ sg13g2_DFCNQD1
Xins_499_ RST clknet_3_7__leaf_CLK ins_075_ R[49] VDD VSS
+ sg13g2_DFCNQD1
Xins_500_ RST clknet_3_1__leaf_CLK ins_076_ R[50] VDD VSS
+ sg13g2_DFCNQD1
Xins_501_ RST clknet_3_7__leaf_CLK ins_077_ R[51] VDD VSS
+ sg13g2_DFCNQD1
Xins_502_ RST clknet_3_6__leaf_CLK ins_078_ R[52] VDD VSS
+ sg13g2_DFCNQD1
Xins_503_ RST clknet_3_7__leaf_CLK ins_079_ R[53] VDD VSS
+ sg13g2_DFCNQD1
Xins_504_ RST clknet_3_3__leaf_CLK ins_080_ R[54] VDD VSS
+ sg13g2_DFCNQD1
Xins_505_ RST clknet_3_7__leaf_CLK ins_081_ R[55] VDD VSS
+ sg13g2_DFCNQD1
Xins_506_ RST clknet_3_3__leaf_CLK ins_082_ we VDD VSS sg13g2_DFCNQD1
Xins_507_ RST clknet_3_0__leaf_CLK ins_022_ ins_021_ VDD VSS
+ sg13g2_DFCNQD1
Xins_508_ RST clknet_3_3__leaf_CLK ins_011_ genblk1.counter\[1\]
+ VDD VSS sg13g2_DFCNQD1
Xins_509_ RST clknet_3_2__leaf_CLK ins_013_ genblk1.counter\[2\]
+ VDD VSS sg13g2_DFCNQD1
Xins_510_ RST clknet_3_2__leaf_CLK ins_014_ genblk1.counter\[3\]
+ VDD VSS sg13g2_DFCNQD1
Xins_511_ RST clknet_3_2__leaf_CLK ins_015_ genblk1.counter\[4\]
+ VDD VSS sg13g2_DFCNQD1
Xins_512_ RST clknet_3_2__leaf_CLK ins_016_ encap VDD VSS
+ sg13g2_DFCNQD1
Xins_513_ RST clknet_3_0__leaf_CLK ins_017_ genblk1.counter\[6\]
+ VDD VSS sg13g2_DFCNQD1
Xins_514_ RST clknet_3_0__leaf_CLK ins_018_ genblk1.counter\[7\]
+ VDD VSS sg13g2_DFCNQD1
Xins_515_ RST clknet_3_0__leaf_CLK ins_019_ genblk1.counter\[8\]
+ VDD VSS sg13g2_DFCNQD1
Xins_516_ RST clknet_3_0__leaf_CLK ins_020_ genblk1.counter\[9\]
+ VDD VSS sg13g2_DFCNQD1
Xins_517_ RST clknet_3_0__leaf_CLK ins_001_ genblk1.counter\[10\]
+ VDD VSS sg13g2_DFCNQD1
Xins_518_ RST clknet_3_0__leaf_CLK ins_002_ genblk1.counter\[11\]
+ VDD VSS sg13g2_DFCNQD1
Xins_519_ RST clknet_3_0__leaf_CLK ins_003_ genblk1.counter\[12\]
+ VDD VSS sg13g2_DFCNQD1
Xins_520_ RST clknet_3_0__leaf_CLK ins_004_ genblk1.counter\[13\]
+ VDD VSS sg13g2_DFCNQD1
Xins_521_ RST clknet_3_0__leaf_CLK ins_005_ genblk1.counter\[14\]
+ VDD VSS sg13g2_DFCNQD1
Xins_522_ RST clknet_3_0__leaf_CLK ins_006_ genblk1.counter\[15\]
+ VDD VSS sg13g2_DFCNQD1
Xins_523_ RST clknet_3_1__leaf_CLK ins_007_ genblk1.counter\[16\]
+ VDD VSS sg13g2_DFCNQD1
Xins_524_ RST clknet_3_1__leaf_CLK ins_008_ genblk1.counter\[17\]
+ VDD VSS sg13g2_DFCNQD1
Xins_525_ RST clknet_3_1__leaf_CLK ins_009_ genblk1.counter\[18\]
+ VDD VSS sg13g2_DFCNQD1
Xins_526_ RST clknet_3_1__leaf_CLK ins_010_ genblk1.counter\[19\]
+ VDD VSS sg13g2_DFCNQD1
Xins_527_ RST clknet_3_1__leaf_CLK ins_012_ genblk1.counter\[20\]
+ VDD VSS sg13g2_DFCNQD1
Xins_528_ RST clknet_3_2__leaf_CLK eno enoz VDD VSS sg13g2_DFCNQD1
Xins_529_ RST clknet_3_2__leaf_CLK ins_000_ DOUT_DAT VDD VSS
+ sg13g2_DFCNQD1
Xins_530_ RST clknet_3_1__leaf_CLK ins_083_ R[32] VDD VSS
+ sg13g2_DFCNQD1
Xins_531_ RST clknet_3_5__leaf_CLK ins_084_ R[33] VDD VSS
+ sg13g2_DFCNQD1
Xins_532_ RST clknet_3_5__leaf_CLK ins_085_ R[34] VDD VSS
+ sg13g2_DFCNQD1
Xins_533_ RST clknet_3_7__leaf_CLK ins_086_ R[35] VDD VSS
+ sg13g2_DFCNQD1
Xins_534_ RST clknet_3_4__leaf_CLK ins_087_ R[36] VDD VSS
+ sg13g2_DFCNQD1
Xins_535_ RST clknet_3_7__leaf_CLK ins_088_ R[37] VDD VSS
+ sg13g2_DFCNQD1
Xins_536_ RST clknet_3_7__leaf_CLK ins_089_ R[38] VDD VSS
+ sg13g2_DFCNQD1
Xins_537_ RST clknet_3_4__leaf_CLK ins_090_ R[39] VDD VSS
+ sg13g2_DFCNQD1
Xins_538_ RST clknet_3_5__leaf_CLK ins_091_ R[24] VDD VSS
+ sg13g2_DFCNQD1
Xins_539_ RST clknet_3_4__leaf_CLK ins_092_ R[25] VDD VSS
+ sg13g2_DFCNQD1
Xins_540_ RST clknet_3_4__leaf_CLK ins_093_ R[26] VDD VSS
+ sg13g2_DFCNQD1
Xins_541_ RST clknet_3_5__leaf_CLK ins_094_ R[27] VDD VSS
+ sg13g2_DFCNQD1
Xins_542_ RST clknet_3_4__leaf_CLK ins_095_ R[28] VDD VSS
+ sg13g2_DFCNQD1
Xins_543_ RST clknet_3_4__leaf_CLK ins_096_ R[29] VDD VSS
+ sg13g2_DFCNQD1
Xins_544_ RST clknet_3_4__leaf_CLK ins_097_ R[30] VDD VSS
+ sg13g2_DFCNQD1
Xins_545_ RST clknet_3_4__leaf_CLK ins_098_ R[31] VDD VSS
+ sg13g2_DFCNQD1
Xins_546_ RST clknet_3_6__leaf_CLK ins_099_ R[8] VDD VSS sg13g2_DFCNQD1
Xins_547_ RST clknet_3_7__leaf_CLK ins_100_ R[9] VDD VSS sg13g2_DFCNQD1
Xins_548_ RST clknet_3_3__leaf_CLK ins_101_ R[10] VDD VSS
+ sg13g2_DFCNQD1
Xins_549_ RST clknet_3_6__leaf_CLK ins_102_ R[11] VDD VSS
+ sg13g2_DFCNQD1
Xins_550_ RST clknet_3_6__leaf_CLK ins_103_ R[12] VDD VSS
+ sg13g2_DFCNQD1
Xins_551_ RST clknet_3_6__leaf_CLK ins_104_ R[13] VDD VSS
+ sg13g2_DFCNQD1
Xins_552_ RST clknet_3_3__leaf_CLK ins_105_ R[14] VDD VSS
+ sg13g2_DFCNQD1
Xins_553_ RST clknet_3_6__leaf_CLK ins_106_ R[15] VDD VSS
+ sg13g2_DFCNQD1
Xins_554_ RST clknet_3_0__leaf_CLK ins_107_ re VDD VSS sg13g2_DFCNQD1
Xclkbuf_0_CLK CLK VDD VSS clknet_0_CLK sg13g2_BUFFD1
Xclkbuf_3_0__f_CLK clknet_0_CLK VDD VSS clknet_3_0__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_1__f_CLK clknet_0_CLK VDD VSS clknet_3_1__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_2__f_CLK clknet_0_CLK VDD VSS clknet_3_2__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_3__f_CLK clknet_0_CLK VDD VSS clknet_3_3__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_4__f_CLK clknet_0_CLK VDD VSS clknet_3_4__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_5__f_CLK clknet_0_CLK VDD VSS clknet_3_5__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_6__f_CLK clknet_0_CLK VDD VSS clknet_3_6__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_7__f_CLK clknet_0_CLK VDD VSS clknet_3_7__leaf_CLK
+ sg13g2_BUFFD1
Xclkload0 clknet_3_0__leaf_CLK _unconnected_0 VSS VDD sg13g2_INVD1
Xclkload1 clknet_3_1__leaf_CLK _unconnected_1 VSS VDD sg13g2_INVD1
Xclkload2 clknet_3_2__leaf_CLK _unconnected_2 VSS VDD sg13g2_INVD1
Xclkload3 clknet_3_3__leaf_CLK _unconnected_3 VSS VDD sg13g2_INVD1
Xclkload4 clknet_3_4__leaf_CLK _unconnected_4 VSS VDD sg13g2_INVD1
Xclkload5 clknet_3_5__leaf_CLK _unconnected_5 VSS VDD sg13g2_INVD1
Xclkload6 clknet_3_6__leaf_CLK _unconnected_6 VSS VDD sg13g2_INVD1
XFILLER_0_0 VDD VSS sg13g2_FILL8
XFILLER_0_8 VDD VSS sg13g2_FILL8
XFILLER_0_16 VDD VSS sg13g2_FILL8
XFILLER_0_24 VDD VSS sg13g2_FILL8
XFILLER_0_32 VDD VSS sg13g2_FILL8
XFILLER_0_40 VDD VSS sg13g2_FILL8
XFILLER_0_48 VDD VSS sg13g2_FILL8
XFILLER_0_56 VDD VSS sg13g2_FILL8
XFILLER_0_64 VDD VSS sg13g2_FILL8
XFILLER_0_72 VDD VSS sg13g2_FILL4
XFILLER_0_76 VDD VSS sg13g2_FILL1
XFILLER_0_90 VDD VSS sg13g2_FILL4
XFILLER_0_94 VDD VSS sg13g2_FILL2
XFILLER_0_146 VDD VSS sg13g2_FILL8
XFILLER_0_154 VDD VSS sg13g2_FILL8
XFILLER_0_162 VDD VSS sg13g2_FILL4
XFILLER_0_179 VDD VSS sg13g2_FILL8
XFILLER_0_187 VDD VSS sg13g2_FILL8
XFILLER_0_195 VDD VSS sg13g2_FILL2
XFILLER_0_255 VDD VSS sg13g2_FILL4
XFILLER_0_272 VDD VSS sg13g2_FILL8
XFILLER_0_280 VDD VSS sg13g2_FILL2
XFILLER_0_358 VDD VSS sg13g2_FILL8
XFILLER_0_366 VDD VSS sg13g2_FILL4
XFILLER_0_370 VDD VSS sg13g2_FILL1
XFILLER_0_465 VDD VSS sg13g2_FILL8
XFILLER_0_473 VDD VSS sg13g2_FILL8
XFILLER_0_481 VDD VSS sg13g2_FILL2
XFILLER_0_505 VDD VSS sg13g2_FILL8
XFILLER_0_513 VDD VSS sg13g2_FILL8
XFILLER_0_571 VDD VSS sg13g2_FILL4
XFILLER_0_625 VDD VSS sg13g2_FILL8
XFILLER_0_633 VDD VSS sg13g2_FILL8
XFILLER_0_641 VDD VSS sg13g2_FILL8
XFILLER_0_699 VDD VSS sg13g2_FILL8
XFILLER_0_707 VDD VSS sg13g2_FILL8
XFILLER_0_715 VDD VSS sg13g2_FILL1
XFILLER_0_738 VDD VSS sg13g2_FILL8
XFILLER_0_746 VDD VSS sg13g2_FILL8
XFILLER_0_754 VDD VSS sg13g2_FILL8
XFILLER_0_762 VDD VSS sg13g2_FILL8
XFILLER_0_770 VDD VSS sg13g2_FILL8
XFILLER_0_778 VDD VSS sg13g2_FILL8
XFILLER_0_786 VDD VSS sg13g2_FILL8
XFILLER_0_794 VDD VSS sg13g2_FILL8
XFILLER_0_802 VDD VSS sg13g2_FILL4
XFILLER_0_806 VDD VSS sg13g2_FILL2
XFILLER_1_0 VDD VSS sg13g2_FILL8
XFILLER_1_8 VDD VSS sg13g2_FILL8
XFILLER_1_16 VDD VSS sg13g2_FILL8
XFILLER_1_24 VDD VSS sg13g2_FILL8
XFILLER_1_32 VDD VSS sg13g2_FILL8
XFILLER_1_40 VDD VSS sg13g2_FILL8
XFILLER_1_98 VDD VSS sg13g2_FILL2
XFILLER_1_171 VDD VSS sg13g2_FILL4
XFILLER_1_175 VDD VSS sg13g2_FILL2
XFILLER_1_177 VDD VSS sg13g2_FILL1
XFILLER_1_304 VDD VSS sg13g2_FILL2
XFILLER_1_356 VDD VSS sg13g2_FILL2
XFILLER_1_358 VDD VSS sg13g2_FILL1
XFILLER_1_781 VDD VSS sg13g2_FILL8
XFILLER_1_789 VDD VSS sg13g2_FILL8
XFILLER_1_797 VDD VSS sg13g2_FILL8
XFILLER_1_805 VDD VSS sg13g2_FILL2
XFILLER_1_807 VDD VSS sg13g2_FILL1
XFILLER_2_0 VDD VSS sg13g2_FILL8
XFILLER_2_8 VDD VSS sg13g2_FILL8
XFILLER_2_16 VDD VSS sg13g2_FILL8
XFILLER_2_24 VDD VSS sg13g2_FILL4
XFILLER_2_28 VDD VSS sg13g2_FILL1
XFILLER_2_137 VDD VSS sg13g2_FILL4
XFILLER_2_241 VDD VSS sg13g2_FILL2
XFILLER_2_267 VDD VSS sg13g2_FILL4
XFILLER_2_271 VDD VSS sg13g2_FILL1
XFILLER_2_485 VDD VSS sg13g2_FILL8
XFILLER_2_493 VDD VSS sg13g2_FILL8
XFILLER_2_617 VDD VSS sg13g2_FILL4
XFILLER_2_621 VDD VSS sg13g2_FILL1
XFILLER_2_679 VDD VSS sg13g2_FILL8
XFILLER_2_787 VDD VSS sg13g2_FILL8
XFILLER_2_795 VDD VSS sg13g2_FILL8
XFILLER_2_803 VDD VSS sg13g2_FILL4
XFILLER_2_807 VDD VSS sg13g2_FILL1
XFILLER_3_0 VDD VSS sg13g2_FILL8
XFILLER_3_8 VDD VSS sg13g2_FILL8
XFILLER_3_16 VDD VSS sg13g2_FILL8
XFILLER_3_24 VDD VSS sg13g2_FILL4
XFILLER_3_28 VDD VSS sg13g2_FILL2
XFILLER_3_106 VDD VSS sg13g2_FILL1
XFILLER_3_136 VDD VSS sg13g2_FILL1
XFILLER_3_203 VDD VSS sg13g2_FILL8
XFILLER_3_211 VDD VSS sg13g2_FILL4
XFILLER_3_215 VDD VSS sg13g2_FILL1
XFILLER_3_279 VDD VSS sg13g2_FILL2
XFILLER_3_281 VDD VSS sg13g2_FILL1
XFILLER_3_375 VDD VSS sg13g2_FILL2
XFILLER_3_377 VDD VSS sg13g2_FILL1
XFILLER_3_422 VDD VSS sg13g2_FILL8
XFILLER_3_430 VDD VSS sg13g2_FILL4
XFILLER_3_434 VDD VSS sg13g2_FILL2
XFILLER_3_458 VDD VSS sg13g2_FILL8
XFILLER_3_466 VDD VSS sg13g2_FILL8
XFILLER_3_474 VDD VSS sg13g2_FILL8
XFILLER_3_482 VDD VSS sg13g2_FILL8
XFILLER_3_490 VDD VSS sg13g2_FILL2
XFILLER_3_492 VDD VSS sg13g2_FILL1
XFILLER_3_600 VDD VSS sg13g2_FILL2
XFILLER_3_602 VDD VSS sg13g2_FILL1
XFILLER_3_719 VDD VSS sg13g2_FILL4
XFILLER_3_723 VDD VSS sg13g2_FILL2
XFILLER_3_775 VDD VSS sg13g2_FILL8
XFILLER_3_783 VDD VSS sg13g2_FILL8
XFILLER_3_791 VDD VSS sg13g2_FILL8
XFILLER_3_799 VDD VSS sg13g2_FILL8
XFILLER_3_807 VDD VSS sg13g2_FILL1
XFILLER_4_0 VDD VSS sg13g2_FILL8
XFILLER_4_8 VDD VSS sg13g2_FILL8
XFILLER_4_16 VDD VSS sg13g2_FILL8
XFILLER_4_24 VDD VSS sg13g2_FILL8
XFILLER_4_32 VDD VSS sg13g2_FILL4
XFILLER_4_36 VDD VSS sg13g2_FILL1
XFILLER_4_87 VDD VSS sg13g2_FILL4
XFILLER_4_91 VDD VSS sg13g2_FILL1
XFILLER_4_121 VDD VSS sg13g2_FILL1
XFILLER_4_190 VDD VSS sg13g2_FILL1
XFILLER_4_221 VDD VSS sg13g2_FILL4
XFILLER_4_225 VDD VSS sg13g2_FILL2
XFILLER_4_227 VDD VSS sg13g2_FILL1
XFILLER_4_300 VDD VSS sg13g2_FILL8
XFILLER_4_308 VDD VSS sg13g2_FILL4
XFILLER_4_312 VDD VSS sg13g2_FILL2
XFILLER_4_322 VDD VSS sg13g2_FILL2
XFILLER_4_324 VDD VSS sg13g2_FILL1
XFILLER_4_375 VDD VSS sg13g2_FILL8
XFILLER_4_383 VDD VSS sg13g2_FILL2
XFILLER_4_385 VDD VSS sg13g2_FILL1
XFILLER_4_486 VDD VSS sg13g2_FILL8
XFILLER_4_494 VDD VSS sg13g2_FILL8
XFILLER_4_502 VDD VSS sg13g2_FILL8
XFILLER_4_510 VDD VSS sg13g2_FILL1
XFILLER_4_583 VDD VSS sg13g2_FILL8
XFILLER_4_591 VDD VSS sg13g2_FILL8
XFILLER_4_599 VDD VSS sg13g2_FILL2
XFILLER_4_601 VDD VSS sg13g2_FILL1
XFILLER_4_674 VDD VSS sg13g2_FILL8
XFILLER_4_682 VDD VSS sg13g2_FILL8
XFILLER_4_690 VDD VSS sg13g2_FILL4
XFILLER_4_694 VDD VSS sg13g2_FILL1
XFILLER_4_789 VDD VSS sg13g2_FILL8
XFILLER_4_797 VDD VSS sg13g2_FILL8
XFILLER_4_805 VDD VSS sg13g2_FILL2
XFILLER_4_807 VDD VSS sg13g2_FILL1
XFILLER_5_0 VDD VSS sg13g2_FILL8
XFILLER_5_8 VDD VSS sg13g2_FILL8
XFILLER_5_16 VDD VSS sg13g2_FILL8
XFILLER_5_24 VDD VSS sg13g2_FILL4
XFILLER_5_28 VDD VSS sg13g2_FILL1
XFILLER_5_92 VDD VSS sg13g2_FILL2
XFILLER_5_107 VDD VSS sg13g2_FILL8
XFILLER_5_115 VDD VSS sg13g2_FILL8
XFILLER_5_123 VDD VSS sg13g2_FILL1
XFILLER_5_245 VDD VSS sg13g2_FILL8
XFILLER_5_253 VDD VSS sg13g2_FILL4
XFILLER_5_401 VDD VSS sg13g2_FILL8
XFILLER_5_409 VDD VSS sg13g2_FILL4
XFILLER_5_413 VDD VSS sg13g2_FILL1
XFILLER_5_514 VDD VSS sg13g2_FILL8
XFILLER_5_522 VDD VSS sg13g2_FILL4
XFILLER_5_526 VDD VSS sg13g2_FILL2
XFILLER_5_528 VDD VSS sg13g2_FILL1
XFILLER_5_601 VDD VSS sg13g2_FILL8
XFILLER_5_609 VDD VSS sg13g2_FILL8
XFILLER_5_617 VDD VSS sg13g2_FILL4
XFILLER_5_621 VDD VSS sg13g2_FILL1
XFILLER_5_672 VDD VSS sg13g2_FILL8
XFILLER_5_702 VDD VSS sg13g2_FILL4
XFILLER_5_706 VDD VSS sg13g2_FILL2
XFILLER_5_708 VDD VSS sg13g2_FILL1
XFILLER_5_781 VDD VSS sg13g2_FILL8
XFILLER_5_789 VDD VSS sg13g2_FILL8
XFILLER_5_797 VDD VSS sg13g2_FILL8
XFILLER_5_805 VDD VSS sg13g2_FILL2
XFILLER_5_807 VDD VSS sg13g2_FILL1
XFILLER_6_0 VDD VSS sg13g2_FILL8
XFILLER_6_8 VDD VSS sg13g2_FILL8
XFILLER_6_16 VDD VSS sg13g2_FILL8
XFILLER_6_24 VDD VSS sg13g2_FILL8
XFILLER_6_32 VDD VSS sg13g2_FILL2
XFILLER_6_206 VDD VSS sg13g2_FILL8
XFILLER_6_214 VDD VSS sg13g2_FILL8
XFILLER_6_222 VDD VSS sg13g2_FILL4
XFILLER_6_299 VDD VSS sg13g2_FILL4
XFILLER_6_303 VDD VSS sg13g2_FILL2
XFILLER_6_377 VDD VSS sg13g2_FILL8
XFILLER_6_385 VDD VSS sg13g2_FILL1
XFILLER_6_500 VDD VSS sg13g2_FILL8
XFILLER_6_508 VDD VSS sg13g2_FILL4
XFILLER_6_512 VDD VSS sg13g2_FILL2
XFILLER_6_514 VDD VSS sg13g2_FILL1
XFILLER_6_587 VDD VSS sg13g2_FILL8
XFILLER_6_595 VDD VSS sg13g2_FILL8
XFILLER_6_603 VDD VSS sg13g2_FILL2
XFILLER_6_677 VDD VSS sg13g2_FILL4
XFILLER_6_731 VDD VSS sg13g2_FILL4
XFILLER_6_807 VDD VSS sg13g2_FILL1
XFILLER_7_0 VDD VSS sg13g2_FILL8
XFILLER_7_8 VDD VSS sg13g2_FILL8
XFILLER_7_16 VDD VSS sg13g2_FILL8
XFILLER_7_24 VDD VSS sg13g2_FILL8
XFILLER_7_32 VDD VSS sg13g2_FILL8
XFILLER_7_40 VDD VSS sg13g2_FILL8
XFILLER_7_48 VDD VSS sg13g2_FILL8
XFILLER_7_56 VDD VSS sg13g2_FILL8
XFILLER_7_64 VDD VSS sg13g2_FILL8
XFILLER_7_85 VDD VSS sg13g2_FILL8
XFILLER_7_93 VDD VSS sg13g2_FILL4
XFILLER_7_97 VDD VSS sg13g2_FILL1
XFILLER_7_106 VDD VSS sg13g2_FILL8
XFILLER_7_114 VDD VSS sg13g2_FILL8
XFILLER_7_122 VDD VSS sg13g2_FILL4
XFILLER_7_126 VDD VSS sg13g2_FILL2
XFILLER_7_171 VDD VSS sg13g2_FILL8
XFILLER_7_179 VDD VSS sg13g2_FILL4
XFILLER_7_191 VDD VSS sg13g2_FILL8
XFILLER_7_199 VDD VSS sg13g2_FILL8
XFILLER_7_207 VDD VSS sg13g2_FILL2
XFILLER_7_214 VDD VSS sg13g2_FILL4
XFILLER_7_218 VDD VSS sg13g2_FILL1
XFILLER_7_249 VDD VSS sg13g2_FILL4
XFILLER_7_299 VDD VSS sg13g2_FILL4
XFILLER_7_324 VDD VSS sg13g2_FILL8
XFILLER_7_332 VDD VSS sg13g2_FILL8
XFILLER_7_340 VDD VSS sg13g2_FILL4
XFILLER_7_344 VDD VSS sg13g2_FILL1
XFILLER_7_367 VDD VSS sg13g2_FILL8
XFILLER_7_375 VDD VSS sg13g2_FILL8
XFILLER_7_383 VDD VSS sg13g2_FILL2
XFILLER_7_401 VDD VSS sg13g2_FILL1
XFILLER_7_423 VDD VSS sg13g2_FILL2
XFILLER_7_425 VDD VSS sg13g2_FILL1
XFILLER_7_476 VDD VSS sg13g2_FILL4
XFILLER_7_502 VDD VSS sg13g2_FILL8
XFILLER_7_510 VDD VSS sg13g2_FILL8
XFILLER_7_518 VDD VSS sg13g2_FILL4
XFILLER_7_566 VDD VSS sg13g2_FILL8
XFILLER_7_574 VDD VSS sg13g2_FILL8
XFILLER_7_582 VDD VSS sg13g2_FILL2
XFILLER_7_584 VDD VSS sg13g2_FILL1
XFILLER_7_607 VDD VSS sg13g2_FILL8
XFILLER_7_615 VDD VSS sg13g2_FILL8
XFILLER_7_623 VDD VSS sg13g2_FILL4
XFILLER_7_649 VDD VSS sg13g2_FILL4
XFILLER_7_653 VDD VSS sg13g2_FILL2
XFILLER_7_677 VDD VSS sg13g2_FILL8
XFILLER_7_685 VDD VSS sg13g2_FILL8
XFILLER_7_693 VDD VSS sg13g2_FILL4
XFILLER_7_791 VDD VSS sg13g2_FILL8
XFILLER_7_799 VDD VSS sg13g2_FILL8
XFILLER_7_807 VDD VSS sg13g2_FILL1
XFILLER_8_0 VDD VSS sg13g2_FILL8
XFILLER_8_8 VDD VSS sg13g2_FILL8
XFILLER_8_16 VDD VSS sg13g2_FILL8
XFILLER_8_24 VDD VSS sg13g2_FILL8
XFILLER_8_32 VDD VSS sg13g2_FILL8
XFILLER_8_40 VDD VSS sg13g2_FILL8
XFILLER_8_48 VDD VSS sg13g2_FILL2
XFILLER_8_50 VDD VSS sg13g2_FILL1
XFILLER_8_95 VDD VSS sg13g2_FILL2
XFILLER_8_97 VDD VSS sg13g2_FILL1
XFILLER_8_161 VDD VSS sg13g2_FILL8
XFILLER_8_169 VDD VSS sg13g2_FILL2
XFILLER_8_184 VDD VSS sg13g2_FILL1
XFILLER_8_379 VDD VSS sg13g2_FILL8
XFILLER_8_387 VDD VSS sg13g2_FILL8
XFILLER_8_395 VDD VSS sg13g2_FILL1
XFILLER_8_522 VDD VSS sg13g2_FILL8
XFILLER_8_530 VDD VSS sg13g2_FILL8
XFILLER_8_538 VDD VSS sg13g2_FILL4
XFILLER_8_542 VDD VSS sg13g2_FILL2
XFILLER_8_544 VDD VSS sg13g2_FILL1
XFILLER_8_645 VDD VSS sg13g2_FILL8
XFILLER_8_653 VDD VSS sg13g2_FILL1
XFILLER_8_704 VDD VSS sg13g2_FILL4
XFILLER_8_708 VDD VSS sg13g2_FILL1
XFILLER_8_789 VDD VSS sg13g2_FILL8
XFILLER_8_797 VDD VSS sg13g2_FILL8
XFILLER_8_805 VDD VSS sg13g2_FILL2
XFILLER_8_807 VDD VSS sg13g2_FILL1
XFILLER_9_0 VDD VSS sg13g2_FILL8
XFILLER_9_8 VDD VSS sg13g2_FILL8
XFILLER_9_16 VDD VSS sg13g2_FILL8
XFILLER_9_24 VDD VSS sg13g2_FILL2
XFILLER_9_26 VDD VSS sg13g2_FILL1
XFILLER_9_77 VDD VSS sg13g2_FILL1
XFILLER_9_178 VDD VSS sg13g2_FILL8
XFILLER_9_186 VDD VSS sg13g2_FILL8
XFILLER_9_194 VDD VSS sg13g2_FILL8
XFILLER_9_202 VDD VSS sg13g2_FILL8
XFILLER_9_210 VDD VSS sg13g2_FILL8
XFILLER_9_218 VDD VSS sg13g2_FILL4
XFILLER_9_222 VDD VSS sg13g2_FILL1
XFILLER_9_402 VDD VSS sg13g2_FILL8
XFILLER_9_410 VDD VSS sg13g2_FILL8
XFILLER_9_418 VDD VSS sg13g2_FILL4
XFILLER_9_422 VDD VSS sg13g2_FILL2
XFILLER_9_429 VDD VSS sg13g2_FILL1
XFILLER_9_463 VDD VSS sg13g2_FILL1
XFILLER_9_514 VDD VSS sg13g2_FILL8
XFILLER_9_522 VDD VSS sg13g2_FILL4
XFILLER_9_526 VDD VSS sg13g2_FILL2
XFILLER_9_528 VDD VSS sg13g2_FILL1
XFILLER_9_601 VDD VSS sg13g2_FILL8
XFILLER_9_609 VDD VSS sg13g2_FILL8
XFILLER_9_617 VDD VSS sg13g2_FILL2
XFILLER_9_619 VDD VSS sg13g2_FILL1
XFILLER_9_770 VDD VSS sg13g2_FILL8
XFILLER_9_778 VDD VSS sg13g2_FILL8
XFILLER_9_786 VDD VSS sg13g2_FILL8
XFILLER_9_794 VDD VSS sg13g2_FILL8
XFILLER_9_802 VDD VSS sg13g2_FILL4
XFILLER_9_806 VDD VSS sg13g2_FILL2
XFILLER_10_0 VDD VSS sg13g2_FILL8
XFILLER_10_8 VDD VSS sg13g2_FILL8
XFILLER_10_16 VDD VSS sg13g2_FILL4
XFILLER_10_20 VDD VSS sg13g2_FILL1
XFILLER_10_181 VDD VSS sg13g2_FILL8
XFILLER_10_189 VDD VSS sg13g2_FILL8
XFILLER_10_197 VDD VSS sg13g2_FILL8
XFILLER_10_205 VDD VSS sg13g2_FILL8
XFILLER_10_213 VDD VSS sg13g2_FILL4
XFILLER_10_217 VDD VSS sg13g2_FILL2
XFILLER_10_219 VDD VSS sg13g2_FILL1
XFILLER_10_291 VDD VSS sg13g2_FILL4
XFILLER_10_382 VDD VSS sg13g2_FILL1
XFILLER_10_522 VDD VSS sg13g2_FILL8
XFILLER_10_530 VDD VSS sg13g2_FILL1
XFILLER_10_553 VDD VSS sg13g2_FILL1
XFILLER_10_692 VDD VSS sg13g2_FILL8
XFILLER_10_700 VDD VSS sg13g2_FILL1
XFILLER_10_767 VDD VSS sg13g2_FILL8
XFILLER_10_775 VDD VSS sg13g2_FILL8
XFILLER_10_783 VDD VSS sg13g2_FILL8
XFILLER_10_791 VDD VSS sg13g2_FILL8
XFILLER_10_799 VDD VSS sg13g2_FILL8
XFILLER_10_807 VDD VSS sg13g2_FILL1
XFILLER_11_0 VDD VSS sg13g2_FILL8
XFILLER_11_8 VDD VSS sg13g2_FILL8
XFILLER_11_16 VDD VSS sg13g2_FILL8
XFILLER_11_24 VDD VSS sg13g2_FILL2
XFILLER_11_76 VDD VSS sg13g2_FILL4
XFILLER_11_179 VDD VSS sg13g2_FILL1
XFILLER_11_230 VDD VSS sg13g2_FILL4
XFILLER_11_267 VDD VSS sg13g2_FILL2
XFILLER_11_314 VDD VSS sg13g2_FILL4
XFILLER_11_318 VDD VSS sg13g2_FILL2
XFILLER_11_320 VDD VSS sg13g2_FILL1
XFILLER_11_337 VDD VSS sg13g2_FILL2
XFILLER_11_374 VDD VSS sg13g2_FILL2
XFILLER_11_392 VDD VSS sg13g2_FILL4
XFILLER_11_396 VDD VSS sg13g2_FILL1
XFILLER_11_429 VDD VSS sg13g2_FILL2
XFILLER_11_431 VDD VSS sg13g2_FILL1
XFILLER_11_448 VDD VSS sg13g2_FILL4
XFILLER_11_481 VDD VSS sg13g2_FILL2
XFILLER_11_483 VDD VSS sg13g2_FILL1
XFILLER_11_542 VDD VSS sg13g2_FILL8
XFILLER_11_550 VDD VSS sg13g2_FILL2
XFILLER_11_552 VDD VSS sg13g2_FILL1
XFILLER_11_616 VDD VSS sg13g2_FILL8
XFILLER_11_624 VDD VSS sg13g2_FILL1
XFILLER_11_675 VDD VSS sg13g2_FILL8
XFILLER_11_683 VDD VSS sg13g2_FILL8
XFILLER_11_691 VDD VSS sg13g2_FILL2
XFILLER_11_787 VDD VSS sg13g2_FILL8
XFILLER_11_795 VDD VSS sg13g2_FILL8
XFILLER_11_803 VDD VSS sg13g2_FILL4
XFILLER_11_807 VDD VSS sg13g2_FILL1
XFILLER_12_0 VDD VSS sg13g2_FILL8
XFILLER_12_8 VDD VSS sg13g2_FILL4
XFILLER_12_12 VDD VSS sg13g2_FILL2
XFILLER_12_14 VDD VSS sg13g2_FILL1
XFILLER_12_115 VDD VSS sg13g2_FILL1
XFILLER_12_166 VDD VSS sg13g2_FILL4
XFILLER_12_186 VDD VSS sg13g2_FILL2
XFILLER_12_260 VDD VSS sg13g2_FILL2
XFILLER_12_262 VDD VSS sg13g2_FILL1
XFILLER_12_468 VDD VSS sg13g2_FILL2
XFILLER_12_531 VDD VSS sg13g2_FILL8
XFILLER_12_539 VDD VSS sg13g2_FILL4
XFILLER_12_615 VDD VSS sg13g2_FILL4
XFILLER_12_619 VDD VSS sg13g2_FILL2
XFILLER_12_621 VDD VSS sg13g2_FILL1
XFILLER_12_672 VDD VSS sg13g2_FILL8
XFILLER_12_680 VDD VSS sg13g2_FILL2
XFILLER_12_682 VDD VSS sg13g2_FILL1
XFILLER_12_733 VDD VSS sg13g2_FILL4
XFILLER_12_737 VDD VSS sg13g2_FILL2
XFILLER_12_739 VDD VSS sg13g2_FILL1
XFILLER_12_790 VDD VSS sg13g2_FILL8
XFILLER_12_798 VDD VSS sg13g2_FILL8
XFILLER_12_806 VDD VSS sg13g2_FILL2
XFILLER_13_0 VDD VSS sg13g2_FILL8
XFILLER_13_8 VDD VSS sg13g2_FILL8
XFILLER_13_16 VDD VSS sg13g2_FILL8
XFILLER_13_24 VDD VSS sg13g2_FILL4
XFILLER_13_129 VDD VSS sg13g2_FILL8
XFILLER_13_137 VDD VSS sg13g2_FILL8
XFILLER_13_145 VDD VSS sg13g2_FILL8
XFILLER_13_153 VDD VSS sg13g2_FILL8
XFILLER_13_177 VDD VSS sg13g2_FILL8
XFILLER_13_185 VDD VSS sg13g2_FILL4
XFILLER_13_189 VDD VSS sg13g2_FILL1
XFILLER_13_203 VDD VSS sg13g2_FILL8
XFILLER_13_211 VDD VSS sg13g2_FILL8
XFILLER_13_219 VDD VSS sg13g2_FILL1
XFILLER_13_242 VDD VSS sg13g2_FILL2
XFILLER_13_307 VDD VSS sg13g2_FILL1
XFILLER_13_324 VDD VSS sg13g2_FILL4
XFILLER_13_328 VDD VSS sg13g2_FILL2
XFILLER_13_330 VDD VSS sg13g2_FILL1
XFILLER_13_397 VDD VSS sg13g2_FILL2
XFILLER_13_399 VDD VSS sg13g2_FILL1
XFILLER_13_426 VDD VSS sg13g2_FILL2
XFILLER_13_428 VDD VSS sg13g2_FILL1
XFILLER_13_550 VDD VSS sg13g2_FILL8
XFILLER_13_558 VDD VSS sg13g2_FILL8
XFILLER_13_588 VDD VSS sg13g2_FILL8
XFILLER_13_596 VDD VSS sg13g2_FILL1
XFILLER_13_669 VDD VSS sg13g2_FILL4
XFILLER_13_695 VDD VSS sg13g2_FILL8
XFILLER_13_703 VDD VSS sg13g2_FILL2
XFILLER_13_805 VDD VSS sg13g2_FILL2
XFILLER_13_807 VDD VSS sg13g2_FILL1
.ENDS SPI
.inc "/opt/ext/OpenPDKs/IHP-Open-PDK/ihp-sg13g2/libs.ref/sg13g2_stdcell/cdl/sg13g2_stdcell.cdl"
*.inc sg13g2_stdcell.cdl

** sch_path: xschem/inv1.sch
.subckt inv1 n_RO_control VDD VSS Vin Vout
M1 net1 n_RO_control VDD VDD sg13_lv_pmos w=3.4u l=0.45u ng=1 m=12
M5 Vout Vin net1 VDD sg13_lv_pmos w=3.4u l=0.45u ng=1 m=4
M2 VSS Vin Vout VSS sg13_lv_nmos w=1.3u l=0.45u ng=1 m=4
.ends

** sch_path: xschem/tristate_inv.sch
.subckt tristate_inv VDD VSS Vin Vup Vdn Vout
M5 Vout Vin net1 VDD sg13_lv_pmos w=3.4u l=0.45u ng=1 m=4
M2 net2 Vin Vout VSS sg13_lv_nmos w=1.3u l=0.45u ng=1 m=4
M1 net1 Vup VDD VDD sg13_lv_pmos w=3.4u l=0.45u ng=1 m=12
M3 VSS Vdn net2 VSS sg13_lv_nmos w=1.3u l=0.45u ng=1 m=12
.ends

** sch_path: xschem/inverter_RO_rel.sch
.subckt inverter_RO_rel VDD Vin Vout VSS
M3 Vout Vin VDD VDD sg13_lv_pmos w=3.4u l=0.45u ng=1 m=4
M1 VSS Vin Vout VSS sg13_lv_nmos w=1.3u l=0.45u ng=1 m=4
.ends

** sch_path: xschem/tgate_force.sch
.subckt tgate_force nclk VDD Vin Vout VSS clk
M3 Vout nclk Vin VDD sg13_lv_pmos w=3.4u l=0.45u ng=1 m=4
M4 Vout clk Vin VSS sg13_lv_nmos w=1.3u l=0.45u ng=1 m=4
.ends

** sch_path: xschem/tgate_force10.sch
.subckt tgate_force10 nclk VDD Vin Vout VSS clk
*.PININFO nclk:B clk:B VDD:B VSS:B Vout:B Vin:B
M1 Vout nclk Vin VDD sg13_lv_pmos w=3.4u l=0.45u ng=1 m=12
M3 Vout clk Vin VSS sg13_lv_nmos w=1.3u l=0.45u ng=1 m=12
.ends

** sch_path: xschem/tgate.sch
.subckt tgate nclk VDD Vin Vout VSS clk
M3 Vout nclk Vin VDD sg13_lv_pmos l=0.45u w=3.4u ng=1 m=1
M1 Vout clk Vin VSS sg13_lv_nmos l=0.45u w=1.3u ng=1 m=1
.ends

** sch_path: xschem/rovcel1.sch
.subckt rovcel1 DUT_Header DUT_Footer Drain_Force Drain_Sense RO_control n_RO_control VDD VSS Vin Vout
x4 VDD VSS Vin DUT_Header DUT_Footer Vout tristate_inv
x1 RO_control VDD Vout Drain_Force VSS n_RO_control tgate_force
x3 RO_control VDD Vout Drain_Sense VSS n_RO_control tgate
.ends

** sch_path: xschem/rovcel2.sch
.subckt rovcel2 VDD VSS Vout Vin
x5 VDD Vin Vout VSS inverter_RO_rel
x1 VDD VDD Vout net2 VSS VSS tgate
x3 VDD VDD Vout net1 VSS VSS tgate
.ends

** sch_path: xschem/rovcel3.sch
.subckt rovcel3 VDD VSS Vin n_RO_control Vout RO_control DUT_gate
x4 VDD VSS Vin n_RO_control RO_control Vout tristate_inv
x1 RO_control VDD Vout net1 VSS n_RO_control tgate
x5 RO_control VDD Vout DUT_gate VSS n_RO_control tgate
.ends

** sch_path: xschem/rovcel4.sch
.subckt rovcel4 VDD VSS Vin n_RO_control Vout
x4 n_RO_control VDD VSS Vin Vout inv1
x1 VDD VDD Vout VSS VSS VSS tgate
x5 VDD VDD Vout net1 VSS VSS tgate
.ends

** sch_path: xschem/top_RO_core_13.sch
.subckt top_RO_core_13 VDD VSS n_RO_control RO_control DUT_gate Vout DUT_Header DUT_Footer Drain_Force Drain_Sense extra_load
*.iopin VDD
*.iopin VSS
*.iopin n_RO_control
*.iopin RO_control
*.iopin DUT_gate
*.iopin extra_load
*.iopin DUT_Header
*.iopin DUT_Footer
*.iopin Drain_Force
*.iopin Drain_Sense
*.iopin Vout
x1 VDD VSS A[9] A[8] rovcel2
x7 VDD VSS A[9] n_RO_control A_10 RO_control DUT_gate rovcel3
x2 DUT_Header DUT_Footer Drain_Force Drain_Sense RO_control n_RO_control VDD VSS A_10 extra_load rovcel1
x3 VDD VSS extra_load n_RO_control A_12 rovcel4
x4 VDD VSS Vout A_12 rovcel2
x5[1] VDD VSS A[8] A[7] rovcel2
x5[2] VDD VSS A[7] A[6] rovcel2
x5[3] VDD VSS A[6] A[5] rovcel2
x5[4] VDD VSS A[5] A[4] rovcel2
x5[5] VDD VSS A[4] A[3] rovcel2
x5[6] VDD VSS A[3] A[2] rovcel2
x5[7] VDD VSS A[2] A[1] rovcel2
x5[8] VDD VSS A[1] Vout rovcel2
.ends

** sch_path: xschem/div_sg13g2_stdcells.sch
.subckt div_sg13g2_stdcells VDD OUT IN GND RSTB
x2 q2 qn2 q1 qn2 RSTB VDD GND sg13g2_dfrbp_1
x1 q1 qn1 IN qn1 RSTB VDD GND sg13g2_dfrbp_1
x3 q3 qn3 q2 qn3 RSTB VDD GND sg13g2_dfrbp_1
x4 q4 qn4 q3 qn4 RSTB VDD GND sg13g2_dfrbp_1
x5 OUT qn5 q4 qn5 RSTB VDD GND sg13g2_dfrbp_1
.ends
.end

** sch_path: xschem/top_13.sch
.subckt top_13 n_RO_control RO_control DUT_gate DUT_Footer DUT_Header Drain_Sense Drain_Force VDD VSS RSTB extra_load OUT
*.iopin n_RO_control
*.iopin RO_control
*.iopin DUT_gate
*.iopin DUT_Footer
*.iopin DUT_Header
*.iopin Drain_Sense
*.iopin Drain_Force
*.iopin VDD
*.iopin VSS
*.iopin RSTB
*.iopin extra_load
*.iopin OUT
x1 VDD VSS n_RO_control RO_control DUT_gate net1 DUT_Header DUT_Footer Drain_Force Drain_Sense extra_load top_RO_core_13
x2 VDD OUT net1 VSS RSTB div_sg13g2_stdcells
.ends

** sch_path: xschem/top_RO_core_101.sch
.subckt top_RO_core_101 VDD VSS n_RO_control RO_control DUT_gate Vout DUT_Header DUT_Footer Drain_Force Drain_Sense extra_load
*.iopin VDD
*.iopin VSS
*.iopin n_RO_control
*.iopin RO_control
*.iopin DUT_gate
*.iopin extra_load
*.iopin DUT_Header
*.iopin DUT_Footer
*.iopin Drain_Force
*.iopin Drain_Sense
*.iopin Vout
x1 VDD VSS A[97] A[96] rovcel2
x7 VDD VSS Vout A[100] rovcel2
x3[1] VDD VSS A[96] A[95] rovcel2
x3[2] VDD VSS A[95] A[94] rovcel2
x3[3] VDD VSS A[94] A[93] rovcel2
x3[4] VDD VSS A[93] A[92] rovcel2
x3[5] VDD VSS A[92] A[91] rovcel2
x3[6] VDD VSS A[91] A[90] rovcel2
x3[7] VDD VSS A[90] A[89] rovcel2
x3[8] VDD VSS A[89] A[88] rovcel2
x3[9] VDD VSS A[88] A[87] rovcel2
x3[10] VDD VSS A[87] A[86] rovcel2
x3[11] VDD VSS A[86] A[85] rovcel2
x3[12] VDD VSS A[85] A[84] rovcel2
x3[13] VDD VSS A[84] A[83] rovcel2
x3[14] VDD VSS A[83] A[82] rovcel2
x3[15] VDD VSS A[82] A[81] rovcel2
x3[16] VDD VSS A[81] A[80] rovcel2
x3[17] VDD VSS A[80] A[79] rovcel2
x3[18] VDD VSS A[79] A[78] rovcel2
x3[19] VDD VSS A[78] A[77] rovcel2
x3[20] VDD VSS A[77] A[76] rovcel2
x3[21] VDD VSS A[76] A[75] rovcel2
x3[22] VDD VSS A[75] A[74] rovcel2
x3[23] VDD VSS A[74] A[73] rovcel2
x3[24] VDD VSS A[73] A[72] rovcel2
x3[25] VDD VSS A[72] A[71] rovcel2
x3[26] VDD VSS A[71] A[70] rovcel2
x3[27] VDD VSS A[70] A[69] rovcel2
x3[28] VDD VSS A[69] A[68] rovcel2
x3[29] VDD VSS A[68] A[67] rovcel2
x3[30] VDD VSS A[67] A[66] rovcel2
x3[31] VDD VSS A[66] A[65] rovcel2
x3[32] VDD VSS A[65] A[64] rovcel2
x3[33] VDD VSS A[64] A[63] rovcel2
x3[34] VDD VSS A[63] A[62] rovcel2
x3[35] VDD VSS A[62] A[61] rovcel2
x3[36] VDD VSS A[61] A[60] rovcel2
x3[37] VDD VSS A[60] A[59] rovcel2
x3[38] VDD VSS A[59] A[58] rovcel2
x3[39] VDD VSS A[58] A[57] rovcel2
x3[40] VDD VSS A[57] A[56] rovcel2
x3[41] VDD VSS A[56] A[55] rovcel2
x3[42] VDD VSS A[55] A[54] rovcel2
x3[43] VDD VSS A[54] A[53] rovcel2
x3[44] VDD VSS A[53] A[52] rovcel2
x3[45] VDD VSS A[52] A[51] rovcel2
x3[46] VDD VSS A[51] A[50] rovcel2
x3[47] VDD VSS A[50] A[49] rovcel2
x3[48] VDD VSS A[49] A[48] rovcel2
x3[49] VDD VSS A[48] A[47] rovcel2
x3[50] VDD VSS A[47] A[46] rovcel2
x3[51] VDD VSS A[46] A[45] rovcel2
x3[52] VDD VSS A[45] A[44] rovcel2
x3[53] VDD VSS A[44] A[43] rovcel2
x3[54] VDD VSS A[43] A[42] rovcel2
x3[55] VDD VSS A[42] A[41] rovcel2
x3[56] VDD VSS A[41] A[40] rovcel2
x3[57] VDD VSS A[40] A[39] rovcel2
x3[58] VDD VSS A[39] A[38] rovcel2
x3[59] VDD VSS A[38] A[37] rovcel2
x3[60] VDD VSS A[37] A[36] rovcel2
x3[61] VDD VSS A[36] A[35] rovcel2
x3[62] VDD VSS A[35] A[34] rovcel2
x3[63] VDD VSS A[34] A[33] rovcel2
x3[64] VDD VSS A[33] A[32] rovcel2
x3[65] VDD VSS A[32] A[31] rovcel2
x3[66] VDD VSS A[31] A[30] rovcel2
x3[67] VDD VSS A[30] A[29] rovcel2
x3[68] VDD VSS A[29] A[28] rovcel2
x3[69] VDD VSS A[28] A[27] rovcel2
x3[70] VDD VSS A[27] A[26] rovcel2
x3[71] VDD VSS A[26] A[25] rovcel2
x3[72] VDD VSS A[25] A[24] rovcel2
x3[73] VDD VSS A[24] A[23] rovcel2
x3[74] VDD VSS A[23] A[22] rovcel2
x3[75] VDD VSS A[22] A[21] rovcel2
x3[76] VDD VSS A[21] A[20] rovcel2
x3[77] VDD VSS A[20] A[19] rovcel2
x3[78] VDD VSS A[19] A[18] rovcel2
x3[79] VDD VSS A[18] A[17] rovcel2
x3[80] VDD VSS A[17] A[16] rovcel2
x3[81] VDD VSS A[16] A[15] rovcel2
x3[82] VDD VSS A[15] A[14] rovcel2
x3[83] VDD VSS A[14] A[13] rovcel2
x3[84] VDD VSS A[13] A[12] rovcel2
x3[85] VDD VSS A[12] A[11] rovcel2
x3[86] VDD VSS A[11] A[10] rovcel2
x3[87] VDD VSS A[10] A[9] rovcel2
x3[88] VDD VSS A[9] A[8] rovcel2
x3[89] VDD VSS A[8] A[7] rovcel2
x3[90] VDD VSS A[7] A[6] rovcel2
x3[91] VDD VSS A[6] A[5] rovcel2
x3[92] VDD VSS A[5] A[4] rovcel2
x3[93] VDD VSS A[4] A[3] rovcel2
x3[94] VDD VSS A[3] A[2] rovcel2
x3[95] VDD VSS A[2] A[1] rovcel2
x3[96] VDD VSS A[1] Vout rovcel2
x3 VDD VSS A[97] n_RO_control A[98] RO_control DUT_gate rovcel3
x2 DUT_Header DUT_Footer Drain_Force Drain_Sense RO_control n_RO_control VDD VSS A[98] extra_load rovcel1
x4 VDD VSS extra_load n_RO_control A[100] rovcel4
.ends

** sch_path: xschem/top_101.sch
.subckt top_101 n_RO_control RO_control DUT_gate DUT_Footer DUT_Header Drain_Sense Drain_Force VDD VSS RSTB extra_load OUT
*.iopin n_RO_control
*.iopin RO_control
*.iopin DUT_gate
*.iopin DUT_Footer
*.iopin DUT_Header
*.iopin Drain_Sense
*.iopin Drain_Force
*.iopin VDD
*.iopin VSS
*.iopin RSTB
*.iopin extra_load
*.iopin OUT
x2 VDD OUT net1 VSS RSTB div_sg13g2_stdcells
x1 VDD VSS n_RO_control RO_control DUT_gate net1 DUT_Header DUT_Footer Drain_Force Drain_Sense extra_load top_RO_core_101
.ends
* CDL Netlist generated by OpenROAD

*.BUSDELIMITER [

.SUBCKT asicone_202508 AVDD RO2VDD ROVDD VDD VDDIO VSS VSSIO
+ pad_RO_101_DUT_gate_pad pad_RO_101_Drain_Force_pad pad_RO_101_Drain_Sense_pad
+ pad_RO_101_Vout_pad pad_RO_101_extra_load_pad pad_RO_13_DUT_gate_pad
+ pad_RO_13_Drain_Force_pad pad_RO_13_Drain_Sense_pad pad_RO_13_Vout_pad
+ pad_RO_13_extra_load_pad pad_RO_RST_B_pad pad_adc_clk_pad
+ pad_adc_go_pad pad_adc_result_0_pad pad_adc_result_1_pad pad_adc_result_2_pad
+ pad_adc_result_3_pad pad_adc_result_4_pad pad_adc_rst_pad
+ pad_adc_sample_pad pad_adc_valid_pad pad_adc_vin_pad pad_adc_vip_pad
+ pad_adc_vrefn_pad pad_adc_vrefp_pad pad_cs_pad pad_miso_pad
+ pad_mosi_pad pad_sclk_pad
XCORNER_1 VDDIO VSSIO VDD VSS VSS sg13g2_Corner
XCORNER_2 VDDIO VSSIO VDD VSS VSS sg13g2_Corner
XCORNER_3 VDDIO VSSIO VDD VSS VSS sg13g2_Corner
XCORNER_4 VDDIO VSSIO VDD VSS VSS sg13g2_Corner
XFILLER_0 VDDIO VSSIO VDD VSS VSS sg13g2_Filler4000
XFILLER_1 VDDIO VSSIO VDD VSS VSS sg13g2_Filler200
XFILLER_2 VDDIO VSSIO VDD VSS VSS sg13g2_Filler4000
XFILLER_3 VDDIO VSSIO VDD VSS VSS sg13g2_Filler200
XFILLER_4 VDDIO VSSIO VDD VSS VSS sg13g2_Filler4000
XFILLER_5 VDDIO VSSIO VDD VSS VSS sg13g2_Filler200
XFILLER_6 VDDIO VSSIO VDD VSS VSS sg13g2_Filler4000
XFILLER_7 VDDIO VSSIO VDD VSS VSS sg13g2_Filler200
Xadc AVDD pad_adc_clk_p2c pad_adc_go_p2c pad_adc_result_0_c2p
+ pad_adc_result_1_c2p pad_adc_result_2_c2p pad_adc_result_3_c2p
+ pad_adc_result_4_c2p pad_adc_rst_p2c pad_adc_sample_c2p pad_adc_valid_c2p
+ VDD pad_adc_vin_padres pad_adc_vip_padres pad_adc_vrefp_padres
+ pad_adc_vrefn_padres VSS SARADC
Xbd_pad_RO2_VDD sg13g2_bpd70
Xbd_pad_RO_101_DUT_gate sg13g2_bpd70
Xbd_pad_RO_101_Drain_Force sg13g2_bpd70
Xbd_pad_RO_101_Drain_Sense sg13g2_bpd70
Xbd_pad_RO_101_Vout sg13g2_bpd70
Xbd_pad_RO_101_extra_load sg13g2_bpd70
Xbd_pad_RO_13_DUT_gate sg13g2_bpd70
Xbd_pad_RO_13_Drain_Force sg13g2_bpd70
Xbd_pad_RO_13_Drain_Sense sg13g2_bpd70
Xbd_pad_RO_13_Vout sg13g2_bpd70
Xbd_pad_RO_13_extra_load sg13g2_bpd70
Xbd_pad_RO_RST_B sg13g2_bpd70
Xbd_pad_RO_VDD sg13g2_bpd70
Xbd_pad_RO_VSS sg13g2_bpd70
Xbd_pad_adc_avdd sg13g2_bpd70
Xbd_pad_adc_clk sg13g2_bpd70
Xbd_pad_adc_go sg13g2_bpd70
Xbd_pad_adc_result_0 sg13g2_bpd70
Xbd_pad_adc_result_1 sg13g2_bpd70
Xbd_pad_adc_result_2 sg13g2_bpd70
Xbd_pad_adc_result_3 sg13g2_bpd70
Xbd_pad_adc_result_4 sg13g2_bpd70
Xbd_pad_adc_rst sg13g2_bpd70
Xbd_pad_adc_sample sg13g2_bpd70
Xbd_pad_adc_valid sg13g2_bpd70
Xbd_pad_adc_vin sg13g2_bpd70
Xbd_pad_adc_vip sg13g2_bpd70
Xbd_pad_adc_vrefn sg13g2_bpd70
Xbd_pad_adc_vrefp sg13g2_bpd70
Xbd_pad_adc_vss sg13g2_bpd70
Xbd_pad_cs sg13g2_bpd70
Xbd_pad_miso sg13g2_bpd70
Xbd_pad_mosi sg13g2_bpd70
Xbd_pad_sclk sg13g2_bpd70
Xbd_vdd_north_0 sg13g2_bpd70
Xbd_vddpst_north_0 sg13g2_bpd70
Xbd_vss_north_0 sg13g2_bpd70
Xbd_vsspst_north_0 sg13g2_bpd70
Xbuf_spi_32 R[0] VDD VSS RD[32] sg13g2_BUFFD1
Xbuf_spi_33 R[1] VDD VSS RD[33] sg13g2_BUFFD1
Xbuf_spi_34 R[2] VDD VSS RD[34] sg13g2_BUFFD1
Xbuf_spi_35 R[3] VDD VSS RD[35] sg13g2_BUFFD1
Xbuf_spi_36 R[4] VDD VSS RD[36] sg13g2_BUFFD1
Xbuf_spi_37 R[5] VDD VSS RD[37] sg13g2_BUFFD1
Xbuf_spi_38 R[6] VDD VSS RD[38] sg13g2_BUFFD1
Xbuf_spi_39 R[7] VDD VSS RD[39] sg13g2_BUFFD1
Xbuf_spi_40 R[8] VDD VSS RD[40] sg13g2_BUFFD1
Xbuf_spi_41 R[9] VDD VSS RD[41] sg13g2_BUFFD1
Xbuf_spi_42 R[10] VDD VSS RD[42] sg13g2_BUFFD1
Xbuf_spi_43 R[11] VDD VSS RD[43] sg13g2_BUFFD1
Xbuf_spi_44 R[12] VDD VSS RD[44] sg13g2_BUFFD1
Xbuf_spi_45 R[13] VDD VSS RD[45] sg13g2_BUFFD1
Xbuf_spi_46 R[14] VDD VSS RD[46] sg13g2_BUFFD1
Xbuf_spi_47 R[15] VDD VSS RD[47] sg13g2_BUFFD1
Xpad_RO2_VDD VDDIO VSSIO RO2VDD pad_RO2_VDD_padres VDD VSS
+ VSS sg13g2_IOPadAnalog
Xpad_RO_101_DUT_gate VDDIO VSSIO pad_RO_101_DUT_gate_p2c pad_RO_101_DUT_gate_pad
+ VDD VSS VSS sg13g2_IOPadIn
Xpad_RO_101_Drain_Force VDDIO VSSIO pad_RO_101_Drain_Force_pad
+ pad_RO_101_Drain_Force_padres VDD VSS VSS sg13g2_IOPadAnalog
Xpad_RO_101_Drain_Sense VDDIO VSSIO pad_RO_101_Drain_Sense_pad
+ pad_RO_101_Drain_Sense_padres VDD VSS VSS sg13g2_IOPadAnalog
Xpad_RO_101_Vout pad_RO_101_Vout_c2p VDDIO VSSIO pad_RO_101_Vout_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_RO_101_extra_load VDDIO VSSIO pad_RO_101_extra_load_pad
+ pad_RO_101_extra_load_padres VDD VSS VSS sg13g2_IOPadAnalog
Xpad_RO_13_DUT_gate VDDIO VSSIO pad_RO_13_DUT_gate_p2c pad_RO_13_DUT_gate_pad
+ VDD VSS VSS sg13g2_IOPadIn
Xpad_RO_13_Drain_Force VDDIO VSSIO pad_RO_13_Drain_Force_pad
+ pad_RO_13_Drain_Force_padres VDD VSS VSS sg13g2_IOPadAnalog
Xpad_RO_13_Drain_Sense VDDIO VSSIO pad_RO_13_Drain_Sense_pad
+ pad_RO_13_Drain_Sense_padres VDD VSS VSS sg13g2_IOPadAnalog
Xpad_RO_13_Vout pad_RO_13_Vout_c2p VDDIO VSSIO pad_RO_13_Vout_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_RO_13_extra_load VDDIO VSSIO pad_RO_13_extra_load_pad
+ pad_RO_13_extra_load_padres VDD VSS VSS sg13g2_IOPadAnalog
Xpad_RO_RST_B VDDIO VSSIO pad_RO_RST_B_p2c pad_RO_RST_B_pad
+ VDD VSS VSS sg13g2_IOPadIn
Xpad_RO_VDD VDDIO VSSIO ROVDD pad_RO_VDD_padres VDD VSS VSS
+ sg13g2_IOPadAnalog
Xpad_RO_VSS VDDIO VSSIO VDD VSS VSS sg13g2_IOPadVssExt
Xpad_adc_avdd VDDIO VSSIO AVDD pad_adc_avdd_padres VDD VSS
+ VSS sg13g2_IOPadAnalog
Xpad_adc_clk VDDIO VSSIO pad_adc_clk_p2c pad_adc_clk_pad VDD
+ VSS VSS sg13g2_IOPadIn
Xpad_adc_go VDDIO VSSIO pad_adc_go_p2c pad_adc_go_pad VDD
+ VSS VSS sg13g2_IOPadIn
Xpad_adc_result_0 pad_adc_result_0_c2p VDDIO VSSIO pad_adc_result_0_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_result_1 pad_adc_result_1_c2p VDDIO VSSIO pad_adc_result_1_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_result_2 pad_adc_result_2_c2p VDDIO VSSIO pad_adc_result_2_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_result_3 pad_adc_result_3_c2p VDDIO VSSIO pad_adc_result_3_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_result_4 pad_adc_result_4_c2p VDDIO VSSIO pad_adc_result_4_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_rst VDDIO VSSIO pad_adc_rst_p2c pad_adc_rst_pad VDD
+ VSS VSS sg13g2_IOPadIn
Xpad_adc_sample pad_adc_sample_c2p VDDIO VSSIO pad_adc_sample_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_valid pad_adc_valid_c2p VDDIO VSSIO pad_adc_valid_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_vin VDDIO VSSIO pad_adc_vin_pad pad_adc_vin_padres
+ VDD VSS VSS sg13g2_IOPadAnalog
Xpad_adc_vip VDDIO VSSIO pad_adc_vip_pad pad_adc_vip_padres
+ VDD VSS VSS sg13g2_IOPadAnalog
Xpad_adc_vrefn VDDIO VSSIO pad_adc_vrefn_pad pad_adc_vrefn_padres
+ VDD VSS VSS sg13g2_IOPadAnalog
Xpad_adc_vrefp VDDIO VSSIO pad_adc_vrefp_pad pad_adc_vrefp_padres
+ VDD VSS VSS sg13g2_IOPadAnalog
Xpad_adc_vss VDDIO VSSIO VDD VSS VSS sg13g2_IOPadVssExt
Xpad_cs VDDIO VSSIO pad_cs_p2c pad_cs_pad VDD VSS VSS sg13g2_IOPadIn
Xpad_miso pad_miso_c2p VDDIO VSSIO pad_miso_pad VDD VSS VSS
+ sg13g2_IOPadOut16mA
Xpad_mosi VDDIO VSSIO pad_mosi_p2c pad_mosi_pad VDD VSS VSS
+ sg13g2_IOPadIn
Xpad_sclk VDDIO VSSIO pad_sclk_p2c pad_sclk_pad VDD VSS VSS
+ sg13g2_IOPadIn
Xpad_vdd_north_0 VDDIO VSSIO VDD VSS VSS sg13g2_IOPadVddExt
Xpad_vddpst_north_0 VDDIO VSSIO VDD VSS VSS sg13g2_IOPadIOVdd
Xpad_vss_north_0 VDDIO VSSIO VDD VSS VSS sg13g2_IOPadVssExt
Xpad_vsspst_north_0 VDDIO VSSIO VDD VSS VSS sg13g2_IOPadIOVss
Xro_101 R[0] R[1] pad_RO_101_DUT_gate_p2c R[2] R[3] pad_RO_101_Drain_Sense_padres
+ pad_RO_101_Drain_Force_padres ROVDD VSS pad_RO_RST_B_p2c pad_RO_101_extra_load_padres
+ pad_RO_101_Vout_c2p top_101
Xro_13 R[8] R[9] pad_RO_13_DUT_gate_p2c R[10] R[11] pad_RO_13_Drain_Sense_padres
+ pad_RO_13_Drain_Force_padres RO2VDD VSS pad_RO_RST_B_p2c pad_RO_13_extra_load_padres
+ pad_RO_13_Vout_c2p top_13
Xspi pad_cs_p2c pad_sclk_p2c pad_mosi_p2c pad_miso_c2p _unconnected_0
+ RD[0] RD[10] RD[11] RD[12] RD[13] RD[14] RD[15] RD[16] RD[17]
+ RD[18] RD[19] RD[1] RD[20] RD[21] RD[22] RD[23] RD[24] RD[25]
+ RD[26] RD[27] RD[28] RD[29] RD[2] RD[30] RD[31] RD[32] RD[33]
+ RD[34] RD[35] RD[36] RD[37] RD[38] RD[39] RD[3] RD[40] RD[41]
+ RD[42] RD[43] RD[44] RD[45] RD[46] RD[47] RD[4] RD[5] RD[6]
+ RD[7] RD[8] RD[9] pad_adc_rst_p2c R[0] R[10] R[11] R[12] R[13]
+ R[14] R[15] R[16] R[17] R[18] R[19] R[1] R[20] R[21] R[22]
+ R[23] R[24] R[25] R[26] R[27] R[28] R[29] R[2] R[30] R[31]
+ R[32] R[33] R[34] R[35] R[36] R[37] R[38] R[39] R[3] R[40]
+ R[41] R[42] R[43] R[44] R[45] R[46] R[47] R[48] R[49] R[4]
+ R[50] R[51] R[52] R[53] R[54] R[55] R[56] R[57] R[58] R[59]
+ R[5] R[60] R[61] R[62] R[63] R[6] R[7] R[8] R[9] VSS VDD SPI
Xspi_adc_result_0 RESULT[0] VDD VSS RD[0] sg13g2_BUFFD1
Xspi_adc_result_1 RESULT[1] VDD VSS RD[1] sg13g2_BUFFD1
Xspi_adc_result_2 RESULT[2] VDD VSS RD[2] sg13g2_BUFFD1
Xspi_adc_result_3 RESULT[3] VDD VSS RD[3] sg13g2_BUFFD1
Xspi_adc_result_4 RESULT[4] VDD VSS RD[4] sg13g2_BUFFD1
Xspi_adc_sample pad_adc_sample_c2p VDD VSS RD[9] sg13g2_BUFFD1
Xspi_adc_valid pad_adc_valid_c2p VDD VSS RD[8] sg13g2_BUFFD1
Xtie_spi_0 VDD VSS RD[5] sg13g2_TIEL
Xtie_spi_1 VDD VSS RD[6] sg13g2_TIEL
Xtie_spi_10 VDD VSS RD[10] sg13g2_TIEL
Xtie_spi_11 VDD VSS RD[11] sg13g2_TIEL
Xtie_spi_12 VDD VSS RD[12] sg13g2_TIEL
Xtie_spi_13 VDD VSS RD[13] sg13g2_TIEL
Xtie_spi_14 VDD VSS RD[14] sg13g2_TIEL
Xtie_spi_15 VDD VSS RD[15] sg13g2_TIEL
Xtie_spi_16 VDD VSS RD[16] sg13g2_TIEL
Xtie_spi_17 VDD VSS RD[17] sg13g2_TIEH
Xtie_spi_18 VDD VSS RD[18] sg13g2_TIEL
Xtie_spi_19 VDD VSS RD[19] sg13g2_TIEH
Xtie_spi_2 VDD VSS RD[7] sg13g2_TIEL
Xtie_spi_20 VDD VSS RD[20] sg13g2_TIEL
Xtie_spi_21 VDD VSS RD[21] sg13g2_TIEH
Xtie_spi_22 VDD VSS RD[22] sg13g2_TIEL
Xtie_spi_23 VDD VSS RD[23] sg13g2_TIEH
Xtie_spi_24 VDD VSS RD[24] sg13g2_TIEH
Xtie_spi_25 VDD VSS RD[25] sg13g2_TIEL
Xtie_spi_26 VDD VSS RD[26] sg13g2_TIEH
Xtie_spi_27 VDD VSS RD[27] sg13g2_TIEL
Xtie_spi_28 VDD VSS RD[28] sg13g2_TIEH
Xtie_spi_29 VDD VSS RD[29] sg13g2_TIEL
Xtie_spi_30 VDD VSS RD[30] sg13g2_TIEH
Xtie_spi_31 VDD VSS RD[31] sg13g2_TIEL
XANTENNA_1 pad_adc_sample_c2p VDD VSS sg13g2_ANTENNA
XANTENNA_2 pad_adc_sample_c2p VDD VSS sg13g2_ANTENNA
XSTDFILL0_0 VDD VSS sg13g2_FILL8
XSTDFILL0_8 VDD VSS sg13g2_FILL8
XSTDFILL0_16 VDD VSS sg13g2_FILL8
XSTDFILL0_24 VDD VSS sg13g2_FILL8
XSTDFILL0_32 VDD VSS sg13g2_FILL8
XSTDFILL0_40 VDD VSS sg13g2_FILL8
XSTDFILL0_48 VDD VSS sg13g2_FILL8
XSTDFILL0_56 VDD VSS sg13g2_FILL8
XSTDFILL0_64 VDD VSS sg13g2_FILL8
XSTDFILL0_72 VDD VSS sg13g2_FILL8
XSTDFILL0_80 VDD VSS sg13g2_FILL8
XSTDFILL0_88 VDD VSS sg13g2_FILL8
XSTDFILL0_96 VDD VSS sg13g2_FILL8
XSTDFILL0_104 VDD VSS sg13g2_FILL8
XSTDFILL0_112 VDD VSS sg13g2_FILL8
XSTDFILL0_120 VDD VSS sg13g2_FILL8
XSTDFILL0_128 VDD VSS sg13g2_FILL4
XSTDFILL0_1835 VDD VSS sg13g2_FILL8
XSTDFILL0_1843 VDD VSS sg13g2_FILL8
XSTDFILL0_1851 VDD VSS sg13g2_FILL8
XSTDFILL0_1859 VDD VSS sg13g2_FILL8
XSTDFILL0_1867 VDD VSS sg13g2_FILL8
XSTDFILL0_1875 VDD VSS sg13g2_FILL8
XSTDFILL0_1883 VDD VSS sg13g2_FILL8
XSTDFILL0_1891 VDD VSS sg13g2_FILL8
XSTDFILL0_1899 VDD VSS sg13g2_FILL8
XSTDFILL0_1907 VDD VSS sg13g2_FILL8
XSTDFILL0_1915 VDD VSS sg13g2_FILL8
XSTDFILL0_1923 VDD VSS sg13g2_FILL8
XSTDFILL0_1931 VDD VSS sg13g2_FILL8
XSTDFILL0_1939 VDD VSS sg13g2_FILL8
XSTDFILL0_1947 VDD VSS sg13g2_FILL8
XSTDFILL0_1955 VDD VSS sg13g2_FILL8
XSTDFILL0_1963 VDD VSS sg13g2_FILL8
XSTDFILL0_1971 VDD VSS sg13g2_FILL8
XSTDFILL0_1979 VDD VSS sg13g2_FILL8
XSTDFILL0_1987 VDD VSS sg13g2_FILL8
XSTDFILL0_1995 VDD VSS sg13g2_FILL8
XSTDFILL0_2003 VDD VSS sg13g2_FILL8
XSTDFILL0_2011 VDD VSS sg13g2_FILL8
XSTDFILL0_2019 VDD VSS sg13g2_FILL8
XSTDFILL0_2027 VDD VSS sg13g2_FILL8
XSTDFILL0_2035 VDD VSS sg13g2_FILL8
XSTDFILL0_2043 VDD VSS sg13g2_FILL8
XSTDFILL0_2051 VDD VSS sg13g2_FILL8
XSTDFILL0_2059 VDD VSS sg13g2_FILL8
XSTDFILL0_2067 VDD VSS sg13g2_FILL8
XSTDFILL0_2075 VDD VSS sg13g2_FILL8
XSTDFILL0_2083 VDD VSS sg13g2_FILL8
XSTDFILL0_2091 VDD VSS sg13g2_FILL8
XSTDFILL0_2099 VDD VSS sg13g2_FILL8
XSTDFILL0_2107 VDD VSS sg13g2_FILL8
XSTDFILL0_2115 VDD VSS sg13g2_FILL8
XSTDFILL0_2123 VDD VSS sg13g2_FILL8
XSTDFILL0_2131 VDD VSS sg13g2_FILL8
XSTDFILL0_2139 VDD VSS sg13g2_FILL8
XSTDFILL0_2147 VDD VSS sg13g2_FILL4
XSTDFILL0_2151 VDD VSS sg13g2_FILL2
XSTDFILL0_2153 VDD VSS sg13g2_FILL1
XSTDFILL1_0 VDD VSS sg13g2_FILL8
XSTDFILL1_8 VDD VSS sg13g2_FILL8
XSTDFILL1_16 VDD VSS sg13g2_FILL8
XSTDFILL1_24 VDD VSS sg13g2_FILL8
XSTDFILL1_32 VDD VSS sg13g2_FILL8
XSTDFILL1_40 VDD VSS sg13g2_FILL8
XSTDFILL1_48 VDD VSS sg13g2_FILL8
XSTDFILL1_56 VDD VSS sg13g2_FILL8
XSTDFILL1_64 VDD VSS sg13g2_FILL8
XSTDFILL1_72 VDD VSS sg13g2_FILL8
XSTDFILL1_80 VDD VSS sg13g2_FILL8
XSTDFILL1_88 VDD VSS sg13g2_FILL8
XSTDFILL1_96 VDD VSS sg13g2_FILL8
XSTDFILL1_104 VDD VSS sg13g2_FILL8
XSTDFILL1_112 VDD VSS sg13g2_FILL8
XSTDFILL1_120 VDD VSS sg13g2_FILL8
XSTDFILL1_128 VDD VSS sg13g2_FILL4
XSTDFILL1_1835 VDD VSS sg13g2_FILL8
XSTDFILL1_1843 VDD VSS sg13g2_FILL8
XSTDFILL1_1851 VDD VSS sg13g2_FILL8
XSTDFILL1_1859 VDD VSS sg13g2_FILL8
XSTDFILL1_1867 VDD VSS sg13g2_FILL8
XSTDFILL1_1875 VDD VSS sg13g2_FILL8
XSTDFILL1_1883 VDD VSS sg13g2_FILL8
XSTDFILL1_1891 VDD VSS sg13g2_FILL8
XSTDFILL1_1899 VDD VSS sg13g2_FILL8
XSTDFILL1_1907 VDD VSS sg13g2_FILL8
XSTDFILL1_1915 VDD VSS sg13g2_FILL8
XSTDFILL1_1923 VDD VSS sg13g2_FILL8
XSTDFILL1_1931 VDD VSS sg13g2_FILL8
XSTDFILL1_1939 VDD VSS sg13g2_FILL8
XSTDFILL1_1947 VDD VSS sg13g2_FILL8
XSTDFILL1_1955 VDD VSS sg13g2_FILL8
XSTDFILL1_1963 VDD VSS sg13g2_FILL8
XSTDFILL1_1971 VDD VSS sg13g2_FILL8
XSTDFILL1_1979 VDD VSS sg13g2_FILL8
XSTDFILL1_1987 VDD VSS sg13g2_FILL8
XSTDFILL1_1995 VDD VSS sg13g2_FILL8
XSTDFILL1_2003 VDD VSS sg13g2_FILL8
XSTDFILL1_2011 VDD VSS sg13g2_FILL8
XSTDFILL1_2019 VDD VSS sg13g2_FILL8
XSTDFILL1_2027 VDD VSS sg13g2_FILL8
XSTDFILL1_2035 VDD VSS sg13g2_FILL8
XSTDFILL1_2043 VDD VSS sg13g2_FILL8
XSTDFILL1_2051 VDD VSS sg13g2_FILL8
XSTDFILL1_2059 VDD VSS sg13g2_FILL8
XSTDFILL1_2067 VDD VSS sg13g2_FILL8
XSTDFILL1_2075 VDD VSS sg13g2_FILL8
XSTDFILL1_2083 VDD VSS sg13g2_FILL8
XSTDFILL1_2091 VDD VSS sg13g2_FILL8
XSTDFILL1_2099 VDD VSS sg13g2_FILL8
XSTDFILL1_2107 VDD VSS sg13g2_FILL8
XSTDFILL1_2115 VDD VSS sg13g2_FILL8
XSTDFILL1_2123 VDD VSS sg13g2_FILL8
XSTDFILL1_2131 VDD VSS sg13g2_FILL8
XSTDFILL1_2139 VDD VSS sg13g2_FILL8
XSTDFILL1_2147 VDD VSS sg13g2_FILL4
XSTDFILL1_2151 VDD VSS sg13g2_FILL2
XSTDFILL1_2153 VDD VSS sg13g2_FILL1
XSTDFILL2_0 VDD VSS sg13g2_FILL8
XSTDFILL2_8 VDD VSS sg13g2_FILL8
XSTDFILL2_16 VDD VSS sg13g2_FILL8
XSTDFILL2_24 VDD VSS sg13g2_FILL8
XSTDFILL2_32 VDD VSS sg13g2_FILL8
XSTDFILL2_40 VDD VSS sg13g2_FILL8
XSTDFILL2_48 VDD VSS sg13g2_FILL8
XSTDFILL2_56 VDD VSS sg13g2_FILL8
XSTDFILL2_64 VDD VSS sg13g2_FILL8
XSTDFILL2_72 VDD VSS sg13g2_FILL8
XSTDFILL2_80 VDD VSS sg13g2_FILL8
XSTDFILL2_88 VDD VSS sg13g2_FILL8
XSTDFILL2_96 VDD VSS sg13g2_FILL8
XSTDFILL2_104 VDD VSS sg13g2_FILL8
XSTDFILL2_112 VDD VSS sg13g2_FILL8
XSTDFILL2_120 VDD VSS sg13g2_FILL8
XSTDFILL2_128 VDD VSS sg13g2_FILL4
XSTDFILL2_1835 VDD VSS sg13g2_FILL8
XSTDFILL2_1843 VDD VSS sg13g2_FILL8
XSTDFILL2_1851 VDD VSS sg13g2_FILL8
XSTDFILL2_1859 VDD VSS sg13g2_FILL8
XSTDFILL2_1867 VDD VSS sg13g2_FILL8
XSTDFILL2_1875 VDD VSS sg13g2_FILL8
XSTDFILL2_1883 VDD VSS sg13g2_FILL8
XSTDFILL2_1891 VDD VSS sg13g2_FILL8
XSTDFILL2_1899 VDD VSS sg13g2_FILL8
XSTDFILL2_1907 VDD VSS sg13g2_FILL8
XSTDFILL2_1915 VDD VSS sg13g2_FILL8
XSTDFILL2_1923 VDD VSS sg13g2_FILL8
XSTDFILL2_1931 VDD VSS sg13g2_FILL8
XSTDFILL2_1939 VDD VSS sg13g2_FILL8
XSTDFILL2_1947 VDD VSS sg13g2_FILL8
XSTDFILL2_1955 VDD VSS sg13g2_FILL8
XSTDFILL2_1963 VDD VSS sg13g2_FILL8
XSTDFILL2_1971 VDD VSS sg13g2_FILL8
XSTDFILL2_1979 VDD VSS sg13g2_FILL8
XSTDFILL2_1987 VDD VSS sg13g2_FILL8
XSTDFILL2_1995 VDD VSS sg13g2_FILL8
XSTDFILL2_2003 VDD VSS sg13g2_FILL8
XSTDFILL2_2011 VDD VSS sg13g2_FILL8
XSTDFILL2_2019 VDD VSS sg13g2_FILL8
XSTDFILL2_2027 VDD VSS sg13g2_FILL8
XSTDFILL2_2035 VDD VSS sg13g2_FILL8
XSTDFILL2_2043 VDD VSS sg13g2_FILL8
XSTDFILL2_2051 VDD VSS sg13g2_FILL8
XSTDFILL2_2059 VDD VSS sg13g2_FILL8
XSTDFILL2_2067 VDD VSS sg13g2_FILL8
XSTDFILL2_2075 VDD VSS sg13g2_FILL8
XSTDFILL2_2083 VDD VSS sg13g2_FILL8
XSTDFILL2_2091 VDD VSS sg13g2_FILL8
XSTDFILL2_2099 VDD VSS sg13g2_FILL8
XSTDFILL2_2107 VDD VSS sg13g2_FILL8
XSTDFILL2_2115 VDD VSS sg13g2_FILL8
XSTDFILL2_2123 VDD VSS sg13g2_FILL8
XSTDFILL2_2131 VDD VSS sg13g2_FILL8
XSTDFILL2_2139 VDD VSS sg13g2_FILL8
XSTDFILL2_2147 VDD VSS sg13g2_FILL4
XSTDFILL2_2151 VDD VSS sg13g2_FILL2
XSTDFILL2_2153 VDD VSS sg13g2_FILL1
XSTDFILL3_0 VDD VSS sg13g2_FILL8
XSTDFILL3_8 VDD VSS sg13g2_FILL8
XSTDFILL3_16 VDD VSS sg13g2_FILL8
XSTDFILL3_24 VDD VSS sg13g2_FILL8
XSTDFILL3_32 VDD VSS sg13g2_FILL8
XSTDFILL3_40 VDD VSS sg13g2_FILL8
XSTDFILL3_48 VDD VSS sg13g2_FILL8
XSTDFILL3_56 VDD VSS sg13g2_FILL8
XSTDFILL3_64 VDD VSS sg13g2_FILL8
XSTDFILL3_72 VDD VSS sg13g2_FILL8
XSTDFILL3_80 VDD VSS sg13g2_FILL8
XSTDFILL3_88 VDD VSS sg13g2_FILL8
XSTDFILL3_96 VDD VSS sg13g2_FILL8
XSTDFILL3_104 VDD VSS sg13g2_FILL8
XSTDFILL3_112 VDD VSS sg13g2_FILL8
XSTDFILL3_120 VDD VSS sg13g2_FILL8
XSTDFILL3_128 VDD VSS sg13g2_FILL4
XSTDFILL3_1835 VDD VSS sg13g2_FILL8
XSTDFILL3_1843 VDD VSS sg13g2_FILL8
XSTDFILL3_1851 VDD VSS sg13g2_FILL8
XSTDFILL3_1859 VDD VSS sg13g2_FILL8
XSTDFILL3_1867 VDD VSS sg13g2_FILL8
XSTDFILL3_1875 VDD VSS sg13g2_FILL8
XSTDFILL3_1883 VDD VSS sg13g2_FILL8
XSTDFILL3_1891 VDD VSS sg13g2_FILL8
XSTDFILL3_1899 VDD VSS sg13g2_FILL8
XSTDFILL3_1907 VDD VSS sg13g2_FILL8
XSTDFILL3_1915 VDD VSS sg13g2_FILL8
XSTDFILL3_1923 VDD VSS sg13g2_FILL8
XSTDFILL3_1931 VDD VSS sg13g2_FILL8
XSTDFILL3_1939 VDD VSS sg13g2_FILL8
XSTDFILL3_1947 VDD VSS sg13g2_FILL8
XSTDFILL3_1955 VDD VSS sg13g2_FILL8
XSTDFILL3_1963 VDD VSS sg13g2_FILL8
XSTDFILL3_1971 VDD VSS sg13g2_FILL8
XSTDFILL3_1979 VDD VSS sg13g2_FILL8
XSTDFILL3_1987 VDD VSS sg13g2_FILL8
XSTDFILL3_1995 VDD VSS sg13g2_FILL8
XSTDFILL3_2003 VDD VSS sg13g2_FILL8
XSTDFILL3_2011 VDD VSS sg13g2_FILL8
XSTDFILL3_2019 VDD VSS sg13g2_FILL8
XSTDFILL3_2027 VDD VSS sg13g2_FILL8
XSTDFILL3_2035 VDD VSS sg13g2_FILL8
XSTDFILL3_2043 VDD VSS sg13g2_FILL8
XSTDFILL3_2051 VDD VSS sg13g2_FILL8
XSTDFILL3_2059 VDD VSS sg13g2_FILL8
XSTDFILL3_2067 VDD VSS sg13g2_FILL8
XSTDFILL3_2075 VDD VSS sg13g2_FILL8
XSTDFILL3_2083 VDD VSS sg13g2_FILL8
XSTDFILL3_2091 VDD VSS sg13g2_FILL8
XSTDFILL3_2099 VDD VSS sg13g2_FILL8
XSTDFILL3_2107 VDD VSS sg13g2_FILL8
XSTDFILL3_2115 VDD VSS sg13g2_FILL8
XSTDFILL3_2123 VDD VSS sg13g2_FILL8
XSTDFILL3_2131 VDD VSS sg13g2_FILL8
XSTDFILL3_2139 VDD VSS sg13g2_FILL8
XSTDFILL3_2147 VDD VSS sg13g2_FILL4
XSTDFILL3_2151 VDD VSS sg13g2_FILL2
XSTDFILL3_2153 VDD VSS sg13g2_FILL1
XSTDFILL4_0 VDD VSS sg13g2_FILL8
XSTDFILL4_8 VDD VSS sg13g2_FILL8
XSTDFILL4_16 VDD VSS sg13g2_FILL8
XSTDFILL4_24 VDD VSS sg13g2_FILL8
XSTDFILL4_32 VDD VSS sg13g2_FILL8
XSTDFILL4_40 VDD VSS sg13g2_FILL8
XSTDFILL4_48 VDD VSS sg13g2_FILL8
XSTDFILL4_56 VDD VSS sg13g2_FILL8
XSTDFILL4_64 VDD VSS sg13g2_FILL8
XSTDFILL4_72 VDD VSS sg13g2_FILL8
XSTDFILL4_80 VDD VSS sg13g2_FILL8
XSTDFILL4_88 VDD VSS sg13g2_FILL8
XSTDFILL4_96 VDD VSS sg13g2_FILL8
XSTDFILL4_104 VDD VSS sg13g2_FILL8
XSTDFILL4_112 VDD VSS sg13g2_FILL8
XSTDFILL4_120 VDD VSS sg13g2_FILL8
XSTDFILL4_128 VDD VSS sg13g2_FILL4
XSTDFILL4_1835 VDD VSS sg13g2_FILL8
XSTDFILL4_1843 VDD VSS sg13g2_FILL8
XSTDFILL4_1851 VDD VSS sg13g2_FILL8
XSTDFILL4_1859 VDD VSS sg13g2_FILL8
XSTDFILL4_1867 VDD VSS sg13g2_FILL8
XSTDFILL4_1875 VDD VSS sg13g2_FILL8
XSTDFILL4_1883 VDD VSS sg13g2_FILL8
XSTDFILL4_1891 VDD VSS sg13g2_FILL8
XSTDFILL4_1899 VDD VSS sg13g2_FILL8
XSTDFILL4_1907 VDD VSS sg13g2_FILL8
XSTDFILL4_1915 VDD VSS sg13g2_FILL8
XSTDFILL4_1923 VDD VSS sg13g2_FILL8
XSTDFILL4_1931 VDD VSS sg13g2_FILL8
XSTDFILL4_1939 VDD VSS sg13g2_FILL8
XSTDFILL4_1947 VDD VSS sg13g2_FILL8
XSTDFILL4_1955 VDD VSS sg13g2_FILL8
XSTDFILL4_1963 VDD VSS sg13g2_FILL8
XSTDFILL4_1971 VDD VSS sg13g2_FILL8
XSTDFILL4_1979 VDD VSS sg13g2_FILL8
XSTDFILL4_1987 VDD VSS sg13g2_FILL8
XSTDFILL4_1995 VDD VSS sg13g2_FILL8
XSTDFILL4_2003 VDD VSS sg13g2_FILL8
XSTDFILL4_2011 VDD VSS sg13g2_FILL8
XSTDFILL4_2019 VDD VSS sg13g2_FILL8
XSTDFILL4_2027 VDD VSS sg13g2_FILL8
XSTDFILL4_2035 VDD VSS sg13g2_FILL8
XSTDFILL4_2043 VDD VSS sg13g2_FILL8
XSTDFILL4_2051 VDD VSS sg13g2_FILL8
XSTDFILL4_2059 VDD VSS sg13g2_FILL8
XSTDFILL4_2067 VDD VSS sg13g2_FILL8
XSTDFILL4_2075 VDD VSS sg13g2_FILL8
XSTDFILL4_2083 VDD VSS sg13g2_FILL8
XSTDFILL4_2091 VDD VSS sg13g2_FILL8
XSTDFILL4_2099 VDD VSS sg13g2_FILL8
XSTDFILL4_2107 VDD VSS sg13g2_FILL8
XSTDFILL4_2115 VDD VSS sg13g2_FILL8
XSTDFILL4_2123 VDD VSS sg13g2_FILL8
XSTDFILL4_2131 VDD VSS sg13g2_FILL8
XSTDFILL4_2139 VDD VSS sg13g2_FILL8
XSTDFILL4_2147 VDD VSS sg13g2_FILL4
XSTDFILL4_2151 VDD VSS sg13g2_FILL2
XSTDFILL4_2153 VDD VSS sg13g2_FILL1
XSTDFILL5_0 VDD VSS sg13g2_FILL8
XSTDFILL5_8 VDD VSS sg13g2_FILL8
XSTDFILL5_16 VDD VSS sg13g2_FILL8
XSTDFILL5_24 VDD VSS sg13g2_FILL8
XSTDFILL5_32 VDD VSS sg13g2_FILL8
XSTDFILL5_40 VDD VSS sg13g2_FILL8
XSTDFILL5_48 VDD VSS sg13g2_FILL8
XSTDFILL5_56 VDD VSS sg13g2_FILL8
XSTDFILL5_64 VDD VSS sg13g2_FILL8
XSTDFILL5_72 VDD VSS sg13g2_FILL8
XSTDFILL5_80 VDD VSS sg13g2_FILL8
XSTDFILL5_88 VDD VSS sg13g2_FILL8
XSTDFILL5_96 VDD VSS sg13g2_FILL8
XSTDFILL5_104 VDD VSS sg13g2_FILL8
XSTDFILL5_112 VDD VSS sg13g2_FILL8
XSTDFILL5_120 VDD VSS sg13g2_FILL8
XSTDFILL5_128 VDD VSS sg13g2_FILL4
XSTDFILL5_1835 VDD VSS sg13g2_FILL8
XSTDFILL5_1843 VDD VSS sg13g2_FILL8
XSTDFILL5_1851 VDD VSS sg13g2_FILL8
XSTDFILL5_1859 VDD VSS sg13g2_FILL8
XSTDFILL5_1867 VDD VSS sg13g2_FILL8
XSTDFILL5_1875 VDD VSS sg13g2_FILL8
XSTDFILL5_1883 VDD VSS sg13g2_FILL8
XSTDFILL5_1891 VDD VSS sg13g2_FILL8
XSTDFILL5_1899 VDD VSS sg13g2_FILL8
XSTDFILL5_1907 VDD VSS sg13g2_FILL8
XSTDFILL5_1915 VDD VSS sg13g2_FILL8
XSTDFILL5_1923 VDD VSS sg13g2_FILL8
XSTDFILL5_1931 VDD VSS sg13g2_FILL8
XSTDFILL5_1939 VDD VSS sg13g2_FILL8
XSTDFILL5_1947 VDD VSS sg13g2_FILL8
XSTDFILL5_1955 VDD VSS sg13g2_FILL8
XSTDFILL5_1963 VDD VSS sg13g2_FILL8
XSTDFILL5_1971 VDD VSS sg13g2_FILL8
XSTDFILL5_1979 VDD VSS sg13g2_FILL8
XSTDFILL5_1987 VDD VSS sg13g2_FILL8
XSTDFILL5_1995 VDD VSS sg13g2_FILL8
XSTDFILL5_2003 VDD VSS sg13g2_FILL8
XSTDFILL5_2011 VDD VSS sg13g2_FILL8
XSTDFILL5_2019 VDD VSS sg13g2_FILL8
XSTDFILL5_2027 VDD VSS sg13g2_FILL8
XSTDFILL5_2035 VDD VSS sg13g2_FILL8
XSTDFILL5_2043 VDD VSS sg13g2_FILL8
XSTDFILL5_2051 VDD VSS sg13g2_FILL8
XSTDFILL5_2059 VDD VSS sg13g2_FILL8
XSTDFILL5_2067 VDD VSS sg13g2_FILL8
XSTDFILL5_2075 VDD VSS sg13g2_FILL8
XSTDFILL5_2083 VDD VSS sg13g2_FILL8
XSTDFILL5_2091 VDD VSS sg13g2_FILL8
XSTDFILL5_2099 VDD VSS sg13g2_FILL8
XSTDFILL5_2107 VDD VSS sg13g2_FILL8
XSTDFILL5_2115 VDD VSS sg13g2_FILL8
XSTDFILL5_2123 VDD VSS sg13g2_FILL8
XSTDFILL5_2131 VDD VSS sg13g2_FILL8
XSTDFILL5_2139 VDD VSS sg13g2_FILL8
XSTDFILL5_2147 VDD VSS sg13g2_FILL4
XSTDFILL5_2151 VDD VSS sg13g2_FILL2
XSTDFILL5_2153 VDD VSS sg13g2_FILL1
XSTDFILL6_0 VDD VSS sg13g2_FILL8
XSTDFILL6_8 VDD VSS sg13g2_FILL8
XSTDFILL6_16 VDD VSS sg13g2_FILL8
XSTDFILL6_24 VDD VSS sg13g2_FILL8
XSTDFILL6_32 VDD VSS sg13g2_FILL8
XSTDFILL6_40 VDD VSS sg13g2_FILL8
XSTDFILL6_48 VDD VSS sg13g2_FILL8
XSTDFILL6_56 VDD VSS sg13g2_FILL8
XSTDFILL6_64 VDD VSS sg13g2_FILL8
XSTDFILL6_72 VDD VSS sg13g2_FILL8
XSTDFILL6_80 VDD VSS sg13g2_FILL8
XSTDFILL6_88 VDD VSS sg13g2_FILL8
XSTDFILL6_96 VDD VSS sg13g2_FILL8
XSTDFILL6_104 VDD VSS sg13g2_FILL8
XSTDFILL6_112 VDD VSS sg13g2_FILL8
XSTDFILL6_120 VDD VSS sg13g2_FILL8
XSTDFILL6_128 VDD VSS sg13g2_FILL4
XSTDFILL6_1835 VDD VSS sg13g2_FILL8
XSTDFILL6_1843 VDD VSS sg13g2_FILL8
XSTDFILL6_1851 VDD VSS sg13g2_FILL8
XSTDFILL6_1859 VDD VSS sg13g2_FILL8
XSTDFILL6_1867 VDD VSS sg13g2_FILL8
XSTDFILL6_1875 VDD VSS sg13g2_FILL8
XSTDFILL6_1883 VDD VSS sg13g2_FILL8
XSTDFILL6_1891 VDD VSS sg13g2_FILL8
XSTDFILL6_1899 VDD VSS sg13g2_FILL8
XSTDFILL6_1907 VDD VSS sg13g2_FILL8
XSTDFILL6_1915 VDD VSS sg13g2_FILL8
XSTDFILL6_1923 VDD VSS sg13g2_FILL8
XSTDFILL6_1931 VDD VSS sg13g2_FILL8
XSTDFILL6_1939 VDD VSS sg13g2_FILL8
XSTDFILL6_1947 VDD VSS sg13g2_FILL8
XSTDFILL6_1955 VDD VSS sg13g2_FILL8
XSTDFILL6_1963 VDD VSS sg13g2_FILL8
XSTDFILL6_1971 VDD VSS sg13g2_FILL8
XSTDFILL6_1979 VDD VSS sg13g2_FILL8
XSTDFILL6_1987 VDD VSS sg13g2_FILL8
XSTDFILL6_1995 VDD VSS sg13g2_FILL8
XSTDFILL6_2003 VDD VSS sg13g2_FILL8
XSTDFILL6_2011 VDD VSS sg13g2_FILL8
XSTDFILL6_2019 VDD VSS sg13g2_FILL8
XSTDFILL6_2027 VDD VSS sg13g2_FILL8
XSTDFILL6_2035 VDD VSS sg13g2_FILL8
XSTDFILL6_2043 VDD VSS sg13g2_FILL8
XSTDFILL6_2051 VDD VSS sg13g2_FILL8
XSTDFILL6_2059 VDD VSS sg13g2_FILL8
XSTDFILL6_2067 VDD VSS sg13g2_FILL8
XSTDFILL6_2075 VDD VSS sg13g2_FILL8
XSTDFILL6_2083 VDD VSS sg13g2_FILL8
XSTDFILL6_2091 VDD VSS sg13g2_FILL8
XSTDFILL6_2099 VDD VSS sg13g2_FILL8
XSTDFILL6_2107 VDD VSS sg13g2_FILL8
XSTDFILL6_2115 VDD VSS sg13g2_FILL8
XSTDFILL6_2123 VDD VSS sg13g2_FILL8
XSTDFILL6_2131 VDD VSS sg13g2_FILL8
XSTDFILL6_2139 VDD VSS sg13g2_FILL8
XSTDFILL6_2147 VDD VSS sg13g2_FILL4
XSTDFILL6_2151 VDD VSS sg13g2_FILL2
XSTDFILL6_2153 VDD VSS sg13g2_FILL1
XSTDFILL7_0 VDD VSS sg13g2_FILL8
XSTDFILL7_8 VDD VSS sg13g2_FILL8
XSTDFILL7_16 VDD VSS sg13g2_FILL8
XSTDFILL7_24 VDD VSS sg13g2_FILL8
XSTDFILL7_32 VDD VSS sg13g2_FILL8
XSTDFILL7_40 VDD VSS sg13g2_FILL8
XSTDFILL7_48 VDD VSS sg13g2_FILL8
XSTDFILL7_56 VDD VSS sg13g2_FILL8
XSTDFILL7_64 VDD VSS sg13g2_FILL8
XSTDFILL7_72 VDD VSS sg13g2_FILL8
XSTDFILL7_80 VDD VSS sg13g2_FILL8
XSTDFILL7_88 VDD VSS sg13g2_FILL8
XSTDFILL7_96 VDD VSS sg13g2_FILL8
XSTDFILL7_104 VDD VSS sg13g2_FILL8
XSTDFILL7_112 VDD VSS sg13g2_FILL8
XSTDFILL7_120 VDD VSS sg13g2_FILL8
XSTDFILL7_128 VDD VSS sg13g2_FILL4
XSTDFILL7_1835 VDD VSS sg13g2_FILL8
XSTDFILL7_1843 VDD VSS sg13g2_FILL8
XSTDFILL7_1851 VDD VSS sg13g2_FILL8
XSTDFILL7_1859 VDD VSS sg13g2_FILL8
XSTDFILL7_1867 VDD VSS sg13g2_FILL8
XSTDFILL7_1875 VDD VSS sg13g2_FILL8
XSTDFILL7_1883 VDD VSS sg13g2_FILL8
XSTDFILL7_1891 VDD VSS sg13g2_FILL8
XSTDFILL7_1899 VDD VSS sg13g2_FILL8
XSTDFILL7_1907 VDD VSS sg13g2_FILL8
XSTDFILL7_1915 VDD VSS sg13g2_FILL8
XSTDFILL7_1923 VDD VSS sg13g2_FILL8
XSTDFILL7_1931 VDD VSS sg13g2_FILL8
XSTDFILL7_1939 VDD VSS sg13g2_FILL8
XSTDFILL7_1947 VDD VSS sg13g2_FILL8
XSTDFILL7_1955 VDD VSS sg13g2_FILL8
XSTDFILL7_1963 VDD VSS sg13g2_FILL8
XSTDFILL7_1971 VDD VSS sg13g2_FILL8
XSTDFILL7_1979 VDD VSS sg13g2_FILL8
XSTDFILL7_1987 VDD VSS sg13g2_FILL8
XSTDFILL7_1995 VDD VSS sg13g2_FILL8
XSTDFILL7_2003 VDD VSS sg13g2_FILL8
XSTDFILL7_2011 VDD VSS sg13g2_FILL8
XSTDFILL7_2019 VDD VSS sg13g2_FILL8
XSTDFILL7_2027 VDD VSS sg13g2_FILL8
XSTDFILL7_2035 VDD VSS sg13g2_FILL8
XSTDFILL7_2043 VDD VSS sg13g2_FILL8
XSTDFILL7_2051 VDD VSS sg13g2_FILL8
XSTDFILL7_2059 VDD VSS sg13g2_FILL8
XSTDFILL7_2067 VDD VSS sg13g2_FILL8
XSTDFILL7_2075 VDD VSS sg13g2_FILL8
XSTDFILL7_2083 VDD VSS sg13g2_FILL8
XSTDFILL7_2091 VDD VSS sg13g2_FILL8
XSTDFILL7_2099 VDD VSS sg13g2_FILL8
XSTDFILL7_2107 VDD VSS sg13g2_FILL8
XSTDFILL7_2115 VDD VSS sg13g2_FILL8
XSTDFILL7_2123 VDD VSS sg13g2_FILL8
XSTDFILL7_2131 VDD VSS sg13g2_FILL8
XSTDFILL7_2139 VDD VSS sg13g2_FILL8
XSTDFILL7_2147 VDD VSS sg13g2_FILL4
XSTDFILL7_2151 VDD VSS sg13g2_FILL2
XSTDFILL7_2153 VDD VSS sg13g2_FILL1
XSTDFILL8_0 VDD VSS sg13g2_FILL8
XSTDFILL8_8 VDD VSS sg13g2_FILL8
XSTDFILL8_16 VDD VSS sg13g2_FILL8
XSTDFILL8_24 VDD VSS sg13g2_FILL8
XSTDFILL8_32 VDD VSS sg13g2_FILL8
XSTDFILL8_40 VDD VSS sg13g2_FILL8
XSTDFILL8_48 VDD VSS sg13g2_FILL8
XSTDFILL8_56 VDD VSS sg13g2_FILL8
XSTDFILL8_64 VDD VSS sg13g2_FILL8
XSTDFILL8_72 VDD VSS sg13g2_FILL8
XSTDFILL8_80 VDD VSS sg13g2_FILL8
XSTDFILL8_88 VDD VSS sg13g2_FILL8
XSTDFILL8_96 VDD VSS sg13g2_FILL8
XSTDFILL8_104 VDD VSS sg13g2_FILL8
XSTDFILL8_112 VDD VSS sg13g2_FILL8
XSTDFILL8_120 VDD VSS sg13g2_FILL8
XSTDFILL8_128 VDD VSS sg13g2_FILL4
XSTDFILL8_1835 VDD VSS sg13g2_FILL8
XSTDFILL8_1843 VDD VSS sg13g2_FILL8
XSTDFILL8_1851 VDD VSS sg13g2_FILL8
XSTDFILL8_1859 VDD VSS sg13g2_FILL8
XSTDFILL8_1867 VDD VSS sg13g2_FILL8
XSTDFILL8_1875 VDD VSS sg13g2_FILL8
XSTDFILL8_1883 VDD VSS sg13g2_FILL8
XSTDFILL8_1891 VDD VSS sg13g2_FILL8
XSTDFILL8_1899 VDD VSS sg13g2_FILL8
XSTDFILL8_1907 VDD VSS sg13g2_FILL8
XSTDFILL8_1915 VDD VSS sg13g2_FILL8
XSTDFILL8_1923 VDD VSS sg13g2_FILL8
XSTDFILL8_1931 VDD VSS sg13g2_FILL8
XSTDFILL8_1939 VDD VSS sg13g2_FILL8
XSTDFILL8_1947 VDD VSS sg13g2_FILL8
XSTDFILL8_1955 VDD VSS sg13g2_FILL8
XSTDFILL8_1963 VDD VSS sg13g2_FILL8
XSTDFILL8_1971 VDD VSS sg13g2_FILL8
XSTDFILL8_1979 VDD VSS sg13g2_FILL8
XSTDFILL8_1987 VDD VSS sg13g2_FILL8
XSTDFILL8_1995 VDD VSS sg13g2_FILL8
XSTDFILL8_2003 VDD VSS sg13g2_FILL8
XSTDFILL8_2011 VDD VSS sg13g2_FILL8
XSTDFILL8_2019 VDD VSS sg13g2_FILL8
XSTDFILL8_2027 VDD VSS sg13g2_FILL8
XSTDFILL8_2035 VDD VSS sg13g2_FILL8
XSTDFILL8_2043 VDD VSS sg13g2_FILL8
XSTDFILL8_2051 VDD VSS sg13g2_FILL8
XSTDFILL8_2059 VDD VSS sg13g2_FILL8
XSTDFILL8_2067 VDD VSS sg13g2_FILL8
XSTDFILL8_2075 VDD VSS sg13g2_FILL8
XSTDFILL8_2083 VDD VSS sg13g2_FILL8
XSTDFILL8_2091 VDD VSS sg13g2_FILL8
XSTDFILL8_2099 VDD VSS sg13g2_FILL8
XSTDFILL8_2107 VDD VSS sg13g2_FILL8
XSTDFILL8_2115 VDD VSS sg13g2_FILL8
XSTDFILL8_2123 VDD VSS sg13g2_FILL8
XSTDFILL8_2131 VDD VSS sg13g2_FILL8
XSTDFILL8_2139 VDD VSS sg13g2_FILL8
XSTDFILL8_2147 VDD VSS sg13g2_FILL4
XSTDFILL8_2151 VDD VSS sg13g2_FILL2
XSTDFILL8_2153 VDD VSS sg13g2_FILL1
XSTDFILL9_0 VDD VSS sg13g2_FILL8
XSTDFILL9_8 VDD VSS sg13g2_FILL8
XSTDFILL9_16 VDD VSS sg13g2_FILL8
XSTDFILL9_24 VDD VSS sg13g2_FILL8
XSTDFILL9_32 VDD VSS sg13g2_FILL8
XSTDFILL9_40 VDD VSS sg13g2_FILL8
XSTDFILL9_48 VDD VSS sg13g2_FILL8
XSTDFILL9_56 VDD VSS sg13g2_FILL8
XSTDFILL9_64 VDD VSS sg13g2_FILL8
XSTDFILL9_72 VDD VSS sg13g2_FILL8
XSTDFILL9_80 VDD VSS sg13g2_FILL8
XSTDFILL9_88 VDD VSS sg13g2_FILL8
XSTDFILL9_96 VDD VSS sg13g2_FILL8
XSTDFILL9_104 VDD VSS sg13g2_FILL8
XSTDFILL9_112 VDD VSS sg13g2_FILL8
XSTDFILL9_120 VDD VSS sg13g2_FILL8
XSTDFILL9_128 VDD VSS sg13g2_FILL4
XSTDFILL9_1835 VDD VSS sg13g2_FILL8
XSTDFILL9_1843 VDD VSS sg13g2_FILL8
XSTDFILL9_1851 VDD VSS sg13g2_FILL8
XSTDFILL9_1859 VDD VSS sg13g2_FILL8
XSTDFILL9_1867 VDD VSS sg13g2_FILL8
XSTDFILL9_1875 VDD VSS sg13g2_FILL8
XSTDFILL9_1883 VDD VSS sg13g2_FILL8
XSTDFILL9_1891 VDD VSS sg13g2_FILL8
XSTDFILL9_1899 VDD VSS sg13g2_FILL8
XSTDFILL9_1907 VDD VSS sg13g2_FILL8
XSTDFILL9_1915 VDD VSS sg13g2_FILL8
XSTDFILL9_1923 VDD VSS sg13g2_FILL8
XSTDFILL9_1931 VDD VSS sg13g2_FILL8
XSTDFILL9_1939 VDD VSS sg13g2_FILL8
XSTDFILL9_1947 VDD VSS sg13g2_FILL8
XSTDFILL9_1955 VDD VSS sg13g2_FILL8
XSTDFILL9_1963 VDD VSS sg13g2_FILL8
XSTDFILL9_1971 VDD VSS sg13g2_FILL8
XSTDFILL9_1979 VDD VSS sg13g2_FILL8
XSTDFILL9_1987 VDD VSS sg13g2_FILL8
XSTDFILL9_1995 VDD VSS sg13g2_FILL8
XSTDFILL9_2003 VDD VSS sg13g2_FILL8
XSTDFILL9_2011 VDD VSS sg13g2_FILL8
XSTDFILL9_2019 VDD VSS sg13g2_FILL8
XSTDFILL9_2027 VDD VSS sg13g2_FILL8
XSTDFILL9_2035 VDD VSS sg13g2_FILL8
XSTDFILL9_2043 VDD VSS sg13g2_FILL8
XSTDFILL9_2051 VDD VSS sg13g2_FILL8
XSTDFILL9_2059 VDD VSS sg13g2_FILL8
XSTDFILL9_2067 VDD VSS sg13g2_FILL8
XSTDFILL9_2075 VDD VSS sg13g2_FILL8
XSTDFILL9_2083 VDD VSS sg13g2_FILL8
XSTDFILL9_2091 VDD VSS sg13g2_FILL8
XSTDFILL9_2099 VDD VSS sg13g2_FILL8
XSTDFILL9_2107 VDD VSS sg13g2_FILL8
XSTDFILL9_2115 VDD VSS sg13g2_FILL8
XSTDFILL9_2123 VDD VSS sg13g2_FILL8
XSTDFILL9_2131 VDD VSS sg13g2_FILL8
XSTDFILL9_2139 VDD VSS sg13g2_FILL8
XSTDFILL9_2147 VDD VSS sg13g2_FILL4
XSTDFILL9_2151 VDD VSS sg13g2_FILL2
XSTDFILL9_2153 VDD VSS sg13g2_FILL1
XSTDFILL10_0 VDD VSS sg13g2_FILL8
XSTDFILL10_8 VDD VSS sg13g2_FILL8
XSTDFILL10_16 VDD VSS sg13g2_FILL8
XSTDFILL10_24 VDD VSS sg13g2_FILL8
XSTDFILL10_32 VDD VSS sg13g2_FILL8
XSTDFILL10_40 VDD VSS sg13g2_FILL8
XSTDFILL10_48 VDD VSS sg13g2_FILL8
XSTDFILL10_56 VDD VSS sg13g2_FILL8
XSTDFILL10_64 VDD VSS sg13g2_FILL8
XSTDFILL10_72 VDD VSS sg13g2_FILL8
XSTDFILL10_80 VDD VSS sg13g2_FILL8
XSTDFILL10_88 VDD VSS sg13g2_FILL8
XSTDFILL10_96 VDD VSS sg13g2_FILL8
XSTDFILL10_104 VDD VSS sg13g2_FILL8
XSTDFILL10_112 VDD VSS sg13g2_FILL8
XSTDFILL10_120 VDD VSS sg13g2_FILL8
XSTDFILL10_128 VDD VSS sg13g2_FILL4
XSTDFILL10_1835 VDD VSS sg13g2_FILL8
XSTDFILL10_1843 VDD VSS sg13g2_FILL8
XSTDFILL10_1851 VDD VSS sg13g2_FILL8
XSTDFILL10_1859 VDD VSS sg13g2_FILL8
XSTDFILL10_1867 VDD VSS sg13g2_FILL8
XSTDFILL10_1875 VDD VSS sg13g2_FILL8
XSTDFILL10_1883 VDD VSS sg13g2_FILL8
XSTDFILL10_1891 VDD VSS sg13g2_FILL8
XSTDFILL10_1899 VDD VSS sg13g2_FILL8
XSTDFILL10_1907 VDD VSS sg13g2_FILL8
XSTDFILL10_1915 VDD VSS sg13g2_FILL8
XSTDFILL10_1923 VDD VSS sg13g2_FILL8
XSTDFILL10_1931 VDD VSS sg13g2_FILL8
XSTDFILL10_1939 VDD VSS sg13g2_FILL8
XSTDFILL10_1947 VDD VSS sg13g2_FILL8
XSTDFILL10_1955 VDD VSS sg13g2_FILL8
XSTDFILL10_1963 VDD VSS sg13g2_FILL8
XSTDFILL10_1971 VDD VSS sg13g2_FILL8
XSTDFILL10_1979 VDD VSS sg13g2_FILL8
XSTDFILL10_1987 VDD VSS sg13g2_FILL8
XSTDFILL10_1995 VDD VSS sg13g2_FILL8
XSTDFILL10_2003 VDD VSS sg13g2_FILL8
XSTDFILL10_2011 VDD VSS sg13g2_FILL8
XSTDFILL10_2019 VDD VSS sg13g2_FILL8
XSTDFILL10_2027 VDD VSS sg13g2_FILL8
XSTDFILL10_2035 VDD VSS sg13g2_FILL8
XSTDFILL10_2043 VDD VSS sg13g2_FILL8
XSTDFILL10_2051 VDD VSS sg13g2_FILL8
XSTDFILL10_2059 VDD VSS sg13g2_FILL8
XSTDFILL10_2067 VDD VSS sg13g2_FILL8
XSTDFILL10_2075 VDD VSS sg13g2_FILL8
XSTDFILL10_2083 VDD VSS sg13g2_FILL8
XSTDFILL10_2091 VDD VSS sg13g2_FILL8
XSTDFILL10_2099 VDD VSS sg13g2_FILL8
XSTDFILL10_2107 VDD VSS sg13g2_FILL8
XSTDFILL10_2115 VDD VSS sg13g2_FILL8
XSTDFILL10_2123 VDD VSS sg13g2_FILL8
XSTDFILL10_2131 VDD VSS sg13g2_FILL8
XSTDFILL10_2139 VDD VSS sg13g2_FILL8
XSTDFILL10_2147 VDD VSS sg13g2_FILL4
XSTDFILL10_2151 VDD VSS sg13g2_FILL2
XSTDFILL10_2153 VDD VSS sg13g2_FILL1
XSTDFILL11_0 VDD VSS sg13g2_FILL8
XSTDFILL11_8 VDD VSS sg13g2_FILL8
XSTDFILL11_16 VDD VSS sg13g2_FILL8
XSTDFILL11_24 VDD VSS sg13g2_FILL8
XSTDFILL11_32 VDD VSS sg13g2_FILL8
XSTDFILL11_40 VDD VSS sg13g2_FILL8
XSTDFILL11_48 VDD VSS sg13g2_FILL8
XSTDFILL11_56 VDD VSS sg13g2_FILL8
XSTDFILL11_64 VDD VSS sg13g2_FILL8
XSTDFILL11_72 VDD VSS sg13g2_FILL8
XSTDFILL11_80 VDD VSS sg13g2_FILL8
XSTDFILL11_88 VDD VSS sg13g2_FILL8
XSTDFILL11_96 VDD VSS sg13g2_FILL8
XSTDFILL11_104 VDD VSS sg13g2_FILL8
XSTDFILL11_112 VDD VSS sg13g2_FILL8
XSTDFILL11_120 VDD VSS sg13g2_FILL8
XSTDFILL11_128 VDD VSS sg13g2_FILL4
XSTDFILL11_1835 VDD VSS sg13g2_FILL8
XSTDFILL11_1843 VDD VSS sg13g2_FILL8
XSTDFILL11_1851 VDD VSS sg13g2_FILL8
XSTDFILL11_1859 VDD VSS sg13g2_FILL8
XSTDFILL11_1867 VDD VSS sg13g2_FILL8
XSTDFILL11_1875 VDD VSS sg13g2_FILL8
XSTDFILL11_1883 VDD VSS sg13g2_FILL8
XSTDFILL11_1891 VDD VSS sg13g2_FILL8
XSTDFILL11_1899 VDD VSS sg13g2_FILL8
XSTDFILL11_1907 VDD VSS sg13g2_FILL8
XSTDFILL11_1915 VDD VSS sg13g2_FILL8
XSTDFILL11_1923 VDD VSS sg13g2_FILL8
XSTDFILL11_1931 VDD VSS sg13g2_FILL8
XSTDFILL11_1939 VDD VSS sg13g2_FILL8
XSTDFILL11_1947 VDD VSS sg13g2_FILL8
XSTDFILL11_1955 VDD VSS sg13g2_FILL8
XSTDFILL11_1963 VDD VSS sg13g2_FILL8
XSTDFILL11_1971 VDD VSS sg13g2_FILL8
XSTDFILL11_1979 VDD VSS sg13g2_FILL8
XSTDFILL11_1987 VDD VSS sg13g2_FILL8
XSTDFILL11_1995 VDD VSS sg13g2_FILL8
XSTDFILL11_2003 VDD VSS sg13g2_FILL8
XSTDFILL11_2011 VDD VSS sg13g2_FILL8
XSTDFILL11_2019 VDD VSS sg13g2_FILL8
XSTDFILL11_2027 VDD VSS sg13g2_FILL8
XSTDFILL11_2035 VDD VSS sg13g2_FILL8
XSTDFILL11_2043 VDD VSS sg13g2_FILL8
XSTDFILL11_2051 VDD VSS sg13g2_FILL8
XSTDFILL11_2059 VDD VSS sg13g2_FILL8
XSTDFILL11_2067 VDD VSS sg13g2_FILL8
XSTDFILL11_2075 VDD VSS sg13g2_FILL8
XSTDFILL11_2083 VDD VSS sg13g2_FILL8
XSTDFILL11_2091 VDD VSS sg13g2_FILL8
XSTDFILL11_2099 VDD VSS sg13g2_FILL8
XSTDFILL11_2107 VDD VSS sg13g2_FILL8
XSTDFILL11_2115 VDD VSS sg13g2_FILL8
XSTDFILL11_2123 VDD VSS sg13g2_FILL8
XSTDFILL11_2131 VDD VSS sg13g2_FILL8
XSTDFILL11_2139 VDD VSS sg13g2_FILL8
XSTDFILL11_2147 VDD VSS sg13g2_FILL4
XSTDFILL11_2151 VDD VSS sg13g2_FILL2
XSTDFILL11_2153 VDD VSS sg13g2_FILL1
XSTDFILL12_0 VDD VSS sg13g2_FILL8
XSTDFILL12_8 VDD VSS sg13g2_FILL8
XSTDFILL12_16 VDD VSS sg13g2_FILL8
XSTDFILL12_24 VDD VSS sg13g2_FILL8
XSTDFILL12_32 VDD VSS sg13g2_FILL8
XSTDFILL12_40 VDD VSS sg13g2_FILL8
XSTDFILL12_48 VDD VSS sg13g2_FILL8
XSTDFILL12_56 VDD VSS sg13g2_FILL8
XSTDFILL12_64 VDD VSS sg13g2_FILL8
XSTDFILL12_72 VDD VSS sg13g2_FILL8
XSTDFILL12_80 VDD VSS sg13g2_FILL8
XSTDFILL12_88 VDD VSS sg13g2_FILL8
XSTDFILL12_96 VDD VSS sg13g2_FILL8
XSTDFILL12_104 VDD VSS sg13g2_FILL8
XSTDFILL12_112 VDD VSS sg13g2_FILL8
XSTDFILL12_120 VDD VSS sg13g2_FILL8
XSTDFILL12_128 VDD VSS sg13g2_FILL4
XSTDFILL12_1835 VDD VSS sg13g2_FILL8
XSTDFILL12_1843 VDD VSS sg13g2_FILL8
XSTDFILL12_1851 VDD VSS sg13g2_FILL8
XSTDFILL12_1859 VDD VSS sg13g2_FILL8
XSTDFILL12_1867 VDD VSS sg13g2_FILL8
XSTDFILL12_1875 VDD VSS sg13g2_FILL8
XSTDFILL12_1883 VDD VSS sg13g2_FILL8
XSTDFILL12_1891 VDD VSS sg13g2_FILL8
XSTDFILL12_1899 VDD VSS sg13g2_FILL8
XSTDFILL12_1907 VDD VSS sg13g2_FILL8
XSTDFILL12_1915 VDD VSS sg13g2_FILL8
XSTDFILL12_1923 VDD VSS sg13g2_FILL8
XSTDFILL12_1931 VDD VSS sg13g2_FILL8
XSTDFILL12_1939 VDD VSS sg13g2_FILL8
XSTDFILL12_1947 VDD VSS sg13g2_FILL8
XSTDFILL12_1955 VDD VSS sg13g2_FILL8
XSTDFILL12_1963 VDD VSS sg13g2_FILL8
XSTDFILL12_1971 VDD VSS sg13g2_FILL8
XSTDFILL12_1979 VDD VSS sg13g2_FILL8
XSTDFILL12_1987 VDD VSS sg13g2_FILL8
XSTDFILL12_1995 VDD VSS sg13g2_FILL8
XSTDFILL12_2003 VDD VSS sg13g2_FILL8
XSTDFILL12_2011 VDD VSS sg13g2_FILL8
XSTDFILL12_2019 VDD VSS sg13g2_FILL8
XSTDFILL12_2027 VDD VSS sg13g2_FILL8
XSTDFILL12_2035 VDD VSS sg13g2_FILL8
XSTDFILL12_2043 VDD VSS sg13g2_FILL8
XSTDFILL12_2051 VDD VSS sg13g2_FILL8
XSTDFILL12_2059 VDD VSS sg13g2_FILL8
XSTDFILL12_2067 VDD VSS sg13g2_FILL8
XSTDFILL12_2075 VDD VSS sg13g2_FILL8
XSTDFILL12_2083 VDD VSS sg13g2_FILL8
XSTDFILL12_2091 VDD VSS sg13g2_FILL8
XSTDFILL12_2099 VDD VSS sg13g2_FILL8
XSTDFILL12_2107 VDD VSS sg13g2_FILL8
XSTDFILL12_2115 VDD VSS sg13g2_FILL8
XSTDFILL12_2123 VDD VSS sg13g2_FILL8
XSTDFILL12_2131 VDD VSS sg13g2_FILL8
XSTDFILL12_2139 VDD VSS sg13g2_FILL8
XSTDFILL12_2147 VDD VSS sg13g2_FILL4
XSTDFILL12_2151 VDD VSS sg13g2_FILL2
XSTDFILL12_2153 VDD VSS sg13g2_FILL1
XSTDFILL13_0 VDD VSS sg13g2_FILL8
XSTDFILL13_8 VDD VSS sg13g2_FILL8
XSTDFILL13_16 VDD VSS sg13g2_FILL8
XSTDFILL13_24 VDD VSS sg13g2_FILL8
XSTDFILL13_32 VDD VSS sg13g2_FILL8
XSTDFILL13_40 VDD VSS sg13g2_FILL8
XSTDFILL13_48 VDD VSS sg13g2_FILL8
XSTDFILL13_56 VDD VSS sg13g2_FILL8
XSTDFILL13_64 VDD VSS sg13g2_FILL8
XSTDFILL13_72 VDD VSS sg13g2_FILL8
XSTDFILL13_80 VDD VSS sg13g2_FILL8
XSTDFILL13_88 VDD VSS sg13g2_FILL8
XSTDFILL13_96 VDD VSS sg13g2_FILL8
XSTDFILL13_104 VDD VSS sg13g2_FILL8
XSTDFILL13_112 VDD VSS sg13g2_FILL8
XSTDFILL13_120 VDD VSS sg13g2_FILL8
XSTDFILL13_128 VDD VSS sg13g2_FILL4
XSTDFILL13_1835 VDD VSS sg13g2_FILL8
XSTDFILL13_1843 VDD VSS sg13g2_FILL8
XSTDFILL13_1851 VDD VSS sg13g2_FILL8
XSTDFILL13_1859 VDD VSS sg13g2_FILL8
XSTDFILL13_1867 VDD VSS sg13g2_FILL8
XSTDFILL13_1875 VDD VSS sg13g2_FILL8
XSTDFILL13_1883 VDD VSS sg13g2_FILL8
XSTDFILL13_1891 VDD VSS sg13g2_FILL8
XSTDFILL13_1899 VDD VSS sg13g2_FILL8
XSTDFILL13_1907 VDD VSS sg13g2_FILL8
XSTDFILL13_1915 VDD VSS sg13g2_FILL8
XSTDFILL13_1923 VDD VSS sg13g2_FILL8
XSTDFILL13_1931 VDD VSS sg13g2_FILL8
XSTDFILL13_1939 VDD VSS sg13g2_FILL8
XSTDFILL13_1947 VDD VSS sg13g2_FILL8
XSTDFILL13_1955 VDD VSS sg13g2_FILL8
XSTDFILL13_1963 VDD VSS sg13g2_FILL8
XSTDFILL13_1971 VDD VSS sg13g2_FILL8
XSTDFILL13_1979 VDD VSS sg13g2_FILL8
XSTDFILL13_1987 VDD VSS sg13g2_FILL8
XSTDFILL13_1995 VDD VSS sg13g2_FILL8
XSTDFILL13_2003 VDD VSS sg13g2_FILL8
XSTDFILL13_2011 VDD VSS sg13g2_FILL8
XSTDFILL13_2019 VDD VSS sg13g2_FILL8
XSTDFILL13_2027 VDD VSS sg13g2_FILL8
XSTDFILL13_2035 VDD VSS sg13g2_FILL8
XSTDFILL13_2043 VDD VSS sg13g2_FILL8
XSTDFILL13_2051 VDD VSS sg13g2_FILL8
XSTDFILL13_2059 VDD VSS sg13g2_FILL8
XSTDFILL13_2067 VDD VSS sg13g2_FILL8
XSTDFILL13_2075 VDD VSS sg13g2_FILL8
XSTDFILL13_2083 VDD VSS sg13g2_FILL8
XSTDFILL13_2091 VDD VSS sg13g2_FILL8
XSTDFILL13_2099 VDD VSS sg13g2_FILL8
XSTDFILL13_2107 VDD VSS sg13g2_FILL8
XSTDFILL13_2115 VDD VSS sg13g2_FILL8
XSTDFILL13_2123 VDD VSS sg13g2_FILL8
XSTDFILL13_2131 VDD VSS sg13g2_FILL8
XSTDFILL13_2139 VDD VSS sg13g2_FILL8
XSTDFILL13_2147 VDD VSS sg13g2_FILL4
XSTDFILL13_2151 VDD VSS sg13g2_FILL2
XSTDFILL13_2153 VDD VSS sg13g2_FILL1
XSTDFILL14_0 VDD VSS sg13g2_FILL8
XSTDFILL14_8 VDD VSS sg13g2_FILL8
XSTDFILL14_16 VDD VSS sg13g2_FILL8
XSTDFILL14_24 VDD VSS sg13g2_FILL8
XSTDFILL14_32 VDD VSS sg13g2_FILL8
XSTDFILL14_40 VDD VSS sg13g2_FILL8
XSTDFILL14_48 VDD VSS sg13g2_FILL8
XSTDFILL14_56 VDD VSS sg13g2_FILL8
XSTDFILL14_64 VDD VSS sg13g2_FILL8
XSTDFILL14_72 VDD VSS sg13g2_FILL8
XSTDFILL14_80 VDD VSS sg13g2_FILL8
XSTDFILL14_88 VDD VSS sg13g2_FILL8
XSTDFILL14_96 VDD VSS sg13g2_FILL8
XSTDFILL14_104 VDD VSS sg13g2_FILL8
XSTDFILL14_112 VDD VSS sg13g2_FILL8
XSTDFILL14_120 VDD VSS sg13g2_FILL8
XSTDFILL14_128 VDD VSS sg13g2_FILL4
XSTDFILL14_1835 VDD VSS sg13g2_FILL8
XSTDFILL14_1843 VDD VSS sg13g2_FILL8
XSTDFILL14_1851 VDD VSS sg13g2_FILL8
XSTDFILL14_1859 VDD VSS sg13g2_FILL8
XSTDFILL14_1867 VDD VSS sg13g2_FILL8
XSTDFILL14_1875 VDD VSS sg13g2_FILL8
XSTDFILL14_1883 VDD VSS sg13g2_FILL8
XSTDFILL14_1891 VDD VSS sg13g2_FILL8
XSTDFILL14_1899 VDD VSS sg13g2_FILL8
XSTDFILL14_1907 VDD VSS sg13g2_FILL8
XSTDFILL14_1915 VDD VSS sg13g2_FILL8
XSTDFILL14_1923 VDD VSS sg13g2_FILL8
XSTDFILL14_1931 VDD VSS sg13g2_FILL8
XSTDFILL14_1939 VDD VSS sg13g2_FILL8
XSTDFILL14_1947 VDD VSS sg13g2_FILL8
XSTDFILL14_1955 VDD VSS sg13g2_FILL8
XSTDFILL14_1963 VDD VSS sg13g2_FILL8
XSTDFILL14_1971 VDD VSS sg13g2_FILL8
XSTDFILL14_1979 VDD VSS sg13g2_FILL8
XSTDFILL14_1987 VDD VSS sg13g2_FILL8
XSTDFILL14_1995 VDD VSS sg13g2_FILL8
XSTDFILL14_2003 VDD VSS sg13g2_FILL8
XSTDFILL14_2011 VDD VSS sg13g2_FILL8
XSTDFILL14_2019 VDD VSS sg13g2_FILL8
XSTDFILL14_2027 VDD VSS sg13g2_FILL8
XSTDFILL14_2035 VDD VSS sg13g2_FILL8
XSTDFILL14_2043 VDD VSS sg13g2_FILL8
XSTDFILL14_2051 VDD VSS sg13g2_FILL8
XSTDFILL14_2059 VDD VSS sg13g2_FILL8
XSTDFILL14_2067 VDD VSS sg13g2_FILL8
XSTDFILL14_2075 VDD VSS sg13g2_FILL8
XSTDFILL14_2083 VDD VSS sg13g2_FILL8
XSTDFILL14_2091 VDD VSS sg13g2_FILL8
XSTDFILL14_2099 VDD VSS sg13g2_FILL8
XSTDFILL14_2107 VDD VSS sg13g2_FILL8
XSTDFILL14_2115 VDD VSS sg13g2_FILL8
XSTDFILL14_2123 VDD VSS sg13g2_FILL8
XSTDFILL14_2131 VDD VSS sg13g2_FILL8
XSTDFILL14_2139 VDD VSS sg13g2_FILL8
XSTDFILL14_2147 VDD VSS sg13g2_FILL4
XSTDFILL14_2151 VDD VSS sg13g2_FILL2
XSTDFILL14_2153 VDD VSS sg13g2_FILL1
XSTDFILL15_0 VDD VSS sg13g2_FILL8
XSTDFILL15_8 VDD VSS sg13g2_FILL8
XSTDFILL15_16 VDD VSS sg13g2_FILL8
XSTDFILL15_24 VDD VSS sg13g2_FILL8
XSTDFILL15_32 VDD VSS sg13g2_FILL8
XSTDFILL15_40 VDD VSS sg13g2_FILL8
XSTDFILL15_48 VDD VSS sg13g2_FILL8
XSTDFILL15_56 VDD VSS sg13g2_FILL8
XSTDFILL15_64 VDD VSS sg13g2_FILL8
XSTDFILL15_72 VDD VSS sg13g2_FILL8
XSTDFILL15_80 VDD VSS sg13g2_FILL8
XSTDFILL15_88 VDD VSS sg13g2_FILL8
XSTDFILL15_96 VDD VSS sg13g2_FILL8
XSTDFILL15_104 VDD VSS sg13g2_FILL8
XSTDFILL15_112 VDD VSS sg13g2_FILL8
XSTDFILL15_120 VDD VSS sg13g2_FILL8
XSTDFILL15_128 VDD VSS sg13g2_FILL4
XSTDFILL15_1835 VDD VSS sg13g2_FILL8
XSTDFILL15_1843 VDD VSS sg13g2_FILL8
XSTDFILL15_1851 VDD VSS sg13g2_FILL8
XSTDFILL15_1859 VDD VSS sg13g2_FILL8
XSTDFILL15_1867 VDD VSS sg13g2_FILL8
XSTDFILL15_1875 VDD VSS sg13g2_FILL8
XSTDFILL15_1883 VDD VSS sg13g2_FILL8
XSTDFILL15_1891 VDD VSS sg13g2_FILL8
XSTDFILL15_1899 VDD VSS sg13g2_FILL8
XSTDFILL15_1907 VDD VSS sg13g2_FILL8
XSTDFILL15_1915 VDD VSS sg13g2_FILL8
XSTDFILL15_1923 VDD VSS sg13g2_FILL8
XSTDFILL15_1931 VDD VSS sg13g2_FILL8
XSTDFILL15_1939 VDD VSS sg13g2_FILL8
XSTDFILL15_1947 VDD VSS sg13g2_FILL8
XSTDFILL15_1955 VDD VSS sg13g2_FILL8
XSTDFILL15_1963 VDD VSS sg13g2_FILL8
XSTDFILL15_1971 VDD VSS sg13g2_FILL8
XSTDFILL15_1979 VDD VSS sg13g2_FILL8
XSTDFILL15_1987 VDD VSS sg13g2_FILL8
XSTDFILL15_1995 VDD VSS sg13g2_FILL8
XSTDFILL15_2003 VDD VSS sg13g2_FILL8
XSTDFILL15_2011 VDD VSS sg13g2_FILL8
XSTDFILL15_2019 VDD VSS sg13g2_FILL8
XSTDFILL15_2027 VDD VSS sg13g2_FILL8
XSTDFILL15_2035 VDD VSS sg13g2_FILL8
XSTDFILL15_2043 VDD VSS sg13g2_FILL8
XSTDFILL15_2051 VDD VSS sg13g2_FILL8
XSTDFILL15_2059 VDD VSS sg13g2_FILL8
XSTDFILL15_2067 VDD VSS sg13g2_FILL8
XSTDFILL15_2075 VDD VSS sg13g2_FILL8
XSTDFILL15_2083 VDD VSS sg13g2_FILL8
XSTDFILL15_2091 VDD VSS sg13g2_FILL8
XSTDFILL15_2099 VDD VSS sg13g2_FILL8
XSTDFILL15_2107 VDD VSS sg13g2_FILL8
XSTDFILL15_2115 VDD VSS sg13g2_FILL8
XSTDFILL15_2123 VDD VSS sg13g2_FILL8
XSTDFILL15_2131 VDD VSS sg13g2_FILL8
XSTDFILL15_2139 VDD VSS sg13g2_FILL8
XSTDFILL15_2147 VDD VSS sg13g2_FILL4
XSTDFILL15_2151 VDD VSS sg13g2_FILL2
XSTDFILL15_2153 VDD VSS sg13g2_FILL1
XSTDFILL16_0 VDD VSS sg13g2_FILL8
XSTDFILL16_8 VDD VSS sg13g2_FILL8
XSTDFILL16_16 VDD VSS sg13g2_FILL8
XSTDFILL16_24 VDD VSS sg13g2_FILL8
XSTDFILL16_32 VDD VSS sg13g2_FILL8
XSTDFILL16_40 VDD VSS sg13g2_FILL8
XSTDFILL16_48 VDD VSS sg13g2_FILL8
XSTDFILL16_56 VDD VSS sg13g2_FILL8
XSTDFILL16_64 VDD VSS sg13g2_FILL8
XSTDFILL16_72 VDD VSS sg13g2_FILL8
XSTDFILL16_80 VDD VSS sg13g2_FILL8
XSTDFILL16_88 VDD VSS sg13g2_FILL8
XSTDFILL16_96 VDD VSS sg13g2_FILL8
XSTDFILL16_104 VDD VSS sg13g2_FILL8
XSTDFILL16_112 VDD VSS sg13g2_FILL8
XSTDFILL16_120 VDD VSS sg13g2_FILL8
XSTDFILL16_128 VDD VSS sg13g2_FILL4
XSTDFILL16_1835 VDD VSS sg13g2_FILL8
XSTDFILL16_1843 VDD VSS sg13g2_FILL8
XSTDFILL16_1851 VDD VSS sg13g2_FILL8
XSTDFILL16_1859 VDD VSS sg13g2_FILL8
XSTDFILL16_1867 VDD VSS sg13g2_FILL8
XSTDFILL16_1875 VDD VSS sg13g2_FILL8
XSTDFILL16_1883 VDD VSS sg13g2_FILL8
XSTDFILL16_1891 VDD VSS sg13g2_FILL8
XSTDFILL16_1899 VDD VSS sg13g2_FILL8
XSTDFILL16_1907 VDD VSS sg13g2_FILL8
XSTDFILL16_1915 VDD VSS sg13g2_FILL8
XSTDFILL16_1923 VDD VSS sg13g2_FILL8
XSTDFILL16_1931 VDD VSS sg13g2_FILL8
XSTDFILL16_1939 VDD VSS sg13g2_FILL8
XSTDFILL16_1947 VDD VSS sg13g2_FILL8
XSTDFILL16_1955 VDD VSS sg13g2_FILL8
XSTDFILL16_1963 VDD VSS sg13g2_FILL8
XSTDFILL16_1971 VDD VSS sg13g2_FILL8
XSTDFILL16_1979 VDD VSS sg13g2_FILL8
XSTDFILL16_1987 VDD VSS sg13g2_FILL8
XSTDFILL16_1995 VDD VSS sg13g2_FILL8
XSTDFILL16_2003 VDD VSS sg13g2_FILL8
XSTDFILL16_2011 VDD VSS sg13g2_FILL8
XSTDFILL16_2019 VDD VSS sg13g2_FILL8
XSTDFILL16_2027 VDD VSS sg13g2_FILL8
XSTDFILL16_2035 VDD VSS sg13g2_FILL8
XSTDFILL16_2043 VDD VSS sg13g2_FILL8
XSTDFILL16_2051 VDD VSS sg13g2_FILL8
XSTDFILL16_2059 VDD VSS sg13g2_FILL8
XSTDFILL16_2067 VDD VSS sg13g2_FILL8
XSTDFILL16_2075 VDD VSS sg13g2_FILL8
XSTDFILL16_2083 VDD VSS sg13g2_FILL8
XSTDFILL16_2091 VDD VSS sg13g2_FILL8
XSTDFILL16_2099 VDD VSS sg13g2_FILL8
XSTDFILL16_2107 VDD VSS sg13g2_FILL8
XSTDFILL16_2115 VDD VSS sg13g2_FILL8
XSTDFILL16_2123 VDD VSS sg13g2_FILL8
XSTDFILL16_2131 VDD VSS sg13g2_FILL8
XSTDFILL16_2139 VDD VSS sg13g2_FILL8
XSTDFILL16_2147 VDD VSS sg13g2_FILL4
XSTDFILL16_2151 VDD VSS sg13g2_FILL2
XSTDFILL16_2153 VDD VSS sg13g2_FILL1
XSTDFILL17_0 VDD VSS sg13g2_FILL8
XSTDFILL17_8 VDD VSS sg13g2_FILL8
XSTDFILL17_16 VDD VSS sg13g2_FILL8
XSTDFILL17_24 VDD VSS sg13g2_FILL8
XSTDFILL17_32 VDD VSS sg13g2_FILL8
XSTDFILL17_40 VDD VSS sg13g2_FILL8
XSTDFILL17_48 VDD VSS sg13g2_FILL8
XSTDFILL17_56 VDD VSS sg13g2_FILL8
XSTDFILL17_64 VDD VSS sg13g2_FILL8
XSTDFILL17_72 VDD VSS sg13g2_FILL8
XSTDFILL17_80 VDD VSS sg13g2_FILL8
XSTDFILL17_88 VDD VSS sg13g2_FILL8
XSTDFILL17_96 VDD VSS sg13g2_FILL8
XSTDFILL17_104 VDD VSS sg13g2_FILL8
XSTDFILL17_112 VDD VSS sg13g2_FILL8
XSTDFILL17_120 VDD VSS sg13g2_FILL8
XSTDFILL17_128 VDD VSS sg13g2_FILL4
XSTDFILL17_1835 VDD VSS sg13g2_FILL8
XSTDFILL17_1843 VDD VSS sg13g2_FILL8
XSTDFILL17_1851 VDD VSS sg13g2_FILL8
XSTDFILL17_1859 VDD VSS sg13g2_FILL8
XSTDFILL17_1867 VDD VSS sg13g2_FILL8
XSTDFILL17_1875 VDD VSS sg13g2_FILL8
XSTDFILL17_1883 VDD VSS sg13g2_FILL8
XSTDFILL17_1891 VDD VSS sg13g2_FILL8
XSTDFILL17_1899 VDD VSS sg13g2_FILL8
XSTDFILL17_1907 VDD VSS sg13g2_FILL8
XSTDFILL17_1915 VDD VSS sg13g2_FILL8
XSTDFILL17_1923 VDD VSS sg13g2_FILL8
XSTDFILL17_1931 VDD VSS sg13g2_FILL8
XSTDFILL17_1939 VDD VSS sg13g2_FILL8
XSTDFILL17_1947 VDD VSS sg13g2_FILL8
XSTDFILL17_1955 VDD VSS sg13g2_FILL8
XSTDFILL17_1963 VDD VSS sg13g2_FILL8
XSTDFILL17_1971 VDD VSS sg13g2_FILL8
XSTDFILL17_1979 VDD VSS sg13g2_FILL8
XSTDFILL17_1987 VDD VSS sg13g2_FILL8
XSTDFILL17_1995 VDD VSS sg13g2_FILL8
XSTDFILL17_2003 VDD VSS sg13g2_FILL8
XSTDFILL17_2011 VDD VSS sg13g2_FILL8
XSTDFILL17_2019 VDD VSS sg13g2_FILL8
XSTDFILL17_2027 VDD VSS sg13g2_FILL8
XSTDFILL17_2035 VDD VSS sg13g2_FILL8
XSTDFILL17_2043 VDD VSS sg13g2_FILL8
XSTDFILL17_2051 VDD VSS sg13g2_FILL8
XSTDFILL17_2059 VDD VSS sg13g2_FILL8
XSTDFILL17_2067 VDD VSS sg13g2_FILL8
XSTDFILL17_2075 VDD VSS sg13g2_FILL8
XSTDFILL17_2083 VDD VSS sg13g2_FILL8
XSTDFILL17_2091 VDD VSS sg13g2_FILL8
XSTDFILL17_2099 VDD VSS sg13g2_FILL8
XSTDFILL17_2107 VDD VSS sg13g2_FILL8
XSTDFILL17_2115 VDD VSS sg13g2_FILL8
XSTDFILL17_2123 VDD VSS sg13g2_FILL8
XSTDFILL17_2131 VDD VSS sg13g2_FILL8
XSTDFILL17_2139 VDD VSS sg13g2_FILL8
XSTDFILL17_2147 VDD VSS sg13g2_FILL4
XSTDFILL17_2151 VDD VSS sg13g2_FILL2
XSTDFILL17_2153 VDD VSS sg13g2_FILL1
XSTDFILL18_0 VDD VSS sg13g2_FILL8
XSTDFILL18_8 VDD VSS sg13g2_FILL8
XSTDFILL18_16 VDD VSS sg13g2_FILL8
XSTDFILL18_24 VDD VSS sg13g2_FILL8
XSTDFILL18_32 VDD VSS sg13g2_FILL8
XSTDFILL18_40 VDD VSS sg13g2_FILL8
XSTDFILL18_48 VDD VSS sg13g2_FILL8
XSTDFILL18_56 VDD VSS sg13g2_FILL8
XSTDFILL18_64 VDD VSS sg13g2_FILL8
XSTDFILL18_72 VDD VSS sg13g2_FILL8
XSTDFILL18_80 VDD VSS sg13g2_FILL8
XSTDFILL18_88 VDD VSS sg13g2_FILL8
XSTDFILL18_96 VDD VSS sg13g2_FILL8
XSTDFILL18_104 VDD VSS sg13g2_FILL8
XSTDFILL18_112 VDD VSS sg13g2_FILL8
XSTDFILL18_120 VDD VSS sg13g2_FILL8
XSTDFILL18_128 VDD VSS sg13g2_FILL4
XSTDFILL18_1835 VDD VSS sg13g2_FILL8
XSTDFILL18_1843 VDD VSS sg13g2_FILL8
XSTDFILL18_1851 VDD VSS sg13g2_FILL8
XSTDFILL18_1859 VDD VSS sg13g2_FILL8
XSTDFILL18_1867 VDD VSS sg13g2_FILL8
XSTDFILL18_1875 VDD VSS sg13g2_FILL8
XSTDFILL18_1883 VDD VSS sg13g2_FILL8
XSTDFILL18_1891 VDD VSS sg13g2_FILL8
XSTDFILL18_1899 VDD VSS sg13g2_FILL8
XSTDFILL18_1907 VDD VSS sg13g2_FILL8
XSTDFILL18_1915 VDD VSS sg13g2_FILL8
XSTDFILL18_1923 VDD VSS sg13g2_FILL8
XSTDFILL18_1931 VDD VSS sg13g2_FILL8
XSTDFILL18_1939 VDD VSS sg13g2_FILL8
XSTDFILL18_1947 VDD VSS sg13g2_FILL8
XSTDFILL18_1955 VDD VSS sg13g2_FILL8
XSTDFILL18_1963 VDD VSS sg13g2_FILL8
XSTDFILL18_1971 VDD VSS sg13g2_FILL8
XSTDFILL18_1979 VDD VSS sg13g2_FILL8
XSTDFILL18_1987 VDD VSS sg13g2_FILL8
XSTDFILL18_1995 VDD VSS sg13g2_FILL8
XSTDFILL18_2003 VDD VSS sg13g2_FILL8
XSTDFILL18_2011 VDD VSS sg13g2_FILL8
XSTDFILL18_2019 VDD VSS sg13g2_FILL8
XSTDFILL18_2027 VDD VSS sg13g2_FILL8
XSTDFILL18_2035 VDD VSS sg13g2_FILL8
XSTDFILL18_2043 VDD VSS sg13g2_FILL8
XSTDFILL18_2051 VDD VSS sg13g2_FILL8
XSTDFILL18_2059 VDD VSS sg13g2_FILL8
XSTDFILL18_2067 VDD VSS sg13g2_FILL8
XSTDFILL18_2075 VDD VSS sg13g2_FILL8
XSTDFILL18_2083 VDD VSS sg13g2_FILL8
XSTDFILL18_2091 VDD VSS sg13g2_FILL8
XSTDFILL18_2099 VDD VSS sg13g2_FILL8
XSTDFILL18_2107 VDD VSS sg13g2_FILL8
XSTDFILL18_2115 VDD VSS sg13g2_FILL8
XSTDFILL18_2123 VDD VSS sg13g2_FILL8
XSTDFILL18_2131 VDD VSS sg13g2_FILL8
XSTDFILL18_2139 VDD VSS sg13g2_FILL8
XSTDFILL18_2147 VDD VSS sg13g2_FILL4
XSTDFILL18_2151 VDD VSS sg13g2_FILL2
XSTDFILL18_2153 VDD VSS sg13g2_FILL1
XSTDFILL19_0 VDD VSS sg13g2_FILL8
XSTDFILL19_8 VDD VSS sg13g2_FILL8
XSTDFILL19_16 VDD VSS sg13g2_FILL8
XSTDFILL19_24 VDD VSS sg13g2_FILL8
XSTDFILL19_32 VDD VSS sg13g2_FILL8
XSTDFILL19_40 VDD VSS sg13g2_FILL8
XSTDFILL19_48 VDD VSS sg13g2_FILL8
XSTDFILL19_56 VDD VSS sg13g2_FILL8
XSTDFILL19_64 VDD VSS sg13g2_FILL8
XSTDFILL19_72 VDD VSS sg13g2_FILL8
XSTDFILL19_80 VDD VSS sg13g2_FILL8
XSTDFILL19_88 VDD VSS sg13g2_FILL8
XSTDFILL19_96 VDD VSS sg13g2_FILL8
XSTDFILL19_104 VDD VSS sg13g2_FILL8
XSTDFILL19_112 VDD VSS sg13g2_FILL8
XSTDFILL19_120 VDD VSS sg13g2_FILL8
XSTDFILL19_128 VDD VSS sg13g2_FILL4
XSTDFILL19_1835 VDD VSS sg13g2_FILL8
XSTDFILL19_1843 VDD VSS sg13g2_FILL8
XSTDFILL19_1851 VDD VSS sg13g2_FILL8
XSTDFILL19_1859 VDD VSS sg13g2_FILL8
XSTDFILL19_1867 VDD VSS sg13g2_FILL8
XSTDFILL19_1875 VDD VSS sg13g2_FILL8
XSTDFILL19_1883 VDD VSS sg13g2_FILL8
XSTDFILL19_1891 VDD VSS sg13g2_FILL8
XSTDFILL19_1899 VDD VSS sg13g2_FILL8
XSTDFILL19_1907 VDD VSS sg13g2_FILL8
XSTDFILL19_1915 VDD VSS sg13g2_FILL8
XSTDFILL19_1923 VDD VSS sg13g2_FILL8
XSTDFILL19_1931 VDD VSS sg13g2_FILL8
XSTDFILL19_1939 VDD VSS sg13g2_FILL8
XSTDFILL19_1947 VDD VSS sg13g2_FILL8
XSTDFILL19_1955 VDD VSS sg13g2_FILL8
XSTDFILL19_1963 VDD VSS sg13g2_FILL8
XSTDFILL19_1971 VDD VSS sg13g2_FILL8
XSTDFILL19_1979 VDD VSS sg13g2_FILL8
XSTDFILL19_1987 VDD VSS sg13g2_FILL8
XSTDFILL19_1995 VDD VSS sg13g2_FILL8
XSTDFILL19_2003 VDD VSS sg13g2_FILL8
XSTDFILL19_2011 VDD VSS sg13g2_FILL8
XSTDFILL19_2019 VDD VSS sg13g2_FILL8
XSTDFILL19_2027 VDD VSS sg13g2_FILL8
XSTDFILL19_2035 VDD VSS sg13g2_FILL8
XSTDFILL19_2043 VDD VSS sg13g2_FILL8
XSTDFILL19_2051 VDD VSS sg13g2_FILL8
XSTDFILL19_2059 VDD VSS sg13g2_FILL8
XSTDFILL19_2067 VDD VSS sg13g2_FILL8
XSTDFILL19_2075 VDD VSS sg13g2_FILL8
XSTDFILL19_2083 VDD VSS sg13g2_FILL8
XSTDFILL19_2091 VDD VSS sg13g2_FILL8
XSTDFILL19_2099 VDD VSS sg13g2_FILL8
XSTDFILL19_2107 VDD VSS sg13g2_FILL8
XSTDFILL19_2115 VDD VSS sg13g2_FILL8
XSTDFILL19_2123 VDD VSS sg13g2_FILL8
XSTDFILL19_2131 VDD VSS sg13g2_FILL8
XSTDFILL19_2139 VDD VSS sg13g2_FILL8
XSTDFILL19_2147 VDD VSS sg13g2_FILL4
XSTDFILL19_2151 VDD VSS sg13g2_FILL2
XSTDFILL19_2153 VDD VSS sg13g2_FILL1
XSTDFILL20_0 VDD VSS sg13g2_FILL8
XSTDFILL20_8 VDD VSS sg13g2_FILL8
XSTDFILL20_16 VDD VSS sg13g2_FILL8
XSTDFILL20_24 VDD VSS sg13g2_FILL8
XSTDFILL20_32 VDD VSS sg13g2_FILL8
XSTDFILL20_40 VDD VSS sg13g2_FILL8
XSTDFILL20_48 VDD VSS sg13g2_FILL8
XSTDFILL20_56 VDD VSS sg13g2_FILL8
XSTDFILL20_64 VDD VSS sg13g2_FILL8
XSTDFILL20_72 VDD VSS sg13g2_FILL8
XSTDFILL20_80 VDD VSS sg13g2_FILL8
XSTDFILL20_88 VDD VSS sg13g2_FILL8
XSTDFILL20_96 VDD VSS sg13g2_FILL8
XSTDFILL20_104 VDD VSS sg13g2_FILL8
XSTDFILL20_112 VDD VSS sg13g2_FILL8
XSTDFILL20_120 VDD VSS sg13g2_FILL8
XSTDFILL20_128 VDD VSS sg13g2_FILL4
XSTDFILL20_1835 VDD VSS sg13g2_FILL8
XSTDFILL20_1843 VDD VSS sg13g2_FILL8
XSTDFILL20_1851 VDD VSS sg13g2_FILL8
XSTDFILL20_1859 VDD VSS sg13g2_FILL8
XSTDFILL20_1867 VDD VSS sg13g2_FILL8
XSTDFILL20_1875 VDD VSS sg13g2_FILL8
XSTDFILL20_1883 VDD VSS sg13g2_FILL8
XSTDFILL20_1891 VDD VSS sg13g2_FILL8
XSTDFILL20_1899 VDD VSS sg13g2_FILL8
XSTDFILL20_1907 VDD VSS sg13g2_FILL8
XSTDFILL20_1915 VDD VSS sg13g2_FILL8
XSTDFILL20_1923 VDD VSS sg13g2_FILL8
XSTDFILL20_1931 VDD VSS sg13g2_FILL8
XSTDFILL20_1939 VDD VSS sg13g2_FILL8
XSTDFILL20_1947 VDD VSS sg13g2_FILL8
XSTDFILL20_1955 VDD VSS sg13g2_FILL8
XSTDFILL20_1963 VDD VSS sg13g2_FILL8
XSTDFILL20_1971 VDD VSS sg13g2_FILL8
XSTDFILL20_1979 VDD VSS sg13g2_FILL8
XSTDFILL20_1987 VDD VSS sg13g2_FILL8
XSTDFILL20_1995 VDD VSS sg13g2_FILL8
XSTDFILL20_2003 VDD VSS sg13g2_FILL8
XSTDFILL20_2011 VDD VSS sg13g2_FILL8
XSTDFILL20_2019 VDD VSS sg13g2_FILL8
XSTDFILL20_2027 VDD VSS sg13g2_FILL8
XSTDFILL20_2035 VDD VSS sg13g2_FILL8
XSTDFILL20_2043 VDD VSS sg13g2_FILL8
XSTDFILL20_2051 VDD VSS sg13g2_FILL8
XSTDFILL20_2059 VDD VSS sg13g2_FILL8
XSTDFILL20_2067 VDD VSS sg13g2_FILL8
XSTDFILL20_2075 VDD VSS sg13g2_FILL8
XSTDFILL20_2083 VDD VSS sg13g2_FILL8
XSTDFILL20_2091 VDD VSS sg13g2_FILL8
XSTDFILL20_2099 VDD VSS sg13g2_FILL8
XSTDFILL20_2107 VDD VSS sg13g2_FILL8
XSTDFILL20_2115 VDD VSS sg13g2_FILL8
XSTDFILL20_2123 VDD VSS sg13g2_FILL8
XSTDFILL20_2131 VDD VSS sg13g2_FILL8
XSTDFILL20_2139 VDD VSS sg13g2_FILL8
XSTDFILL20_2147 VDD VSS sg13g2_FILL4
XSTDFILL20_2151 VDD VSS sg13g2_FILL2
XSTDFILL20_2153 VDD VSS sg13g2_FILL1
XSTDFILL21_0 VDD VSS sg13g2_FILL8
XSTDFILL21_8 VDD VSS sg13g2_FILL8
XSTDFILL21_16 VDD VSS sg13g2_FILL8
XSTDFILL21_24 VDD VSS sg13g2_FILL8
XSTDFILL21_32 VDD VSS sg13g2_FILL8
XSTDFILL21_40 VDD VSS sg13g2_FILL8
XSTDFILL21_48 VDD VSS sg13g2_FILL8
XSTDFILL21_56 VDD VSS sg13g2_FILL8
XSTDFILL21_64 VDD VSS sg13g2_FILL8
XSTDFILL21_72 VDD VSS sg13g2_FILL8
XSTDFILL21_80 VDD VSS sg13g2_FILL8
XSTDFILL21_88 VDD VSS sg13g2_FILL8
XSTDFILL21_96 VDD VSS sg13g2_FILL8
XSTDFILL21_104 VDD VSS sg13g2_FILL8
XSTDFILL21_112 VDD VSS sg13g2_FILL8
XSTDFILL21_120 VDD VSS sg13g2_FILL8
XSTDFILL21_128 VDD VSS sg13g2_FILL4
XSTDFILL21_1835 VDD VSS sg13g2_FILL8
XSTDFILL21_1843 VDD VSS sg13g2_FILL8
XSTDFILL21_1851 VDD VSS sg13g2_FILL8
XSTDFILL21_1859 VDD VSS sg13g2_FILL8
XSTDFILL21_1867 VDD VSS sg13g2_FILL8
XSTDFILL21_1875 VDD VSS sg13g2_FILL8
XSTDFILL21_1883 VDD VSS sg13g2_FILL8
XSTDFILL21_1891 VDD VSS sg13g2_FILL8
XSTDFILL21_1899 VDD VSS sg13g2_FILL8
XSTDFILL21_1907 VDD VSS sg13g2_FILL8
XSTDFILL21_1915 VDD VSS sg13g2_FILL8
XSTDFILL21_1923 VDD VSS sg13g2_FILL8
XSTDFILL21_1931 VDD VSS sg13g2_FILL8
XSTDFILL21_1939 VDD VSS sg13g2_FILL8
XSTDFILL21_1947 VDD VSS sg13g2_FILL8
XSTDFILL21_1955 VDD VSS sg13g2_FILL8
XSTDFILL21_1963 VDD VSS sg13g2_FILL8
XSTDFILL21_1971 VDD VSS sg13g2_FILL8
XSTDFILL21_1979 VDD VSS sg13g2_FILL8
XSTDFILL21_1987 VDD VSS sg13g2_FILL8
XSTDFILL21_1995 VDD VSS sg13g2_FILL8
XSTDFILL21_2003 VDD VSS sg13g2_FILL8
XSTDFILL21_2011 VDD VSS sg13g2_FILL8
XSTDFILL21_2019 VDD VSS sg13g2_FILL8
XSTDFILL21_2027 VDD VSS sg13g2_FILL8
XSTDFILL21_2035 VDD VSS sg13g2_FILL8
XSTDFILL21_2043 VDD VSS sg13g2_FILL8
XSTDFILL21_2051 VDD VSS sg13g2_FILL8
XSTDFILL21_2059 VDD VSS sg13g2_FILL8
XSTDFILL21_2067 VDD VSS sg13g2_FILL8
XSTDFILL21_2075 VDD VSS sg13g2_FILL8
XSTDFILL21_2083 VDD VSS sg13g2_FILL8
XSTDFILL21_2091 VDD VSS sg13g2_FILL8
XSTDFILL21_2099 VDD VSS sg13g2_FILL8
XSTDFILL21_2107 VDD VSS sg13g2_FILL8
XSTDFILL21_2115 VDD VSS sg13g2_FILL8
XSTDFILL21_2123 VDD VSS sg13g2_FILL8
XSTDFILL21_2131 VDD VSS sg13g2_FILL8
XSTDFILL21_2139 VDD VSS sg13g2_FILL8
XSTDFILL21_2147 VDD VSS sg13g2_FILL4
XSTDFILL21_2151 VDD VSS sg13g2_FILL2
XSTDFILL21_2153 VDD VSS sg13g2_FILL1
XSTDFILL22_0 VDD VSS sg13g2_FILL8
XSTDFILL22_8 VDD VSS sg13g2_FILL8
XSTDFILL22_16 VDD VSS sg13g2_FILL8
XSTDFILL22_24 VDD VSS sg13g2_FILL8
XSTDFILL22_32 VDD VSS sg13g2_FILL8
XSTDFILL22_40 VDD VSS sg13g2_FILL8
XSTDFILL22_48 VDD VSS sg13g2_FILL8
XSTDFILL22_56 VDD VSS sg13g2_FILL8
XSTDFILL22_64 VDD VSS sg13g2_FILL8
XSTDFILL22_72 VDD VSS sg13g2_FILL8
XSTDFILL22_80 VDD VSS sg13g2_FILL8
XSTDFILL22_88 VDD VSS sg13g2_FILL8
XSTDFILL22_96 VDD VSS sg13g2_FILL8
XSTDFILL22_104 VDD VSS sg13g2_FILL8
XSTDFILL22_112 VDD VSS sg13g2_FILL8
XSTDFILL22_120 VDD VSS sg13g2_FILL8
XSTDFILL22_128 VDD VSS sg13g2_FILL4
XSTDFILL22_1835 VDD VSS sg13g2_FILL8
XSTDFILL22_1843 VDD VSS sg13g2_FILL8
XSTDFILL22_1851 VDD VSS sg13g2_FILL8
XSTDFILL22_1859 VDD VSS sg13g2_FILL8
XSTDFILL22_1867 VDD VSS sg13g2_FILL8
XSTDFILL22_1875 VDD VSS sg13g2_FILL8
XSTDFILL22_1883 VDD VSS sg13g2_FILL8
XSTDFILL22_1891 VDD VSS sg13g2_FILL8
XSTDFILL22_1899 VDD VSS sg13g2_FILL8
XSTDFILL22_1907 VDD VSS sg13g2_FILL8
XSTDFILL22_1915 VDD VSS sg13g2_FILL8
XSTDFILL22_1923 VDD VSS sg13g2_FILL8
XSTDFILL22_1931 VDD VSS sg13g2_FILL8
XSTDFILL22_1939 VDD VSS sg13g2_FILL8
XSTDFILL22_1947 VDD VSS sg13g2_FILL8
XSTDFILL22_1955 VDD VSS sg13g2_FILL8
XSTDFILL22_1963 VDD VSS sg13g2_FILL8
XSTDFILL22_1971 VDD VSS sg13g2_FILL8
XSTDFILL22_1979 VDD VSS sg13g2_FILL8
XSTDFILL22_1987 VDD VSS sg13g2_FILL8
XSTDFILL22_1995 VDD VSS sg13g2_FILL8
XSTDFILL22_2003 VDD VSS sg13g2_FILL8
XSTDFILL22_2011 VDD VSS sg13g2_FILL8
XSTDFILL22_2019 VDD VSS sg13g2_FILL8
XSTDFILL22_2027 VDD VSS sg13g2_FILL8
XSTDFILL22_2035 VDD VSS sg13g2_FILL8
XSTDFILL22_2043 VDD VSS sg13g2_FILL8
XSTDFILL22_2051 VDD VSS sg13g2_FILL8
XSTDFILL22_2059 VDD VSS sg13g2_FILL8
XSTDFILL22_2067 VDD VSS sg13g2_FILL8
XSTDFILL22_2075 VDD VSS sg13g2_FILL8
XSTDFILL22_2083 VDD VSS sg13g2_FILL8
XSTDFILL22_2091 VDD VSS sg13g2_FILL8
XSTDFILL22_2099 VDD VSS sg13g2_FILL8
XSTDFILL22_2107 VDD VSS sg13g2_FILL8
XSTDFILL22_2115 VDD VSS sg13g2_FILL8
XSTDFILL22_2123 VDD VSS sg13g2_FILL8
XSTDFILL22_2131 VDD VSS sg13g2_FILL8
XSTDFILL22_2139 VDD VSS sg13g2_FILL8
XSTDFILL22_2147 VDD VSS sg13g2_FILL4
XSTDFILL22_2151 VDD VSS sg13g2_FILL2
XSTDFILL22_2153 VDD VSS sg13g2_FILL1
XSTDFILL23_0 VDD VSS sg13g2_FILL8
XSTDFILL23_8 VDD VSS sg13g2_FILL8
XSTDFILL23_16 VDD VSS sg13g2_FILL8
XSTDFILL23_24 VDD VSS sg13g2_FILL8
XSTDFILL23_32 VDD VSS sg13g2_FILL8
XSTDFILL23_40 VDD VSS sg13g2_FILL8
XSTDFILL23_48 VDD VSS sg13g2_FILL8
XSTDFILL23_56 VDD VSS sg13g2_FILL8
XSTDFILL23_64 VDD VSS sg13g2_FILL8
XSTDFILL23_72 VDD VSS sg13g2_FILL8
XSTDFILL23_80 VDD VSS sg13g2_FILL8
XSTDFILL23_88 VDD VSS sg13g2_FILL8
XSTDFILL23_96 VDD VSS sg13g2_FILL8
XSTDFILL23_104 VDD VSS sg13g2_FILL8
XSTDFILL23_112 VDD VSS sg13g2_FILL8
XSTDFILL23_120 VDD VSS sg13g2_FILL8
XSTDFILL23_128 VDD VSS sg13g2_FILL4
XSTDFILL23_1835 VDD VSS sg13g2_FILL8
XSTDFILL23_1843 VDD VSS sg13g2_FILL8
XSTDFILL23_1851 VDD VSS sg13g2_FILL8
XSTDFILL23_1859 VDD VSS sg13g2_FILL8
XSTDFILL23_1867 VDD VSS sg13g2_FILL8
XSTDFILL23_1875 VDD VSS sg13g2_FILL8
XSTDFILL23_1883 VDD VSS sg13g2_FILL8
XSTDFILL23_1891 VDD VSS sg13g2_FILL8
XSTDFILL23_1899 VDD VSS sg13g2_FILL8
XSTDFILL23_1907 VDD VSS sg13g2_FILL8
XSTDFILL23_1915 VDD VSS sg13g2_FILL8
XSTDFILL23_1923 VDD VSS sg13g2_FILL8
XSTDFILL23_1931 VDD VSS sg13g2_FILL8
XSTDFILL23_1939 VDD VSS sg13g2_FILL8
XSTDFILL23_1947 VDD VSS sg13g2_FILL8
XSTDFILL23_1955 VDD VSS sg13g2_FILL8
XSTDFILL23_1963 VDD VSS sg13g2_FILL8
XSTDFILL23_1971 VDD VSS sg13g2_FILL8
XSTDFILL23_1979 VDD VSS sg13g2_FILL8
XSTDFILL23_1987 VDD VSS sg13g2_FILL8
XSTDFILL23_1995 VDD VSS sg13g2_FILL8
XSTDFILL23_2003 VDD VSS sg13g2_FILL8
XSTDFILL23_2011 VDD VSS sg13g2_FILL8
XSTDFILL23_2019 VDD VSS sg13g2_FILL8
XSTDFILL23_2027 VDD VSS sg13g2_FILL8
XSTDFILL23_2035 VDD VSS sg13g2_FILL8
XSTDFILL23_2043 VDD VSS sg13g2_FILL8
XSTDFILL23_2051 VDD VSS sg13g2_FILL8
XSTDFILL23_2059 VDD VSS sg13g2_FILL8
XSTDFILL23_2067 VDD VSS sg13g2_FILL8
XSTDFILL23_2075 VDD VSS sg13g2_FILL8
XSTDFILL23_2083 VDD VSS sg13g2_FILL8
XSTDFILL23_2091 VDD VSS sg13g2_FILL8
XSTDFILL23_2099 VDD VSS sg13g2_FILL8
XSTDFILL23_2107 VDD VSS sg13g2_FILL8
XSTDFILL23_2115 VDD VSS sg13g2_FILL8
XSTDFILL23_2123 VDD VSS sg13g2_FILL8
XSTDFILL23_2131 VDD VSS sg13g2_FILL8
XSTDFILL23_2139 VDD VSS sg13g2_FILL8
XSTDFILL23_2147 VDD VSS sg13g2_FILL4
XSTDFILL23_2151 VDD VSS sg13g2_FILL2
XSTDFILL23_2153 VDD VSS sg13g2_FILL1
XSTDFILL24_0 VDD VSS sg13g2_FILL8
XSTDFILL24_8 VDD VSS sg13g2_FILL8
XSTDFILL24_16 VDD VSS sg13g2_FILL8
XSTDFILL24_24 VDD VSS sg13g2_FILL8
XSTDFILL24_32 VDD VSS sg13g2_FILL8
XSTDFILL24_40 VDD VSS sg13g2_FILL8
XSTDFILL24_48 VDD VSS sg13g2_FILL8
XSTDFILL24_56 VDD VSS sg13g2_FILL8
XSTDFILL24_64 VDD VSS sg13g2_FILL8
XSTDFILL24_72 VDD VSS sg13g2_FILL8
XSTDFILL24_80 VDD VSS sg13g2_FILL8
XSTDFILL24_88 VDD VSS sg13g2_FILL8
XSTDFILL24_96 VDD VSS sg13g2_FILL8
XSTDFILL24_104 VDD VSS sg13g2_FILL8
XSTDFILL24_112 VDD VSS sg13g2_FILL8
XSTDFILL24_120 VDD VSS sg13g2_FILL8
XSTDFILL24_128 VDD VSS sg13g2_FILL4
XSTDFILL24_1835 VDD VSS sg13g2_FILL8
XSTDFILL24_1843 VDD VSS sg13g2_FILL8
XSTDFILL24_1851 VDD VSS sg13g2_FILL8
XSTDFILL24_1859 VDD VSS sg13g2_FILL8
XSTDFILL24_1867 VDD VSS sg13g2_FILL8
XSTDFILL24_1875 VDD VSS sg13g2_FILL8
XSTDFILL24_1883 VDD VSS sg13g2_FILL8
XSTDFILL24_1891 VDD VSS sg13g2_FILL8
XSTDFILL24_1899 VDD VSS sg13g2_FILL8
XSTDFILL24_1907 VDD VSS sg13g2_FILL8
XSTDFILL24_1915 VDD VSS sg13g2_FILL8
XSTDFILL24_1923 VDD VSS sg13g2_FILL8
XSTDFILL24_1931 VDD VSS sg13g2_FILL8
XSTDFILL24_1939 VDD VSS sg13g2_FILL8
XSTDFILL24_1947 VDD VSS sg13g2_FILL8
XSTDFILL24_1955 VDD VSS sg13g2_FILL8
XSTDFILL24_1963 VDD VSS sg13g2_FILL8
XSTDFILL24_1971 VDD VSS sg13g2_FILL8
XSTDFILL24_1979 VDD VSS sg13g2_FILL8
XSTDFILL24_1987 VDD VSS sg13g2_FILL8
XSTDFILL24_1995 VDD VSS sg13g2_FILL8
XSTDFILL24_2003 VDD VSS sg13g2_FILL8
XSTDFILL24_2011 VDD VSS sg13g2_FILL8
XSTDFILL24_2019 VDD VSS sg13g2_FILL8
XSTDFILL24_2027 VDD VSS sg13g2_FILL8
XSTDFILL24_2035 VDD VSS sg13g2_FILL8
XSTDFILL24_2043 VDD VSS sg13g2_FILL8
XSTDFILL24_2051 VDD VSS sg13g2_FILL8
XSTDFILL24_2059 VDD VSS sg13g2_FILL8
XSTDFILL24_2067 VDD VSS sg13g2_FILL8
XSTDFILL24_2075 VDD VSS sg13g2_FILL8
XSTDFILL24_2083 VDD VSS sg13g2_FILL8
XSTDFILL24_2091 VDD VSS sg13g2_FILL8
XSTDFILL24_2099 VDD VSS sg13g2_FILL8
XSTDFILL24_2107 VDD VSS sg13g2_FILL8
XSTDFILL24_2115 VDD VSS sg13g2_FILL8
XSTDFILL24_2123 VDD VSS sg13g2_FILL8
XSTDFILL24_2131 VDD VSS sg13g2_FILL8
XSTDFILL24_2139 VDD VSS sg13g2_FILL8
XSTDFILL24_2147 VDD VSS sg13g2_FILL4
XSTDFILL24_2151 VDD VSS sg13g2_FILL2
XSTDFILL24_2153 VDD VSS sg13g2_FILL1
XSTDFILL25_0 VDD VSS sg13g2_FILL8
XSTDFILL25_8 VDD VSS sg13g2_FILL8
XSTDFILL25_16 VDD VSS sg13g2_FILL8
XSTDFILL25_24 VDD VSS sg13g2_FILL8
XSTDFILL25_32 VDD VSS sg13g2_FILL8
XSTDFILL25_40 VDD VSS sg13g2_FILL8
XSTDFILL25_48 VDD VSS sg13g2_FILL8
XSTDFILL25_56 VDD VSS sg13g2_FILL8
XSTDFILL25_64 VDD VSS sg13g2_FILL8
XSTDFILL25_72 VDD VSS sg13g2_FILL8
XSTDFILL25_80 VDD VSS sg13g2_FILL8
XSTDFILL25_88 VDD VSS sg13g2_FILL8
XSTDFILL25_96 VDD VSS sg13g2_FILL8
XSTDFILL25_104 VDD VSS sg13g2_FILL8
XSTDFILL25_112 VDD VSS sg13g2_FILL8
XSTDFILL25_120 VDD VSS sg13g2_FILL8
XSTDFILL25_128 VDD VSS sg13g2_FILL4
XSTDFILL25_1835 VDD VSS sg13g2_FILL8
XSTDFILL25_1843 VDD VSS sg13g2_FILL8
XSTDFILL25_1851 VDD VSS sg13g2_FILL8
XSTDFILL25_1859 VDD VSS sg13g2_FILL8
XSTDFILL25_1867 VDD VSS sg13g2_FILL8
XSTDFILL25_1875 VDD VSS sg13g2_FILL8
XSTDFILL25_1883 VDD VSS sg13g2_FILL8
XSTDFILL25_1891 VDD VSS sg13g2_FILL8
XSTDFILL25_1899 VDD VSS sg13g2_FILL8
XSTDFILL25_1907 VDD VSS sg13g2_FILL8
XSTDFILL25_1915 VDD VSS sg13g2_FILL8
XSTDFILL25_1923 VDD VSS sg13g2_FILL8
XSTDFILL25_1931 VDD VSS sg13g2_FILL8
XSTDFILL25_1939 VDD VSS sg13g2_FILL8
XSTDFILL25_1947 VDD VSS sg13g2_FILL8
XSTDFILL25_1955 VDD VSS sg13g2_FILL8
XSTDFILL25_1963 VDD VSS sg13g2_FILL8
XSTDFILL25_1971 VDD VSS sg13g2_FILL8
XSTDFILL25_1979 VDD VSS sg13g2_FILL8
XSTDFILL25_1987 VDD VSS sg13g2_FILL8
XSTDFILL25_1995 VDD VSS sg13g2_FILL8
XSTDFILL25_2003 VDD VSS sg13g2_FILL8
XSTDFILL25_2011 VDD VSS sg13g2_FILL8
XSTDFILL25_2019 VDD VSS sg13g2_FILL8
XSTDFILL25_2027 VDD VSS sg13g2_FILL8
XSTDFILL25_2035 VDD VSS sg13g2_FILL8
XSTDFILL25_2043 VDD VSS sg13g2_FILL8
XSTDFILL25_2051 VDD VSS sg13g2_FILL8
XSTDFILL25_2059 VDD VSS sg13g2_FILL8
XSTDFILL25_2067 VDD VSS sg13g2_FILL8
XSTDFILL25_2075 VDD VSS sg13g2_FILL8
XSTDFILL25_2083 VDD VSS sg13g2_FILL8
XSTDFILL25_2091 VDD VSS sg13g2_FILL8
XSTDFILL25_2099 VDD VSS sg13g2_FILL8
XSTDFILL25_2107 VDD VSS sg13g2_FILL8
XSTDFILL25_2115 VDD VSS sg13g2_FILL8
XSTDFILL25_2123 VDD VSS sg13g2_FILL8
XSTDFILL25_2131 VDD VSS sg13g2_FILL8
XSTDFILL25_2139 VDD VSS sg13g2_FILL8
XSTDFILL25_2147 VDD VSS sg13g2_FILL4
XSTDFILL25_2151 VDD VSS sg13g2_FILL2
XSTDFILL25_2153 VDD VSS sg13g2_FILL1
XSTDFILL26_0 VDD VSS sg13g2_FILL8
XSTDFILL26_8 VDD VSS sg13g2_FILL8
XSTDFILL26_16 VDD VSS sg13g2_FILL8
XSTDFILL26_24 VDD VSS sg13g2_FILL8
XSTDFILL26_32 VDD VSS sg13g2_FILL8
XSTDFILL26_40 VDD VSS sg13g2_FILL8
XSTDFILL26_48 VDD VSS sg13g2_FILL8
XSTDFILL26_56 VDD VSS sg13g2_FILL8
XSTDFILL26_64 VDD VSS sg13g2_FILL8
XSTDFILL26_72 VDD VSS sg13g2_FILL8
XSTDFILL26_80 VDD VSS sg13g2_FILL8
XSTDFILL26_88 VDD VSS sg13g2_FILL8
XSTDFILL26_96 VDD VSS sg13g2_FILL8
XSTDFILL26_104 VDD VSS sg13g2_FILL8
XSTDFILL26_112 VDD VSS sg13g2_FILL8
XSTDFILL26_120 VDD VSS sg13g2_FILL8
XSTDFILL26_128 VDD VSS sg13g2_FILL4
XSTDFILL26_1835 VDD VSS sg13g2_FILL8
XSTDFILL26_1843 VDD VSS sg13g2_FILL8
XSTDFILL26_1851 VDD VSS sg13g2_FILL8
XSTDFILL26_1859 VDD VSS sg13g2_FILL8
XSTDFILL26_1867 VDD VSS sg13g2_FILL8
XSTDFILL26_1875 VDD VSS sg13g2_FILL8
XSTDFILL26_1883 VDD VSS sg13g2_FILL8
XSTDFILL26_1891 VDD VSS sg13g2_FILL8
XSTDFILL26_1899 VDD VSS sg13g2_FILL8
XSTDFILL26_1907 VDD VSS sg13g2_FILL8
XSTDFILL26_1915 VDD VSS sg13g2_FILL8
XSTDFILL26_1923 VDD VSS sg13g2_FILL8
XSTDFILL26_1931 VDD VSS sg13g2_FILL8
XSTDFILL26_1939 VDD VSS sg13g2_FILL8
XSTDFILL26_1947 VDD VSS sg13g2_FILL8
XSTDFILL26_1955 VDD VSS sg13g2_FILL8
XSTDFILL26_1963 VDD VSS sg13g2_FILL8
XSTDFILL26_1971 VDD VSS sg13g2_FILL8
XSTDFILL26_1979 VDD VSS sg13g2_FILL8
XSTDFILL26_1987 VDD VSS sg13g2_FILL8
XSTDFILL26_1995 VDD VSS sg13g2_FILL8
XSTDFILL26_2003 VDD VSS sg13g2_FILL8
XSTDFILL26_2011 VDD VSS sg13g2_FILL8
XSTDFILL26_2019 VDD VSS sg13g2_FILL8
XSTDFILL26_2027 VDD VSS sg13g2_FILL8
XSTDFILL26_2035 VDD VSS sg13g2_FILL8
XSTDFILL26_2043 VDD VSS sg13g2_FILL8
XSTDFILL26_2051 VDD VSS sg13g2_FILL8
XSTDFILL26_2059 VDD VSS sg13g2_FILL8
XSTDFILL26_2067 VDD VSS sg13g2_FILL8
XSTDFILL26_2075 VDD VSS sg13g2_FILL8
XSTDFILL26_2083 VDD VSS sg13g2_FILL8
XSTDFILL26_2091 VDD VSS sg13g2_FILL8
XSTDFILL26_2099 VDD VSS sg13g2_FILL8
XSTDFILL26_2107 VDD VSS sg13g2_FILL8
XSTDFILL26_2115 VDD VSS sg13g2_FILL8
XSTDFILL26_2123 VDD VSS sg13g2_FILL8
XSTDFILL26_2131 VDD VSS sg13g2_FILL8
XSTDFILL26_2139 VDD VSS sg13g2_FILL8
XSTDFILL26_2147 VDD VSS sg13g2_FILL4
XSTDFILL26_2151 VDD VSS sg13g2_FILL2
XSTDFILL26_2153 VDD VSS sg13g2_FILL1
XSTDFILL27_0 VDD VSS sg13g2_FILL8
XSTDFILL27_8 VDD VSS sg13g2_FILL8
XSTDFILL27_16 VDD VSS sg13g2_FILL8
XSTDFILL27_24 VDD VSS sg13g2_FILL8
XSTDFILL27_32 VDD VSS sg13g2_FILL8
XSTDFILL27_40 VDD VSS sg13g2_FILL8
XSTDFILL27_48 VDD VSS sg13g2_FILL8
XSTDFILL27_56 VDD VSS sg13g2_FILL8
XSTDFILL27_64 VDD VSS sg13g2_FILL8
XSTDFILL27_72 VDD VSS sg13g2_FILL8
XSTDFILL27_80 VDD VSS sg13g2_FILL8
XSTDFILL27_88 VDD VSS sg13g2_FILL8
XSTDFILL27_96 VDD VSS sg13g2_FILL8
XSTDFILL27_104 VDD VSS sg13g2_FILL8
XSTDFILL27_112 VDD VSS sg13g2_FILL8
XSTDFILL27_120 VDD VSS sg13g2_FILL8
XSTDFILL27_128 VDD VSS sg13g2_FILL4
XSTDFILL27_1835 VDD VSS sg13g2_FILL8
XSTDFILL27_1843 VDD VSS sg13g2_FILL8
XSTDFILL27_1851 VDD VSS sg13g2_FILL8
XSTDFILL27_1859 VDD VSS sg13g2_FILL8
XSTDFILL27_1867 VDD VSS sg13g2_FILL8
XSTDFILL27_1875 VDD VSS sg13g2_FILL8
XSTDFILL27_1883 VDD VSS sg13g2_FILL8
XSTDFILL27_1891 VDD VSS sg13g2_FILL8
XSTDFILL27_1899 VDD VSS sg13g2_FILL8
XSTDFILL27_1907 VDD VSS sg13g2_FILL8
XSTDFILL27_1915 VDD VSS sg13g2_FILL8
XSTDFILL27_1923 VDD VSS sg13g2_FILL8
XSTDFILL27_1931 VDD VSS sg13g2_FILL8
XSTDFILL27_1939 VDD VSS sg13g2_FILL8
XSTDFILL27_1947 VDD VSS sg13g2_FILL8
XSTDFILL27_1955 VDD VSS sg13g2_FILL8
XSTDFILL27_1963 VDD VSS sg13g2_FILL8
XSTDFILL27_1971 VDD VSS sg13g2_FILL8
XSTDFILL27_1979 VDD VSS sg13g2_FILL8
XSTDFILL27_1987 VDD VSS sg13g2_FILL8
XSTDFILL27_1995 VDD VSS sg13g2_FILL8
XSTDFILL27_2003 VDD VSS sg13g2_FILL8
XSTDFILL27_2011 VDD VSS sg13g2_FILL8
XSTDFILL27_2019 VDD VSS sg13g2_FILL8
XSTDFILL27_2027 VDD VSS sg13g2_FILL8
XSTDFILL27_2035 VDD VSS sg13g2_FILL8
XSTDFILL27_2043 VDD VSS sg13g2_FILL8
XSTDFILL27_2051 VDD VSS sg13g2_FILL8
XSTDFILL27_2059 VDD VSS sg13g2_FILL8
XSTDFILL27_2067 VDD VSS sg13g2_FILL8
XSTDFILL27_2075 VDD VSS sg13g2_FILL8
XSTDFILL27_2083 VDD VSS sg13g2_FILL8
XSTDFILL27_2091 VDD VSS sg13g2_FILL8
XSTDFILL27_2099 VDD VSS sg13g2_FILL8
XSTDFILL27_2107 VDD VSS sg13g2_FILL8
XSTDFILL27_2115 VDD VSS sg13g2_FILL8
XSTDFILL27_2123 VDD VSS sg13g2_FILL8
XSTDFILL27_2131 VDD VSS sg13g2_FILL8
XSTDFILL27_2139 VDD VSS sg13g2_FILL8
XSTDFILL27_2147 VDD VSS sg13g2_FILL4
XSTDFILL27_2151 VDD VSS sg13g2_FILL2
XSTDFILL27_2153 VDD VSS sg13g2_FILL1
XSTDFILL28_0 VDD VSS sg13g2_FILL8
XSTDFILL28_8 VDD VSS sg13g2_FILL8
XSTDFILL28_16 VDD VSS sg13g2_FILL8
XSTDFILL28_24 VDD VSS sg13g2_FILL8
XSTDFILL28_32 VDD VSS sg13g2_FILL8
XSTDFILL28_40 VDD VSS sg13g2_FILL8
XSTDFILL28_48 VDD VSS sg13g2_FILL8
XSTDFILL28_56 VDD VSS sg13g2_FILL8
XSTDFILL28_64 VDD VSS sg13g2_FILL8
XSTDFILL28_72 VDD VSS sg13g2_FILL8
XSTDFILL28_80 VDD VSS sg13g2_FILL8
XSTDFILL28_88 VDD VSS sg13g2_FILL8
XSTDFILL28_96 VDD VSS sg13g2_FILL8
XSTDFILL28_104 VDD VSS sg13g2_FILL8
XSTDFILL28_112 VDD VSS sg13g2_FILL8
XSTDFILL28_120 VDD VSS sg13g2_FILL8
XSTDFILL28_128 VDD VSS sg13g2_FILL4
XSTDFILL28_1835 VDD VSS sg13g2_FILL8
XSTDFILL28_1843 VDD VSS sg13g2_FILL8
XSTDFILL28_1851 VDD VSS sg13g2_FILL8
XSTDFILL28_1859 VDD VSS sg13g2_FILL8
XSTDFILL28_1867 VDD VSS sg13g2_FILL8
XSTDFILL28_1875 VDD VSS sg13g2_FILL8
XSTDFILL28_1883 VDD VSS sg13g2_FILL8
XSTDFILL28_1891 VDD VSS sg13g2_FILL8
XSTDFILL28_1899 VDD VSS sg13g2_FILL8
XSTDFILL28_1907 VDD VSS sg13g2_FILL8
XSTDFILL28_1915 VDD VSS sg13g2_FILL8
XSTDFILL28_1923 VDD VSS sg13g2_FILL8
XSTDFILL28_1931 VDD VSS sg13g2_FILL8
XSTDFILL28_1939 VDD VSS sg13g2_FILL8
XSTDFILL28_1947 VDD VSS sg13g2_FILL8
XSTDFILL28_1955 VDD VSS sg13g2_FILL8
XSTDFILL28_1963 VDD VSS sg13g2_FILL8
XSTDFILL28_1971 VDD VSS sg13g2_FILL8
XSTDFILL28_1979 VDD VSS sg13g2_FILL8
XSTDFILL28_1987 VDD VSS sg13g2_FILL8
XSTDFILL28_1995 VDD VSS sg13g2_FILL8
XSTDFILL28_2003 VDD VSS sg13g2_FILL8
XSTDFILL28_2011 VDD VSS sg13g2_FILL8
XSTDFILL28_2019 VDD VSS sg13g2_FILL8
XSTDFILL28_2027 VDD VSS sg13g2_FILL8
XSTDFILL28_2035 VDD VSS sg13g2_FILL8
XSTDFILL28_2043 VDD VSS sg13g2_FILL8
XSTDFILL28_2051 VDD VSS sg13g2_FILL8
XSTDFILL28_2059 VDD VSS sg13g2_FILL8
XSTDFILL28_2067 VDD VSS sg13g2_FILL8
XSTDFILL28_2075 VDD VSS sg13g2_FILL8
XSTDFILL28_2083 VDD VSS sg13g2_FILL8
XSTDFILL28_2091 VDD VSS sg13g2_FILL8
XSTDFILL28_2099 VDD VSS sg13g2_FILL8
XSTDFILL28_2107 VDD VSS sg13g2_FILL8
XSTDFILL28_2115 VDD VSS sg13g2_FILL8
XSTDFILL28_2123 VDD VSS sg13g2_FILL8
XSTDFILL28_2131 VDD VSS sg13g2_FILL8
XSTDFILL28_2139 VDD VSS sg13g2_FILL8
XSTDFILL28_2147 VDD VSS sg13g2_FILL4
XSTDFILL28_2151 VDD VSS sg13g2_FILL2
XSTDFILL28_2153 VDD VSS sg13g2_FILL1
XSTDFILL29_0 VDD VSS sg13g2_FILL8
XSTDFILL29_8 VDD VSS sg13g2_FILL8
XSTDFILL29_16 VDD VSS sg13g2_FILL8
XSTDFILL29_24 VDD VSS sg13g2_FILL8
XSTDFILL29_32 VDD VSS sg13g2_FILL8
XSTDFILL29_40 VDD VSS sg13g2_FILL8
XSTDFILL29_48 VDD VSS sg13g2_FILL8
XSTDFILL29_56 VDD VSS sg13g2_FILL8
XSTDFILL29_64 VDD VSS sg13g2_FILL8
XSTDFILL29_72 VDD VSS sg13g2_FILL8
XSTDFILL29_80 VDD VSS sg13g2_FILL8
XSTDFILL29_88 VDD VSS sg13g2_FILL8
XSTDFILL29_96 VDD VSS sg13g2_FILL8
XSTDFILL29_104 VDD VSS sg13g2_FILL8
XSTDFILL29_112 VDD VSS sg13g2_FILL8
XSTDFILL29_120 VDD VSS sg13g2_FILL8
XSTDFILL29_128 VDD VSS sg13g2_FILL4
XSTDFILL29_1835 VDD VSS sg13g2_FILL8
XSTDFILL29_1843 VDD VSS sg13g2_FILL8
XSTDFILL29_1851 VDD VSS sg13g2_FILL8
XSTDFILL29_1859 VDD VSS sg13g2_FILL8
XSTDFILL29_1867 VDD VSS sg13g2_FILL8
XSTDFILL29_1875 VDD VSS sg13g2_FILL8
XSTDFILL29_1883 VDD VSS sg13g2_FILL8
XSTDFILL29_1891 VDD VSS sg13g2_FILL8
XSTDFILL29_1899 VDD VSS sg13g2_FILL8
XSTDFILL29_1907 VDD VSS sg13g2_FILL8
XSTDFILL29_1915 VDD VSS sg13g2_FILL8
XSTDFILL29_1923 VDD VSS sg13g2_FILL8
XSTDFILL29_1931 VDD VSS sg13g2_FILL8
XSTDFILL29_1939 VDD VSS sg13g2_FILL8
XSTDFILL29_1947 VDD VSS sg13g2_FILL8
XSTDFILL29_1955 VDD VSS sg13g2_FILL8
XSTDFILL29_1963 VDD VSS sg13g2_FILL8
XSTDFILL29_1971 VDD VSS sg13g2_FILL8
XSTDFILL29_1979 VDD VSS sg13g2_FILL8
XSTDFILL29_1987 VDD VSS sg13g2_FILL8
XSTDFILL29_1995 VDD VSS sg13g2_FILL8
XSTDFILL29_2003 VDD VSS sg13g2_FILL8
XSTDFILL29_2011 VDD VSS sg13g2_FILL8
XSTDFILL29_2019 VDD VSS sg13g2_FILL8
XSTDFILL29_2027 VDD VSS sg13g2_FILL8
XSTDFILL29_2035 VDD VSS sg13g2_FILL8
XSTDFILL29_2043 VDD VSS sg13g2_FILL8
XSTDFILL29_2051 VDD VSS sg13g2_FILL8
XSTDFILL29_2059 VDD VSS sg13g2_FILL8
XSTDFILL29_2067 VDD VSS sg13g2_FILL8
XSTDFILL29_2075 VDD VSS sg13g2_FILL8
XSTDFILL29_2083 VDD VSS sg13g2_FILL8
XSTDFILL29_2091 VDD VSS sg13g2_FILL8
XSTDFILL29_2099 VDD VSS sg13g2_FILL8
XSTDFILL29_2107 VDD VSS sg13g2_FILL8
XSTDFILL29_2115 VDD VSS sg13g2_FILL8
XSTDFILL29_2123 VDD VSS sg13g2_FILL8
XSTDFILL29_2131 VDD VSS sg13g2_FILL8
XSTDFILL29_2139 VDD VSS sg13g2_FILL8
XSTDFILL29_2147 VDD VSS sg13g2_FILL4
XSTDFILL29_2151 VDD VSS sg13g2_FILL2
XSTDFILL29_2153 VDD VSS sg13g2_FILL1
XSTDFILL30_0 VDD VSS sg13g2_FILL8
XSTDFILL30_8 VDD VSS sg13g2_FILL8
XSTDFILL30_16 VDD VSS sg13g2_FILL8
XSTDFILL30_24 VDD VSS sg13g2_FILL8
XSTDFILL30_32 VDD VSS sg13g2_FILL8
XSTDFILL30_40 VDD VSS sg13g2_FILL8
XSTDFILL30_48 VDD VSS sg13g2_FILL8
XSTDFILL30_56 VDD VSS sg13g2_FILL8
XSTDFILL30_64 VDD VSS sg13g2_FILL8
XSTDFILL30_72 VDD VSS sg13g2_FILL8
XSTDFILL30_80 VDD VSS sg13g2_FILL8
XSTDFILL30_88 VDD VSS sg13g2_FILL8
XSTDFILL30_96 VDD VSS sg13g2_FILL8
XSTDFILL30_104 VDD VSS sg13g2_FILL8
XSTDFILL30_112 VDD VSS sg13g2_FILL8
XSTDFILL30_120 VDD VSS sg13g2_FILL8
XSTDFILL30_128 VDD VSS sg13g2_FILL4
XSTDFILL30_1835 VDD VSS sg13g2_FILL8
XSTDFILL30_1843 VDD VSS sg13g2_FILL8
XSTDFILL30_1851 VDD VSS sg13g2_FILL8
XSTDFILL30_1859 VDD VSS sg13g2_FILL8
XSTDFILL30_1867 VDD VSS sg13g2_FILL8
XSTDFILL30_1875 VDD VSS sg13g2_FILL8
XSTDFILL30_1883 VDD VSS sg13g2_FILL8
XSTDFILL30_1891 VDD VSS sg13g2_FILL8
XSTDFILL30_1899 VDD VSS sg13g2_FILL8
XSTDFILL30_1907 VDD VSS sg13g2_FILL8
XSTDFILL30_1915 VDD VSS sg13g2_FILL8
XSTDFILL30_1923 VDD VSS sg13g2_FILL8
XSTDFILL30_1931 VDD VSS sg13g2_FILL8
XSTDFILL30_1939 VDD VSS sg13g2_FILL8
XSTDFILL30_1947 VDD VSS sg13g2_FILL8
XSTDFILL30_1955 VDD VSS sg13g2_FILL8
XSTDFILL30_1963 VDD VSS sg13g2_FILL8
XSTDFILL30_1971 VDD VSS sg13g2_FILL8
XSTDFILL30_1979 VDD VSS sg13g2_FILL8
XSTDFILL30_1987 VDD VSS sg13g2_FILL8
XSTDFILL30_1995 VDD VSS sg13g2_FILL8
XSTDFILL30_2003 VDD VSS sg13g2_FILL8
XSTDFILL30_2011 VDD VSS sg13g2_FILL8
XSTDFILL30_2019 VDD VSS sg13g2_FILL8
XSTDFILL30_2027 VDD VSS sg13g2_FILL8
XSTDFILL30_2035 VDD VSS sg13g2_FILL8
XSTDFILL30_2043 VDD VSS sg13g2_FILL8
XSTDFILL30_2051 VDD VSS sg13g2_FILL8
XSTDFILL30_2059 VDD VSS sg13g2_FILL8
XSTDFILL30_2067 VDD VSS sg13g2_FILL8
XSTDFILL30_2075 VDD VSS sg13g2_FILL8
XSTDFILL30_2083 VDD VSS sg13g2_FILL8
XSTDFILL30_2091 VDD VSS sg13g2_FILL8
XSTDFILL30_2099 VDD VSS sg13g2_FILL8
XSTDFILL30_2107 VDD VSS sg13g2_FILL8
XSTDFILL30_2115 VDD VSS sg13g2_FILL8
XSTDFILL30_2123 VDD VSS sg13g2_FILL8
XSTDFILL30_2131 VDD VSS sg13g2_FILL8
XSTDFILL30_2139 VDD VSS sg13g2_FILL8
XSTDFILL30_2147 VDD VSS sg13g2_FILL4
XSTDFILL30_2151 VDD VSS sg13g2_FILL2
XSTDFILL30_2153 VDD VSS sg13g2_FILL1
XSTDFILL31_0 VDD VSS sg13g2_FILL8
XSTDFILL31_8 VDD VSS sg13g2_FILL8
XSTDFILL31_16 VDD VSS sg13g2_FILL8
XSTDFILL31_24 VDD VSS sg13g2_FILL8
XSTDFILL31_32 VDD VSS sg13g2_FILL8
XSTDFILL31_40 VDD VSS sg13g2_FILL8
XSTDFILL31_48 VDD VSS sg13g2_FILL8
XSTDFILL31_56 VDD VSS sg13g2_FILL8
XSTDFILL31_64 VDD VSS sg13g2_FILL8
XSTDFILL31_72 VDD VSS sg13g2_FILL8
XSTDFILL31_80 VDD VSS sg13g2_FILL8
XSTDFILL31_88 VDD VSS sg13g2_FILL8
XSTDFILL31_96 VDD VSS sg13g2_FILL8
XSTDFILL31_104 VDD VSS sg13g2_FILL8
XSTDFILL31_112 VDD VSS sg13g2_FILL8
XSTDFILL31_120 VDD VSS sg13g2_FILL8
XSTDFILL31_128 VDD VSS sg13g2_FILL4
XSTDFILL31_1835 VDD VSS sg13g2_FILL8
XSTDFILL31_1843 VDD VSS sg13g2_FILL8
XSTDFILL31_1851 VDD VSS sg13g2_FILL8
XSTDFILL31_1859 VDD VSS sg13g2_FILL8
XSTDFILL31_1867 VDD VSS sg13g2_FILL8
XSTDFILL31_1875 VDD VSS sg13g2_FILL8
XSTDFILL31_1883 VDD VSS sg13g2_FILL8
XSTDFILL31_1891 VDD VSS sg13g2_FILL8
XSTDFILL31_1899 VDD VSS sg13g2_FILL8
XSTDFILL31_1907 VDD VSS sg13g2_FILL8
XSTDFILL31_1915 VDD VSS sg13g2_FILL8
XSTDFILL31_1923 VDD VSS sg13g2_FILL8
XSTDFILL31_1931 VDD VSS sg13g2_FILL8
XSTDFILL31_1939 VDD VSS sg13g2_FILL8
XSTDFILL31_1947 VDD VSS sg13g2_FILL8
XSTDFILL31_1955 VDD VSS sg13g2_FILL8
XSTDFILL31_1963 VDD VSS sg13g2_FILL8
XSTDFILL31_1971 VDD VSS sg13g2_FILL8
XSTDFILL31_1979 VDD VSS sg13g2_FILL8
XSTDFILL31_1987 VDD VSS sg13g2_FILL8
XSTDFILL31_1995 VDD VSS sg13g2_FILL8
XSTDFILL31_2003 VDD VSS sg13g2_FILL8
XSTDFILL31_2011 VDD VSS sg13g2_FILL8
XSTDFILL31_2019 VDD VSS sg13g2_FILL8
XSTDFILL31_2027 VDD VSS sg13g2_FILL8
XSTDFILL31_2035 VDD VSS sg13g2_FILL8
XSTDFILL31_2043 VDD VSS sg13g2_FILL8
XSTDFILL31_2051 VDD VSS sg13g2_FILL8
XSTDFILL31_2059 VDD VSS sg13g2_FILL8
XSTDFILL31_2067 VDD VSS sg13g2_FILL8
XSTDFILL31_2075 VDD VSS sg13g2_FILL8
XSTDFILL31_2083 VDD VSS sg13g2_FILL8
XSTDFILL31_2091 VDD VSS sg13g2_FILL8
XSTDFILL31_2099 VDD VSS sg13g2_FILL8
XSTDFILL31_2107 VDD VSS sg13g2_FILL8
XSTDFILL31_2115 VDD VSS sg13g2_FILL8
XSTDFILL31_2123 VDD VSS sg13g2_FILL8
XSTDFILL31_2131 VDD VSS sg13g2_FILL8
XSTDFILL31_2139 VDD VSS sg13g2_FILL8
XSTDFILL31_2147 VDD VSS sg13g2_FILL4
XSTDFILL31_2151 VDD VSS sg13g2_FILL2
XSTDFILL31_2153 VDD VSS sg13g2_FILL1
XSTDFILL32_0 VDD VSS sg13g2_FILL8
XSTDFILL32_8 VDD VSS sg13g2_FILL8
XSTDFILL32_16 VDD VSS sg13g2_FILL8
XSTDFILL32_24 VDD VSS sg13g2_FILL8
XSTDFILL32_32 VDD VSS sg13g2_FILL8
XSTDFILL32_40 VDD VSS sg13g2_FILL8
XSTDFILL32_48 VDD VSS sg13g2_FILL8
XSTDFILL32_56 VDD VSS sg13g2_FILL8
XSTDFILL32_64 VDD VSS sg13g2_FILL8
XSTDFILL32_72 VDD VSS sg13g2_FILL8
XSTDFILL32_80 VDD VSS sg13g2_FILL8
XSTDFILL32_88 VDD VSS sg13g2_FILL8
XSTDFILL32_96 VDD VSS sg13g2_FILL8
XSTDFILL32_104 VDD VSS sg13g2_FILL8
XSTDFILL32_112 VDD VSS sg13g2_FILL8
XSTDFILL32_120 VDD VSS sg13g2_FILL8
XSTDFILL32_128 VDD VSS sg13g2_FILL4
XSTDFILL32_1835 VDD VSS sg13g2_FILL8
XSTDFILL32_1843 VDD VSS sg13g2_FILL8
XSTDFILL32_1851 VDD VSS sg13g2_FILL8
XSTDFILL32_1859 VDD VSS sg13g2_FILL8
XSTDFILL32_1867 VDD VSS sg13g2_FILL8
XSTDFILL32_1875 VDD VSS sg13g2_FILL8
XSTDFILL32_1883 VDD VSS sg13g2_FILL8
XSTDFILL32_1891 VDD VSS sg13g2_FILL8
XSTDFILL32_1899 VDD VSS sg13g2_FILL8
XSTDFILL32_1907 VDD VSS sg13g2_FILL8
XSTDFILL32_1915 VDD VSS sg13g2_FILL8
XSTDFILL32_1923 VDD VSS sg13g2_FILL8
XSTDFILL32_1931 VDD VSS sg13g2_FILL8
XSTDFILL32_1939 VDD VSS sg13g2_FILL8
XSTDFILL32_1947 VDD VSS sg13g2_FILL8
XSTDFILL32_1955 VDD VSS sg13g2_FILL8
XSTDFILL32_1963 VDD VSS sg13g2_FILL8
XSTDFILL32_1971 VDD VSS sg13g2_FILL8
XSTDFILL32_1979 VDD VSS sg13g2_FILL8
XSTDFILL32_1987 VDD VSS sg13g2_FILL8
XSTDFILL32_1995 VDD VSS sg13g2_FILL8
XSTDFILL32_2003 VDD VSS sg13g2_FILL8
XSTDFILL32_2011 VDD VSS sg13g2_FILL8
XSTDFILL32_2019 VDD VSS sg13g2_FILL8
XSTDFILL32_2027 VDD VSS sg13g2_FILL8
XSTDFILL32_2035 VDD VSS sg13g2_FILL8
XSTDFILL32_2043 VDD VSS sg13g2_FILL8
XSTDFILL32_2051 VDD VSS sg13g2_FILL8
XSTDFILL32_2059 VDD VSS sg13g2_FILL8
XSTDFILL32_2067 VDD VSS sg13g2_FILL8
XSTDFILL32_2075 VDD VSS sg13g2_FILL8
XSTDFILL32_2083 VDD VSS sg13g2_FILL8
XSTDFILL32_2091 VDD VSS sg13g2_FILL8
XSTDFILL32_2099 VDD VSS sg13g2_FILL8
XSTDFILL32_2107 VDD VSS sg13g2_FILL8
XSTDFILL32_2115 VDD VSS sg13g2_FILL8
XSTDFILL32_2123 VDD VSS sg13g2_FILL8
XSTDFILL32_2131 VDD VSS sg13g2_FILL8
XSTDFILL32_2139 VDD VSS sg13g2_FILL8
XSTDFILL32_2147 VDD VSS sg13g2_FILL4
XSTDFILL32_2151 VDD VSS sg13g2_FILL2
XSTDFILL32_2153 VDD VSS sg13g2_FILL1
XSTDFILL33_0 VDD VSS sg13g2_FILL8
XSTDFILL33_8 VDD VSS sg13g2_FILL8
XSTDFILL33_16 VDD VSS sg13g2_FILL8
XSTDFILL33_24 VDD VSS sg13g2_FILL8
XSTDFILL33_32 VDD VSS sg13g2_FILL8
XSTDFILL33_40 VDD VSS sg13g2_FILL8
XSTDFILL33_48 VDD VSS sg13g2_FILL8
XSTDFILL33_56 VDD VSS sg13g2_FILL8
XSTDFILL33_64 VDD VSS sg13g2_FILL8
XSTDFILL33_72 VDD VSS sg13g2_FILL8
XSTDFILL33_80 VDD VSS sg13g2_FILL8
XSTDFILL33_88 VDD VSS sg13g2_FILL8
XSTDFILL33_96 VDD VSS sg13g2_FILL8
XSTDFILL33_104 VDD VSS sg13g2_FILL8
XSTDFILL33_112 VDD VSS sg13g2_FILL8
XSTDFILL33_120 VDD VSS sg13g2_FILL8
XSTDFILL33_128 VDD VSS sg13g2_FILL4
XSTDFILL33_1835 VDD VSS sg13g2_FILL8
XSTDFILL33_1843 VDD VSS sg13g2_FILL8
XSTDFILL33_1851 VDD VSS sg13g2_FILL8
XSTDFILL33_1859 VDD VSS sg13g2_FILL8
XSTDFILL33_1867 VDD VSS sg13g2_FILL8
XSTDFILL33_1875 VDD VSS sg13g2_FILL8
XSTDFILL33_1883 VDD VSS sg13g2_FILL8
XSTDFILL33_1891 VDD VSS sg13g2_FILL8
XSTDFILL33_1899 VDD VSS sg13g2_FILL8
XSTDFILL33_1907 VDD VSS sg13g2_FILL8
XSTDFILL33_1915 VDD VSS sg13g2_FILL8
XSTDFILL33_1923 VDD VSS sg13g2_FILL8
XSTDFILL33_1931 VDD VSS sg13g2_FILL8
XSTDFILL33_1939 VDD VSS sg13g2_FILL8
XSTDFILL33_1947 VDD VSS sg13g2_FILL8
XSTDFILL33_1955 VDD VSS sg13g2_FILL8
XSTDFILL33_1963 VDD VSS sg13g2_FILL8
XSTDFILL33_1971 VDD VSS sg13g2_FILL8
XSTDFILL33_1979 VDD VSS sg13g2_FILL8
XSTDFILL33_1987 VDD VSS sg13g2_FILL8
XSTDFILL33_1995 VDD VSS sg13g2_FILL8
XSTDFILL33_2003 VDD VSS sg13g2_FILL8
XSTDFILL33_2011 VDD VSS sg13g2_FILL8
XSTDFILL33_2019 VDD VSS sg13g2_FILL8
XSTDFILL33_2027 VDD VSS sg13g2_FILL8
XSTDFILL33_2035 VDD VSS sg13g2_FILL8
XSTDFILL33_2043 VDD VSS sg13g2_FILL8
XSTDFILL33_2051 VDD VSS sg13g2_FILL8
XSTDFILL33_2059 VDD VSS sg13g2_FILL8
XSTDFILL33_2067 VDD VSS sg13g2_FILL8
XSTDFILL33_2075 VDD VSS sg13g2_FILL8
XSTDFILL33_2083 VDD VSS sg13g2_FILL8
XSTDFILL33_2091 VDD VSS sg13g2_FILL8
XSTDFILL33_2099 VDD VSS sg13g2_FILL8
XSTDFILL33_2107 VDD VSS sg13g2_FILL8
XSTDFILL33_2115 VDD VSS sg13g2_FILL8
XSTDFILL33_2123 VDD VSS sg13g2_FILL8
XSTDFILL33_2131 VDD VSS sg13g2_FILL8
XSTDFILL33_2139 VDD VSS sg13g2_FILL8
XSTDFILL33_2147 VDD VSS sg13g2_FILL4
XSTDFILL33_2151 VDD VSS sg13g2_FILL2
XSTDFILL33_2153 VDD VSS sg13g2_FILL1
XSTDFILL34_0 VDD VSS sg13g2_FILL8
XSTDFILL34_8 VDD VSS sg13g2_FILL8
XSTDFILL34_16 VDD VSS sg13g2_FILL8
XSTDFILL34_24 VDD VSS sg13g2_FILL8
XSTDFILL34_32 VDD VSS sg13g2_FILL8
XSTDFILL34_40 VDD VSS sg13g2_FILL8
XSTDFILL34_48 VDD VSS sg13g2_FILL8
XSTDFILL34_56 VDD VSS sg13g2_FILL8
XSTDFILL34_64 VDD VSS sg13g2_FILL8
XSTDFILL34_72 VDD VSS sg13g2_FILL8
XSTDFILL34_80 VDD VSS sg13g2_FILL8
XSTDFILL34_88 VDD VSS sg13g2_FILL8
XSTDFILL34_96 VDD VSS sg13g2_FILL8
XSTDFILL34_104 VDD VSS sg13g2_FILL8
XSTDFILL34_112 VDD VSS sg13g2_FILL8
XSTDFILL34_120 VDD VSS sg13g2_FILL8
XSTDFILL34_128 VDD VSS sg13g2_FILL4
XSTDFILL34_1835 VDD VSS sg13g2_FILL8
XSTDFILL34_1843 VDD VSS sg13g2_FILL8
XSTDFILL34_1851 VDD VSS sg13g2_FILL8
XSTDFILL34_1859 VDD VSS sg13g2_FILL8
XSTDFILL34_1867 VDD VSS sg13g2_FILL8
XSTDFILL34_1875 VDD VSS sg13g2_FILL8
XSTDFILL34_1883 VDD VSS sg13g2_FILL8
XSTDFILL34_1891 VDD VSS sg13g2_FILL8
XSTDFILL34_1899 VDD VSS sg13g2_FILL8
XSTDFILL34_1907 VDD VSS sg13g2_FILL8
XSTDFILL34_1915 VDD VSS sg13g2_FILL8
XSTDFILL34_1923 VDD VSS sg13g2_FILL8
XSTDFILL34_1931 VDD VSS sg13g2_FILL8
XSTDFILL34_1939 VDD VSS sg13g2_FILL8
XSTDFILL34_1947 VDD VSS sg13g2_FILL8
XSTDFILL34_1955 VDD VSS sg13g2_FILL8
XSTDFILL34_1963 VDD VSS sg13g2_FILL8
XSTDFILL34_1971 VDD VSS sg13g2_FILL8
XSTDFILL34_1979 VDD VSS sg13g2_FILL8
XSTDFILL34_1987 VDD VSS sg13g2_FILL8
XSTDFILL34_1995 VDD VSS sg13g2_FILL8
XSTDFILL34_2003 VDD VSS sg13g2_FILL8
XSTDFILL34_2011 VDD VSS sg13g2_FILL8
XSTDFILL34_2019 VDD VSS sg13g2_FILL8
XSTDFILL34_2027 VDD VSS sg13g2_FILL8
XSTDFILL34_2035 VDD VSS sg13g2_FILL8
XSTDFILL34_2043 VDD VSS sg13g2_FILL8
XSTDFILL34_2051 VDD VSS sg13g2_FILL8
XSTDFILL34_2059 VDD VSS sg13g2_FILL8
XSTDFILL34_2067 VDD VSS sg13g2_FILL8
XSTDFILL34_2075 VDD VSS sg13g2_FILL8
XSTDFILL34_2083 VDD VSS sg13g2_FILL8
XSTDFILL34_2091 VDD VSS sg13g2_FILL8
XSTDFILL34_2099 VDD VSS sg13g2_FILL8
XSTDFILL34_2107 VDD VSS sg13g2_FILL8
XSTDFILL34_2115 VDD VSS sg13g2_FILL8
XSTDFILL34_2123 VDD VSS sg13g2_FILL8
XSTDFILL34_2131 VDD VSS sg13g2_FILL8
XSTDFILL34_2139 VDD VSS sg13g2_FILL8
XSTDFILL34_2147 VDD VSS sg13g2_FILL4
XSTDFILL34_2151 VDD VSS sg13g2_FILL2
XSTDFILL34_2153 VDD VSS sg13g2_FILL1
XSTDFILL35_0 VDD VSS sg13g2_FILL8
XSTDFILL35_8 VDD VSS sg13g2_FILL8
XSTDFILL35_16 VDD VSS sg13g2_FILL8
XSTDFILL35_24 VDD VSS sg13g2_FILL8
XSTDFILL35_32 VDD VSS sg13g2_FILL8
XSTDFILL35_40 VDD VSS sg13g2_FILL8
XSTDFILL35_48 VDD VSS sg13g2_FILL8
XSTDFILL35_56 VDD VSS sg13g2_FILL8
XSTDFILL35_64 VDD VSS sg13g2_FILL8
XSTDFILL35_72 VDD VSS sg13g2_FILL8
XSTDFILL35_80 VDD VSS sg13g2_FILL8
XSTDFILL35_88 VDD VSS sg13g2_FILL8
XSTDFILL35_96 VDD VSS sg13g2_FILL8
XSTDFILL35_104 VDD VSS sg13g2_FILL8
XSTDFILL35_112 VDD VSS sg13g2_FILL8
XSTDFILL35_120 VDD VSS sg13g2_FILL8
XSTDFILL35_128 VDD VSS sg13g2_FILL4
XSTDFILL35_1835 VDD VSS sg13g2_FILL8
XSTDFILL35_1843 VDD VSS sg13g2_FILL8
XSTDFILL35_1851 VDD VSS sg13g2_FILL8
XSTDFILL35_1859 VDD VSS sg13g2_FILL8
XSTDFILL35_1867 VDD VSS sg13g2_FILL8
XSTDFILL35_1875 VDD VSS sg13g2_FILL8
XSTDFILL35_1883 VDD VSS sg13g2_FILL8
XSTDFILL35_1891 VDD VSS sg13g2_FILL8
XSTDFILL35_1899 VDD VSS sg13g2_FILL8
XSTDFILL35_1907 VDD VSS sg13g2_FILL8
XSTDFILL35_1915 VDD VSS sg13g2_FILL8
XSTDFILL35_1923 VDD VSS sg13g2_FILL8
XSTDFILL35_1931 VDD VSS sg13g2_FILL8
XSTDFILL35_1939 VDD VSS sg13g2_FILL8
XSTDFILL35_1947 VDD VSS sg13g2_FILL8
XSTDFILL35_1955 VDD VSS sg13g2_FILL8
XSTDFILL35_1963 VDD VSS sg13g2_FILL8
XSTDFILL35_1971 VDD VSS sg13g2_FILL8
XSTDFILL35_1979 VDD VSS sg13g2_FILL8
XSTDFILL35_1987 VDD VSS sg13g2_FILL8
XSTDFILL35_1995 VDD VSS sg13g2_FILL8
XSTDFILL35_2003 VDD VSS sg13g2_FILL8
XSTDFILL35_2011 VDD VSS sg13g2_FILL8
XSTDFILL35_2019 VDD VSS sg13g2_FILL8
XSTDFILL35_2027 VDD VSS sg13g2_FILL8
XSTDFILL35_2035 VDD VSS sg13g2_FILL8
XSTDFILL35_2043 VDD VSS sg13g2_FILL8
XSTDFILL35_2051 VDD VSS sg13g2_FILL8
XSTDFILL35_2059 VDD VSS sg13g2_FILL8
XSTDFILL35_2067 VDD VSS sg13g2_FILL8
XSTDFILL35_2075 VDD VSS sg13g2_FILL8
XSTDFILL35_2083 VDD VSS sg13g2_FILL8
XSTDFILL35_2091 VDD VSS sg13g2_FILL8
XSTDFILL35_2099 VDD VSS sg13g2_FILL8
XSTDFILL35_2107 VDD VSS sg13g2_FILL8
XSTDFILL35_2115 VDD VSS sg13g2_FILL8
XSTDFILL35_2123 VDD VSS sg13g2_FILL8
XSTDFILL35_2131 VDD VSS sg13g2_FILL8
XSTDFILL35_2139 VDD VSS sg13g2_FILL8
XSTDFILL35_2147 VDD VSS sg13g2_FILL4
XSTDFILL35_2151 VDD VSS sg13g2_FILL2
XSTDFILL35_2153 VDD VSS sg13g2_FILL1
XSTDFILL36_0 VDD VSS sg13g2_FILL8
XSTDFILL36_8 VDD VSS sg13g2_FILL8
XSTDFILL36_16 VDD VSS sg13g2_FILL8
XSTDFILL36_24 VDD VSS sg13g2_FILL8
XSTDFILL36_32 VDD VSS sg13g2_FILL8
XSTDFILL36_40 VDD VSS sg13g2_FILL8
XSTDFILL36_48 VDD VSS sg13g2_FILL8
XSTDFILL36_56 VDD VSS sg13g2_FILL8
XSTDFILL36_64 VDD VSS sg13g2_FILL8
XSTDFILL36_72 VDD VSS sg13g2_FILL8
XSTDFILL36_80 VDD VSS sg13g2_FILL8
XSTDFILL36_88 VDD VSS sg13g2_FILL8
XSTDFILL36_96 VDD VSS sg13g2_FILL8
XSTDFILL36_104 VDD VSS sg13g2_FILL8
XSTDFILL36_112 VDD VSS sg13g2_FILL8
XSTDFILL36_120 VDD VSS sg13g2_FILL8
XSTDFILL36_128 VDD VSS sg13g2_FILL4
XSTDFILL36_1835 VDD VSS sg13g2_FILL8
XSTDFILL36_1843 VDD VSS sg13g2_FILL8
XSTDFILL36_1851 VDD VSS sg13g2_FILL8
XSTDFILL36_1859 VDD VSS sg13g2_FILL8
XSTDFILL36_1867 VDD VSS sg13g2_FILL8
XSTDFILL36_1875 VDD VSS sg13g2_FILL8
XSTDFILL36_1883 VDD VSS sg13g2_FILL8
XSTDFILL36_1891 VDD VSS sg13g2_FILL8
XSTDFILL36_1899 VDD VSS sg13g2_FILL8
XSTDFILL36_1907 VDD VSS sg13g2_FILL8
XSTDFILL36_1915 VDD VSS sg13g2_FILL8
XSTDFILL36_1923 VDD VSS sg13g2_FILL8
XSTDFILL36_1931 VDD VSS sg13g2_FILL8
XSTDFILL36_1939 VDD VSS sg13g2_FILL8
XSTDFILL36_1947 VDD VSS sg13g2_FILL8
XSTDFILL36_1955 VDD VSS sg13g2_FILL8
XSTDFILL36_1963 VDD VSS sg13g2_FILL8
XSTDFILL36_1971 VDD VSS sg13g2_FILL8
XSTDFILL36_1979 VDD VSS sg13g2_FILL8
XSTDFILL36_1987 VDD VSS sg13g2_FILL8
XSTDFILL36_1995 VDD VSS sg13g2_FILL8
XSTDFILL36_2003 VDD VSS sg13g2_FILL8
XSTDFILL36_2011 VDD VSS sg13g2_FILL8
XSTDFILL36_2019 VDD VSS sg13g2_FILL8
XSTDFILL36_2027 VDD VSS sg13g2_FILL8
XSTDFILL36_2035 VDD VSS sg13g2_FILL8
XSTDFILL36_2043 VDD VSS sg13g2_FILL8
XSTDFILL36_2051 VDD VSS sg13g2_FILL8
XSTDFILL36_2059 VDD VSS sg13g2_FILL8
XSTDFILL36_2067 VDD VSS sg13g2_FILL8
XSTDFILL36_2075 VDD VSS sg13g2_FILL8
XSTDFILL36_2083 VDD VSS sg13g2_FILL8
XSTDFILL36_2091 VDD VSS sg13g2_FILL8
XSTDFILL36_2099 VDD VSS sg13g2_FILL8
XSTDFILL36_2107 VDD VSS sg13g2_FILL8
XSTDFILL36_2115 VDD VSS sg13g2_FILL8
XSTDFILL36_2123 VDD VSS sg13g2_FILL8
XSTDFILL36_2131 VDD VSS sg13g2_FILL8
XSTDFILL36_2139 VDD VSS sg13g2_FILL8
XSTDFILL36_2147 VDD VSS sg13g2_FILL4
XSTDFILL36_2151 VDD VSS sg13g2_FILL2
XSTDFILL36_2153 VDD VSS sg13g2_FILL1
XSTDFILL37_0 VDD VSS sg13g2_FILL8
XSTDFILL37_8 VDD VSS sg13g2_FILL8
XSTDFILL37_16 VDD VSS sg13g2_FILL8
XSTDFILL37_24 VDD VSS sg13g2_FILL8
XSTDFILL37_32 VDD VSS sg13g2_FILL8
XSTDFILL37_40 VDD VSS sg13g2_FILL8
XSTDFILL37_48 VDD VSS sg13g2_FILL8
XSTDFILL37_56 VDD VSS sg13g2_FILL8
XSTDFILL37_64 VDD VSS sg13g2_FILL8
XSTDFILL37_72 VDD VSS sg13g2_FILL8
XSTDFILL37_80 VDD VSS sg13g2_FILL8
XSTDFILL37_88 VDD VSS sg13g2_FILL8
XSTDFILL37_96 VDD VSS sg13g2_FILL8
XSTDFILL37_104 VDD VSS sg13g2_FILL8
XSTDFILL37_112 VDD VSS sg13g2_FILL8
XSTDFILL37_120 VDD VSS sg13g2_FILL8
XSTDFILL37_128 VDD VSS sg13g2_FILL4
XSTDFILL37_1835 VDD VSS sg13g2_FILL8
XSTDFILL37_1843 VDD VSS sg13g2_FILL8
XSTDFILL37_1851 VDD VSS sg13g2_FILL8
XSTDFILL37_1859 VDD VSS sg13g2_FILL8
XSTDFILL37_1867 VDD VSS sg13g2_FILL8
XSTDFILL37_1875 VDD VSS sg13g2_FILL8
XSTDFILL37_1883 VDD VSS sg13g2_FILL8
XSTDFILL37_1891 VDD VSS sg13g2_FILL8
XSTDFILL37_1899 VDD VSS sg13g2_FILL8
XSTDFILL37_1907 VDD VSS sg13g2_FILL8
XSTDFILL37_1915 VDD VSS sg13g2_FILL8
XSTDFILL37_1923 VDD VSS sg13g2_FILL8
XSTDFILL37_1931 VDD VSS sg13g2_FILL8
XSTDFILL37_1939 VDD VSS sg13g2_FILL8
XSTDFILL37_1947 VDD VSS sg13g2_FILL8
XSTDFILL37_1955 VDD VSS sg13g2_FILL8
XSTDFILL37_1963 VDD VSS sg13g2_FILL8
XSTDFILL37_1971 VDD VSS sg13g2_FILL8
XSTDFILL37_1979 VDD VSS sg13g2_FILL8
XSTDFILL37_1987 VDD VSS sg13g2_FILL8
XSTDFILL37_1995 VDD VSS sg13g2_FILL8
XSTDFILL37_2003 VDD VSS sg13g2_FILL8
XSTDFILL37_2011 VDD VSS sg13g2_FILL8
XSTDFILL37_2019 VDD VSS sg13g2_FILL8
XSTDFILL37_2027 VDD VSS sg13g2_FILL8
XSTDFILL37_2035 VDD VSS sg13g2_FILL8
XSTDFILL37_2043 VDD VSS sg13g2_FILL8
XSTDFILL37_2051 VDD VSS sg13g2_FILL8
XSTDFILL37_2059 VDD VSS sg13g2_FILL8
XSTDFILL37_2067 VDD VSS sg13g2_FILL8
XSTDFILL37_2075 VDD VSS sg13g2_FILL8
XSTDFILL37_2083 VDD VSS sg13g2_FILL8
XSTDFILL37_2091 VDD VSS sg13g2_FILL8
XSTDFILL37_2099 VDD VSS sg13g2_FILL8
XSTDFILL37_2107 VDD VSS sg13g2_FILL8
XSTDFILL37_2115 VDD VSS sg13g2_FILL8
XSTDFILL37_2123 VDD VSS sg13g2_FILL8
XSTDFILL37_2131 VDD VSS sg13g2_FILL8
XSTDFILL37_2139 VDD VSS sg13g2_FILL8
XSTDFILL37_2147 VDD VSS sg13g2_FILL4
XSTDFILL37_2151 VDD VSS sg13g2_FILL2
XSTDFILL37_2153 VDD VSS sg13g2_FILL1
XSTDFILL38_0 VDD VSS sg13g2_FILL8
XSTDFILL38_8 VDD VSS sg13g2_FILL8
XSTDFILL38_16 VDD VSS sg13g2_FILL8
XSTDFILL38_24 VDD VSS sg13g2_FILL8
XSTDFILL38_32 VDD VSS sg13g2_FILL8
XSTDFILL38_40 VDD VSS sg13g2_FILL8
XSTDFILL38_48 VDD VSS sg13g2_FILL8
XSTDFILL38_56 VDD VSS sg13g2_FILL8
XSTDFILL38_64 VDD VSS sg13g2_FILL8
XSTDFILL38_72 VDD VSS sg13g2_FILL8
XSTDFILL38_80 VDD VSS sg13g2_FILL8
XSTDFILL38_88 VDD VSS sg13g2_FILL8
XSTDFILL38_96 VDD VSS sg13g2_FILL8
XSTDFILL38_104 VDD VSS sg13g2_FILL8
XSTDFILL38_112 VDD VSS sg13g2_FILL8
XSTDFILL38_120 VDD VSS sg13g2_FILL8
XSTDFILL38_128 VDD VSS sg13g2_FILL4
XSTDFILL38_1835 VDD VSS sg13g2_FILL8
XSTDFILL38_1843 VDD VSS sg13g2_FILL8
XSTDFILL38_1851 VDD VSS sg13g2_FILL8
XSTDFILL38_1859 VDD VSS sg13g2_FILL8
XSTDFILL38_1867 VDD VSS sg13g2_FILL8
XSTDFILL38_1875 VDD VSS sg13g2_FILL8
XSTDFILL38_1883 VDD VSS sg13g2_FILL8
XSTDFILL38_1891 VDD VSS sg13g2_FILL8
XSTDFILL38_1899 VDD VSS sg13g2_FILL8
XSTDFILL38_1907 VDD VSS sg13g2_FILL8
XSTDFILL38_1915 VDD VSS sg13g2_FILL8
XSTDFILL38_1923 VDD VSS sg13g2_FILL8
XSTDFILL38_1931 VDD VSS sg13g2_FILL8
XSTDFILL38_1939 VDD VSS sg13g2_FILL8
XSTDFILL38_1947 VDD VSS sg13g2_FILL8
XSTDFILL38_1955 VDD VSS sg13g2_FILL8
XSTDFILL38_1963 VDD VSS sg13g2_FILL8
XSTDFILL38_1971 VDD VSS sg13g2_FILL8
XSTDFILL38_1979 VDD VSS sg13g2_FILL8
XSTDFILL38_1987 VDD VSS sg13g2_FILL8
XSTDFILL38_1995 VDD VSS sg13g2_FILL8
XSTDFILL38_2003 VDD VSS sg13g2_FILL8
XSTDFILL38_2011 VDD VSS sg13g2_FILL8
XSTDFILL38_2019 VDD VSS sg13g2_FILL8
XSTDFILL38_2027 VDD VSS sg13g2_FILL8
XSTDFILL38_2035 VDD VSS sg13g2_FILL8
XSTDFILL38_2043 VDD VSS sg13g2_FILL8
XSTDFILL38_2051 VDD VSS sg13g2_FILL8
XSTDFILL38_2059 VDD VSS sg13g2_FILL8
XSTDFILL38_2067 VDD VSS sg13g2_FILL8
XSTDFILL38_2075 VDD VSS sg13g2_FILL8
XSTDFILL38_2083 VDD VSS sg13g2_FILL8
XSTDFILL38_2091 VDD VSS sg13g2_FILL8
XSTDFILL38_2099 VDD VSS sg13g2_FILL8
XSTDFILL38_2107 VDD VSS sg13g2_FILL8
XSTDFILL38_2115 VDD VSS sg13g2_FILL8
XSTDFILL38_2123 VDD VSS sg13g2_FILL8
XSTDFILL38_2131 VDD VSS sg13g2_FILL8
XSTDFILL38_2139 VDD VSS sg13g2_FILL8
XSTDFILL38_2147 VDD VSS sg13g2_FILL4
XSTDFILL38_2151 VDD VSS sg13g2_FILL2
XSTDFILL38_2153 VDD VSS sg13g2_FILL1
XSTDFILL39_0 VDD VSS sg13g2_FILL8
XSTDFILL39_8 VDD VSS sg13g2_FILL8
XSTDFILL39_16 VDD VSS sg13g2_FILL8
XSTDFILL39_24 VDD VSS sg13g2_FILL8
XSTDFILL39_32 VDD VSS sg13g2_FILL8
XSTDFILL39_40 VDD VSS sg13g2_FILL8
XSTDFILL39_48 VDD VSS sg13g2_FILL8
XSTDFILL39_56 VDD VSS sg13g2_FILL8
XSTDFILL39_64 VDD VSS sg13g2_FILL8
XSTDFILL39_72 VDD VSS sg13g2_FILL8
XSTDFILL39_80 VDD VSS sg13g2_FILL8
XSTDFILL39_88 VDD VSS sg13g2_FILL8
XSTDFILL39_96 VDD VSS sg13g2_FILL8
XSTDFILL39_104 VDD VSS sg13g2_FILL8
XSTDFILL39_112 VDD VSS sg13g2_FILL8
XSTDFILL39_120 VDD VSS sg13g2_FILL8
XSTDFILL39_128 VDD VSS sg13g2_FILL4
XSTDFILL39_1835 VDD VSS sg13g2_FILL8
XSTDFILL39_1843 VDD VSS sg13g2_FILL8
XSTDFILL39_1851 VDD VSS sg13g2_FILL8
XSTDFILL39_1859 VDD VSS sg13g2_FILL8
XSTDFILL39_1867 VDD VSS sg13g2_FILL8
XSTDFILL39_1875 VDD VSS sg13g2_FILL8
XSTDFILL39_1883 VDD VSS sg13g2_FILL8
XSTDFILL39_1891 VDD VSS sg13g2_FILL8
XSTDFILL39_1899 VDD VSS sg13g2_FILL8
XSTDFILL39_1907 VDD VSS sg13g2_FILL8
XSTDFILL39_1915 VDD VSS sg13g2_FILL8
XSTDFILL39_1923 VDD VSS sg13g2_FILL8
XSTDFILL39_1931 VDD VSS sg13g2_FILL8
XSTDFILL39_1939 VDD VSS sg13g2_FILL8
XSTDFILL39_1947 VDD VSS sg13g2_FILL8
XSTDFILL39_1955 VDD VSS sg13g2_FILL8
XSTDFILL39_1963 VDD VSS sg13g2_FILL8
XSTDFILL39_1971 VDD VSS sg13g2_FILL8
XSTDFILL39_1979 VDD VSS sg13g2_FILL8
XSTDFILL39_1987 VDD VSS sg13g2_FILL8
XSTDFILL39_1995 VDD VSS sg13g2_FILL8
XSTDFILL39_2003 VDD VSS sg13g2_FILL8
XSTDFILL39_2011 VDD VSS sg13g2_FILL8
XSTDFILL39_2019 VDD VSS sg13g2_FILL8
XSTDFILL39_2027 VDD VSS sg13g2_FILL8
XSTDFILL39_2035 VDD VSS sg13g2_FILL8
XSTDFILL39_2043 VDD VSS sg13g2_FILL8
XSTDFILL39_2051 VDD VSS sg13g2_FILL8
XSTDFILL39_2059 VDD VSS sg13g2_FILL8
XSTDFILL39_2067 VDD VSS sg13g2_FILL8
XSTDFILL39_2075 VDD VSS sg13g2_FILL8
XSTDFILL39_2083 VDD VSS sg13g2_FILL8
XSTDFILL39_2091 VDD VSS sg13g2_FILL8
XSTDFILL39_2099 VDD VSS sg13g2_FILL8
XSTDFILL39_2107 VDD VSS sg13g2_FILL8
XSTDFILL39_2115 VDD VSS sg13g2_FILL8
XSTDFILL39_2123 VDD VSS sg13g2_FILL8
XSTDFILL39_2131 VDD VSS sg13g2_FILL8
XSTDFILL39_2139 VDD VSS sg13g2_FILL8
XSTDFILL39_2147 VDD VSS sg13g2_FILL4
XSTDFILL39_2151 VDD VSS sg13g2_FILL2
XSTDFILL39_2153 VDD VSS sg13g2_FILL1
XSTDFILL40_0 VDD VSS sg13g2_FILL8
XSTDFILL40_8 VDD VSS sg13g2_FILL8
XSTDFILL40_16 VDD VSS sg13g2_FILL8
XSTDFILL40_24 VDD VSS sg13g2_FILL8
XSTDFILL40_32 VDD VSS sg13g2_FILL8
XSTDFILL40_40 VDD VSS sg13g2_FILL8
XSTDFILL40_48 VDD VSS sg13g2_FILL8
XSTDFILL40_56 VDD VSS sg13g2_FILL8
XSTDFILL40_64 VDD VSS sg13g2_FILL8
XSTDFILL40_72 VDD VSS sg13g2_FILL8
XSTDFILL40_80 VDD VSS sg13g2_FILL8
XSTDFILL40_88 VDD VSS sg13g2_FILL8
XSTDFILL40_96 VDD VSS sg13g2_FILL8
XSTDFILL40_104 VDD VSS sg13g2_FILL8
XSTDFILL40_112 VDD VSS sg13g2_FILL8
XSTDFILL40_120 VDD VSS sg13g2_FILL8
XSTDFILL40_128 VDD VSS sg13g2_FILL4
XSTDFILL40_1835 VDD VSS sg13g2_FILL8
XSTDFILL40_1843 VDD VSS sg13g2_FILL8
XSTDFILL40_1851 VDD VSS sg13g2_FILL8
XSTDFILL40_1859 VDD VSS sg13g2_FILL8
XSTDFILL40_1867 VDD VSS sg13g2_FILL8
XSTDFILL40_1875 VDD VSS sg13g2_FILL8
XSTDFILL40_1883 VDD VSS sg13g2_FILL8
XSTDFILL40_1891 VDD VSS sg13g2_FILL8
XSTDFILL40_1899 VDD VSS sg13g2_FILL8
XSTDFILL40_1907 VDD VSS sg13g2_FILL8
XSTDFILL40_1915 VDD VSS sg13g2_FILL8
XSTDFILL40_1923 VDD VSS sg13g2_FILL8
XSTDFILL40_1931 VDD VSS sg13g2_FILL8
XSTDFILL40_1939 VDD VSS sg13g2_FILL8
XSTDFILL40_1947 VDD VSS sg13g2_FILL8
XSTDFILL40_1955 VDD VSS sg13g2_FILL8
XSTDFILL40_1963 VDD VSS sg13g2_FILL8
XSTDFILL40_1971 VDD VSS sg13g2_FILL8
XSTDFILL40_1979 VDD VSS sg13g2_FILL8
XSTDFILL40_1987 VDD VSS sg13g2_FILL8
XSTDFILL40_1995 VDD VSS sg13g2_FILL8
XSTDFILL40_2003 VDD VSS sg13g2_FILL8
XSTDFILL40_2011 VDD VSS sg13g2_FILL8
XSTDFILL40_2019 VDD VSS sg13g2_FILL8
XSTDFILL40_2027 VDD VSS sg13g2_FILL8
XSTDFILL40_2035 VDD VSS sg13g2_FILL8
XSTDFILL40_2043 VDD VSS sg13g2_FILL8
XSTDFILL40_2051 VDD VSS sg13g2_FILL8
XSTDFILL40_2059 VDD VSS sg13g2_FILL8
XSTDFILL40_2067 VDD VSS sg13g2_FILL8
XSTDFILL40_2075 VDD VSS sg13g2_FILL8
XSTDFILL40_2083 VDD VSS sg13g2_FILL8
XSTDFILL40_2091 VDD VSS sg13g2_FILL8
XSTDFILL40_2099 VDD VSS sg13g2_FILL8
XSTDFILL40_2107 VDD VSS sg13g2_FILL8
XSTDFILL40_2115 VDD VSS sg13g2_FILL8
XSTDFILL40_2123 VDD VSS sg13g2_FILL8
XSTDFILL40_2131 VDD VSS sg13g2_FILL8
XSTDFILL40_2139 VDD VSS sg13g2_FILL8
XSTDFILL40_2147 VDD VSS sg13g2_FILL4
XSTDFILL40_2151 VDD VSS sg13g2_FILL2
XSTDFILL40_2153 VDD VSS sg13g2_FILL1
XSTDFILL41_0 VDD VSS sg13g2_FILL8
XSTDFILL41_8 VDD VSS sg13g2_FILL8
XSTDFILL41_16 VDD VSS sg13g2_FILL8
XSTDFILL41_24 VDD VSS sg13g2_FILL8
XSTDFILL41_32 VDD VSS sg13g2_FILL8
XSTDFILL41_40 VDD VSS sg13g2_FILL8
XSTDFILL41_48 VDD VSS sg13g2_FILL8
XSTDFILL41_56 VDD VSS sg13g2_FILL8
XSTDFILL41_64 VDD VSS sg13g2_FILL8
XSTDFILL41_72 VDD VSS sg13g2_FILL8
XSTDFILL41_80 VDD VSS sg13g2_FILL8
XSTDFILL41_88 VDD VSS sg13g2_FILL8
XSTDFILL41_96 VDD VSS sg13g2_FILL8
XSTDFILL41_104 VDD VSS sg13g2_FILL8
XSTDFILL41_112 VDD VSS sg13g2_FILL8
XSTDFILL41_120 VDD VSS sg13g2_FILL8
XSTDFILL41_128 VDD VSS sg13g2_FILL4
XSTDFILL41_1835 VDD VSS sg13g2_FILL8
XSTDFILL41_1843 VDD VSS sg13g2_FILL8
XSTDFILL41_1851 VDD VSS sg13g2_FILL8
XSTDFILL41_1859 VDD VSS sg13g2_FILL8
XSTDFILL41_1867 VDD VSS sg13g2_FILL8
XSTDFILL41_1875 VDD VSS sg13g2_FILL8
XSTDFILL41_1883 VDD VSS sg13g2_FILL8
XSTDFILL41_1891 VDD VSS sg13g2_FILL8
XSTDFILL41_1899 VDD VSS sg13g2_FILL8
XSTDFILL41_1907 VDD VSS sg13g2_FILL8
XSTDFILL41_1915 VDD VSS sg13g2_FILL8
XSTDFILL41_1923 VDD VSS sg13g2_FILL8
XSTDFILL41_1931 VDD VSS sg13g2_FILL8
XSTDFILL41_1939 VDD VSS sg13g2_FILL8
XSTDFILL41_1947 VDD VSS sg13g2_FILL8
XSTDFILL41_1955 VDD VSS sg13g2_FILL8
XSTDFILL41_1963 VDD VSS sg13g2_FILL8
XSTDFILL41_1971 VDD VSS sg13g2_FILL8
XSTDFILL41_1979 VDD VSS sg13g2_FILL8
XSTDFILL41_1987 VDD VSS sg13g2_FILL8
XSTDFILL41_1995 VDD VSS sg13g2_FILL8
XSTDFILL41_2003 VDD VSS sg13g2_FILL8
XSTDFILL41_2011 VDD VSS sg13g2_FILL8
XSTDFILL41_2019 VDD VSS sg13g2_FILL8
XSTDFILL41_2027 VDD VSS sg13g2_FILL8
XSTDFILL41_2035 VDD VSS sg13g2_FILL8
XSTDFILL41_2043 VDD VSS sg13g2_FILL8
XSTDFILL41_2051 VDD VSS sg13g2_FILL8
XSTDFILL41_2059 VDD VSS sg13g2_FILL8
XSTDFILL41_2067 VDD VSS sg13g2_FILL8
XSTDFILL41_2075 VDD VSS sg13g2_FILL8
XSTDFILL41_2083 VDD VSS sg13g2_FILL8
XSTDFILL41_2091 VDD VSS sg13g2_FILL8
XSTDFILL41_2099 VDD VSS sg13g2_FILL8
XSTDFILL41_2107 VDD VSS sg13g2_FILL8
XSTDFILL41_2115 VDD VSS sg13g2_FILL8
XSTDFILL41_2123 VDD VSS sg13g2_FILL8
XSTDFILL41_2131 VDD VSS sg13g2_FILL8
XSTDFILL41_2139 VDD VSS sg13g2_FILL8
XSTDFILL41_2147 VDD VSS sg13g2_FILL4
XSTDFILL41_2151 VDD VSS sg13g2_FILL2
XSTDFILL41_2153 VDD VSS sg13g2_FILL1
XSTDFILL42_0 VDD VSS sg13g2_FILL8
XSTDFILL42_8 VDD VSS sg13g2_FILL8
XSTDFILL42_16 VDD VSS sg13g2_FILL8
XSTDFILL42_24 VDD VSS sg13g2_FILL8
XSTDFILL42_32 VDD VSS sg13g2_FILL8
XSTDFILL42_40 VDD VSS sg13g2_FILL8
XSTDFILL42_48 VDD VSS sg13g2_FILL8
XSTDFILL42_56 VDD VSS sg13g2_FILL8
XSTDFILL42_64 VDD VSS sg13g2_FILL8
XSTDFILL42_72 VDD VSS sg13g2_FILL8
XSTDFILL42_80 VDD VSS sg13g2_FILL8
XSTDFILL42_88 VDD VSS sg13g2_FILL8
XSTDFILL42_96 VDD VSS sg13g2_FILL8
XSTDFILL42_104 VDD VSS sg13g2_FILL8
XSTDFILL42_112 VDD VSS sg13g2_FILL8
XSTDFILL42_120 VDD VSS sg13g2_FILL8
XSTDFILL42_128 VDD VSS sg13g2_FILL4
XSTDFILL42_1835 VDD VSS sg13g2_FILL8
XSTDFILL42_1843 VDD VSS sg13g2_FILL8
XSTDFILL42_1851 VDD VSS sg13g2_FILL8
XSTDFILL42_1859 VDD VSS sg13g2_FILL8
XSTDFILL42_1867 VDD VSS sg13g2_FILL8
XSTDFILL42_1875 VDD VSS sg13g2_FILL8
XSTDFILL42_1883 VDD VSS sg13g2_FILL8
XSTDFILL42_1891 VDD VSS sg13g2_FILL8
XSTDFILL42_1899 VDD VSS sg13g2_FILL8
XSTDFILL42_1907 VDD VSS sg13g2_FILL8
XSTDFILL42_1915 VDD VSS sg13g2_FILL8
XSTDFILL42_1923 VDD VSS sg13g2_FILL8
XSTDFILL42_1931 VDD VSS sg13g2_FILL8
XSTDFILL42_1939 VDD VSS sg13g2_FILL8
XSTDFILL42_1947 VDD VSS sg13g2_FILL8
XSTDFILL42_1955 VDD VSS sg13g2_FILL8
XSTDFILL42_1963 VDD VSS sg13g2_FILL8
XSTDFILL42_1971 VDD VSS sg13g2_FILL8
XSTDFILL42_1979 VDD VSS sg13g2_FILL8
XSTDFILL42_1987 VDD VSS sg13g2_FILL8
XSTDFILL42_1995 VDD VSS sg13g2_FILL8
XSTDFILL42_2003 VDD VSS sg13g2_FILL8
XSTDFILL42_2011 VDD VSS sg13g2_FILL8
XSTDFILL42_2019 VDD VSS sg13g2_FILL8
XSTDFILL42_2027 VDD VSS sg13g2_FILL8
XSTDFILL42_2035 VDD VSS sg13g2_FILL8
XSTDFILL42_2043 VDD VSS sg13g2_FILL8
XSTDFILL42_2051 VDD VSS sg13g2_FILL8
XSTDFILL42_2059 VDD VSS sg13g2_FILL8
XSTDFILL42_2067 VDD VSS sg13g2_FILL8
XSTDFILL42_2075 VDD VSS sg13g2_FILL8
XSTDFILL42_2083 VDD VSS sg13g2_FILL8
XSTDFILL42_2091 VDD VSS sg13g2_FILL8
XSTDFILL42_2099 VDD VSS sg13g2_FILL8
XSTDFILL42_2107 VDD VSS sg13g2_FILL8
XSTDFILL42_2115 VDD VSS sg13g2_FILL8
XSTDFILL42_2123 VDD VSS sg13g2_FILL8
XSTDFILL42_2131 VDD VSS sg13g2_FILL8
XSTDFILL42_2139 VDD VSS sg13g2_FILL8
XSTDFILL42_2147 VDD VSS sg13g2_FILL4
XSTDFILL42_2151 VDD VSS sg13g2_FILL2
XSTDFILL42_2153 VDD VSS sg13g2_FILL1
XSTDFILL43_0 VDD VSS sg13g2_FILL8
XSTDFILL43_8 VDD VSS sg13g2_FILL8
XSTDFILL43_16 VDD VSS sg13g2_FILL8
XSTDFILL43_24 VDD VSS sg13g2_FILL8
XSTDFILL43_32 VDD VSS sg13g2_FILL8
XSTDFILL43_40 VDD VSS sg13g2_FILL8
XSTDFILL43_48 VDD VSS sg13g2_FILL8
XSTDFILL43_56 VDD VSS sg13g2_FILL8
XSTDFILL43_64 VDD VSS sg13g2_FILL8
XSTDFILL43_72 VDD VSS sg13g2_FILL8
XSTDFILL43_80 VDD VSS sg13g2_FILL8
XSTDFILL43_88 VDD VSS sg13g2_FILL8
XSTDFILL43_96 VDD VSS sg13g2_FILL8
XSTDFILL43_104 VDD VSS sg13g2_FILL8
XSTDFILL43_112 VDD VSS sg13g2_FILL8
XSTDFILL43_120 VDD VSS sg13g2_FILL8
XSTDFILL43_128 VDD VSS sg13g2_FILL4
XSTDFILL43_1835 VDD VSS sg13g2_FILL8
XSTDFILL43_1843 VDD VSS sg13g2_FILL8
XSTDFILL43_1851 VDD VSS sg13g2_FILL8
XSTDFILL43_1859 VDD VSS sg13g2_FILL8
XSTDFILL43_1867 VDD VSS sg13g2_FILL8
XSTDFILL43_1875 VDD VSS sg13g2_FILL8
XSTDFILL43_1883 VDD VSS sg13g2_FILL8
XSTDFILL43_1891 VDD VSS sg13g2_FILL8
XSTDFILL43_1899 VDD VSS sg13g2_FILL8
XSTDFILL43_1907 VDD VSS sg13g2_FILL8
XSTDFILL43_1915 VDD VSS sg13g2_FILL8
XSTDFILL43_1923 VDD VSS sg13g2_FILL8
XSTDFILL43_1931 VDD VSS sg13g2_FILL8
XSTDFILL43_1939 VDD VSS sg13g2_FILL8
XSTDFILL43_1947 VDD VSS sg13g2_FILL8
XSTDFILL43_1955 VDD VSS sg13g2_FILL8
XSTDFILL43_1963 VDD VSS sg13g2_FILL8
XSTDFILL43_1971 VDD VSS sg13g2_FILL8
XSTDFILL43_1979 VDD VSS sg13g2_FILL8
XSTDFILL43_1987 VDD VSS sg13g2_FILL8
XSTDFILL43_1995 VDD VSS sg13g2_FILL8
XSTDFILL43_2003 VDD VSS sg13g2_FILL8
XSTDFILL43_2011 VDD VSS sg13g2_FILL8
XSTDFILL43_2019 VDD VSS sg13g2_FILL8
XSTDFILL43_2027 VDD VSS sg13g2_FILL8
XSTDFILL43_2035 VDD VSS sg13g2_FILL8
XSTDFILL43_2043 VDD VSS sg13g2_FILL8
XSTDFILL43_2051 VDD VSS sg13g2_FILL8
XSTDFILL43_2059 VDD VSS sg13g2_FILL8
XSTDFILL43_2067 VDD VSS sg13g2_FILL8
XSTDFILL43_2075 VDD VSS sg13g2_FILL8
XSTDFILL43_2083 VDD VSS sg13g2_FILL8
XSTDFILL43_2091 VDD VSS sg13g2_FILL8
XSTDFILL43_2099 VDD VSS sg13g2_FILL8
XSTDFILL43_2107 VDD VSS sg13g2_FILL8
XSTDFILL43_2115 VDD VSS sg13g2_FILL8
XSTDFILL43_2123 VDD VSS sg13g2_FILL8
XSTDFILL43_2131 VDD VSS sg13g2_FILL8
XSTDFILL43_2139 VDD VSS sg13g2_FILL8
XSTDFILL43_2147 VDD VSS sg13g2_FILL4
XSTDFILL43_2151 VDD VSS sg13g2_FILL2
XSTDFILL43_2153 VDD VSS sg13g2_FILL1
XSTDFILL44_0 VDD VSS sg13g2_FILL8
XSTDFILL44_8 VDD VSS sg13g2_FILL8
XSTDFILL44_16 VDD VSS sg13g2_FILL8
XSTDFILL44_24 VDD VSS sg13g2_FILL8
XSTDFILL44_32 VDD VSS sg13g2_FILL8
XSTDFILL44_40 VDD VSS sg13g2_FILL8
XSTDFILL44_48 VDD VSS sg13g2_FILL8
XSTDFILL44_56 VDD VSS sg13g2_FILL8
XSTDFILL44_64 VDD VSS sg13g2_FILL8
XSTDFILL44_72 VDD VSS sg13g2_FILL8
XSTDFILL44_80 VDD VSS sg13g2_FILL8
XSTDFILL44_88 VDD VSS sg13g2_FILL8
XSTDFILL44_96 VDD VSS sg13g2_FILL8
XSTDFILL44_104 VDD VSS sg13g2_FILL8
XSTDFILL44_112 VDD VSS sg13g2_FILL8
XSTDFILL44_120 VDD VSS sg13g2_FILL8
XSTDFILL44_128 VDD VSS sg13g2_FILL4
XSTDFILL44_1835 VDD VSS sg13g2_FILL8
XSTDFILL44_1843 VDD VSS sg13g2_FILL8
XSTDFILL44_1851 VDD VSS sg13g2_FILL8
XSTDFILL44_1859 VDD VSS sg13g2_FILL8
XSTDFILL44_1867 VDD VSS sg13g2_FILL8
XSTDFILL44_1875 VDD VSS sg13g2_FILL8
XSTDFILL44_1883 VDD VSS sg13g2_FILL8
XSTDFILL44_1891 VDD VSS sg13g2_FILL8
XSTDFILL44_1899 VDD VSS sg13g2_FILL8
XSTDFILL44_1907 VDD VSS sg13g2_FILL8
XSTDFILL44_1915 VDD VSS sg13g2_FILL8
XSTDFILL44_1923 VDD VSS sg13g2_FILL8
XSTDFILL44_1931 VDD VSS sg13g2_FILL8
XSTDFILL44_1939 VDD VSS sg13g2_FILL8
XSTDFILL44_1947 VDD VSS sg13g2_FILL8
XSTDFILL44_1955 VDD VSS sg13g2_FILL8
XSTDFILL44_1963 VDD VSS sg13g2_FILL8
XSTDFILL44_1971 VDD VSS sg13g2_FILL8
XSTDFILL44_1979 VDD VSS sg13g2_FILL8
XSTDFILL44_1987 VDD VSS sg13g2_FILL8
XSTDFILL44_1995 VDD VSS sg13g2_FILL8
XSTDFILL44_2003 VDD VSS sg13g2_FILL8
XSTDFILL44_2011 VDD VSS sg13g2_FILL8
XSTDFILL44_2019 VDD VSS sg13g2_FILL8
XSTDFILL44_2027 VDD VSS sg13g2_FILL8
XSTDFILL44_2035 VDD VSS sg13g2_FILL8
XSTDFILL44_2043 VDD VSS sg13g2_FILL8
XSTDFILL44_2051 VDD VSS sg13g2_FILL8
XSTDFILL44_2059 VDD VSS sg13g2_FILL8
XSTDFILL44_2067 VDD VSS sg13g2_FILL8
XSTDFILL44_2075 VDD VSS sg13g2_FILL8
XSTDFILL44_2083 VDD VSS sg13g2_FILL8
XSTDFILL44_2091 VDD VSS sg13g2_FILL8
XSTDFILL44_2099 VDD VSS sg13g2_FILL8
XSTDFILL44_2107 VDD VSS sg13g2_FILL8
XSTDFILL44_2115 VDD VSS sg13g2_FILL8
XSTDFILL44_2123 VDD VSS sg13g2_FILL8
XSTDFILL44_2131 VDD VSS sg13g2_FILL8
XSTDFILL44_2139 VDD VSS sg13g2_FILL8
XSTDFILL44_2147 VDD VSS sg13g2_FILL4
XSTDFILL44_2151 VDD VSS sg13g2_FILL2
XSTDFILL44_2153 VDD VSS sg13g2_FILL1
XSTDFILL45_0 VDD VSS sg13g2_FILL8
XSTDFILL45_8 VDD VSS sg13g2_FILL8
XSTDFILL45_16 VDD VSS sg13g2_FILL8
XSTDFILL45_24 VDD VSS sg13g2_FILL8
XSTDFILL45_32 VDD VSS sg13g2_FILL8
XSTDFILL45_40 VDD VSS sg13g2_FILL8
XSTDFILL45_48 VDD VSS sg13g2_FILL8
XSTDFILL45_56 VDD VSS sg13g2_FILL8
XSTDFILL45_64 VDD VSS sg13g2_FILL8
XSTDFILL45_72 VDD VSS sg13g2_FILL8
XSTDFILL45_80 VDD VSS sg13g2_FILL8
XSTDFILL45_88 VDD VSS sg13g2_FILL8
XSTDFILL45_96 VDD VSS sg13g2_FILL8
XSTDFILL45_104 VDD VSS sg13g2_FILL8
XSTDFILL45_112 VDD VSS sg13g2_FILL8
XSTDFILL45_120 VDD VSS sg13g2_FILL8
XSTDFILL45_128 VDD VSS sg13g2_FILL4
XSTDFILL45_1835 VDD VSS sg13g2_FILL8
XSTDFILL45_1843 VDD VSS sg13g2_FILL8
XSTDFILL45_1851 VDD VSS sg13g2_FILL8
XSTDFILL45_1859 VDD VSS sg13g2_FILL8
XSTDFILL45_1867 VDD VSS sg13g2_FILL8
XSTDFILL45_1875 VDD VSS sg13g2_FILL8
XSTDFILL45_1883 VDD VSS sg13g2_FILL8
XSTDFILL45_1891 VDD VSS sg13g2_FILL8
XSTDFILL45_1899 VDD VSS sg13g2_FILL8
XSTDFILL45_1907 VDD VSS sg13g2_FILL8
XSTDFILL45_1915 VDD VSS sg13g2_FILL8
XSTDFILL45_1923 VDD VSS sg13g2_FILL8
XSTDFILL45_1931 VDD VSS sg13g2_FILL8
XSTDFILL45_1939 VDD VSS sg13g2_FILL8
XSTDFILL45_1947 VDD VSS sg13g2_FILL8
XSTDFILL45_1955 VDD VSS sg13g2_FILL8
XSTDFILL45_1963 VDD VSS sg13g2_FILL8
XSTDFILL45_1971 VDD VSS sg13g2_FILL8
XSTDFILL45_1979 VDD VSS sg13g2_FILL8
XSTDFILL45_1987 VDD VSS sg13g2_FILL8
XSTDFILL45_1995 VDD VSS sg13g2_FILL8
XSTDFILL45_2003 VDD VSS sg13g2_FILL8
XSTDFILL45_2011 VDD VSS sg13g2_FILL8
XSTDFILL45_2019 VDD VSS sg13g2_FILL8
XSTDFILL45_2027 VDD VSS sg13g2_FILL8
XSTDFILL45_2035 VDD VSS sg13g2_FILL8
XSTDFILL45_2043 VDD VSS sg13g2_FILL8
XSTDFILL45_2051 VDD VSS sg13g2_FILL8
XSTDFILL45_2059 VDD VSS sg13g2_FILL8
XSTDFILL45_2067 VDD VSS sg13g2_FILL8
XSTDFILL45_2075 VDD VSS sg13g2_FILL8
XSTDFILL45_2083 VDD VSS sg13g2_FILL8
XSTDFILL45_2091 VDD VSS sg13g2_FILL8
XSTDFILL45_2099 VDD VSS sg13g2_FILL8
XSTDFILL45_2107 VDD VSS sg13g2_FILL8
XSTDFILL45_2115 VDD VSS sg13g2_FILL8
XSTDFILL45_2123 VDD VSS sg13g2_FILL8
XSTDFILL45_2131 VDD VSS sg13g2_FILL8
XSTDFILL45_2139 VDD VSS sg13g2_FILL8
XSTDFILL45_2147 VDD VSS sg13g2_FILL4
XSTDFILL45_2151 VDD VSS sg13g2_FILL2
XSTDFILL45_2153 VDD VSS sg13g2_FILL1
XSTDFILL46_0 VDD VSS sg13g2_FILL8
XSTDFILL46_8 VDD VSS sg13g2_FILL8
XSTDFILL46_16 VDD VSS sg13g2_FILL8
XSTDFILL46_24 VDD VSS sg13g2_FILL8
XSTDFILL46_32 VDD VSS sg13g2_FILL8
XSTDFILL46_40 VDD VSS sg13g2_FILL8
XSTDFILL46_48 VDD VSS sg13g2_FILL8
XSTDFILL46_56 VDD VSS sg13g2_FILL8
XSTDFILL46_64 VDD VSS sg13g2_FILL8
XSTDFILL46_72 VDD VSS sg13g2_FILL8
XSTDFILL46_80 VDD VSS sg13g2_FILL8
XSTDFILL46_88 VDD VSS sg13g2_FILL8
XSTDFILL46_96 VDD VSS sg13g2_FILL8
XSTDFILL46_104 VDD VSS sg13g2_FILL8
XSTDFILL46_112 VDD VSS sg13g2_FILL8
XSTDFILL46_120 VDD VSS sg13g2_FILL8
XSTDFILL46_128 VDD VSS sg13g2_FILL4
XSTDFILL46_1835 VDD VSS sg13g2_FILL8
XSTDFILL46_1843 VDD VSS sg13g2_FILL8
XSTDFILL46_1851 VDD VSS sg13g2_FILL8
XSTDFILL46_1859 VDD VSS sg13g2_FILL8
XSTDFILL46_1867 VDD VSS sg13g2_FILL8
XSTDFILL46_1875 VDD VSS sg13g2_FILL8
XSTDFILL46_1883 VDD VSS sg13g2_FILL8
XSTDFILL46_1891 VDD VSS sg13g2_FILL8
XSTDFILL46_1899 VDD VSS sg13g2_FILL8
XSTDFILL46_1907 VDD VSS sg13g2_FILL8
XSTDFILL46_1915 VDD VSS sg13g2_FILL8
XSTDFILL46_1923 VDD VSS sg13g2_FILL8
XSTDFILL46_1931 VDD VSS sg13g2_FILL8
XSTDFILL46_1939 VDD VSS sg13g2_FILL8
XSTDFILL46_1947 VDD VSS sg13g2_FILL8
XSTDFILL46_1955 VDD VSS sg13g2_FILL8
XSTDFILL46_1963 VDD VSS sg13g2_FILL8
XSTDFILL46_1971 VDD VSS sg13g2_FILL8
XSTDFILL46_1979 VDD VSS sg13g2_FILL8
XSTDFILL46_1987 VDD VSS sg13g2_FILL8
XSTDFILL46_1995 VDD VSS sg13g2_FILL8
XSTDFILL46_2003 VDD VSS sg13g2_FILL8
XSTDFILL46_2011 VDD VSS sg13g2_FILL8
XSTDFILL46_2019 VDD VSS sg13g2_FILL8
XSTDFILL46_2027 VDD VSS sg13g2_FILL8
XSTDFILL46_2035 VDD VSS sg13g2_FILL8
XSTDFILL46_2043 VDD VSS sg13g2_FILL8
XSTDFILL46_2051 VDD VSS sg13g2_FILL8
XSTDFILL46_2059 VDD VSS sg13g2_FILL8
XSTDFILL46_2067 VDD VSS sg13g2_FILL8
XSTDFILL46_2075 VDD VSS sg13g2_FILL8
XSTDFILL46_2083 VDD VSS sg13g2_FILL8
XSTDFILL46_2091 VDD VSS sg13g2_FILL8
XSTDFILL46_2099 VDD VSS sg13g2_FILL8
XSTDFILL46_2107 VDD VSS sg13g2_FILL8
XSTDFILL46_2115 VDD VSS sg13g2_FILL8
XSTDFILL46_2123 VDD VSS sg13g2_FILL8
XSTDFILL46_2131 VDD VSS sg13g2_FILL8
XSTDFILL46_2139 VDD VSS sg13g2_FILL8
XSTDFILL46_2147 VDD VSS sg13g2_FILL4
XSTDFILL46_2151 VDD VSS sg13g2_FILL2
XSTDFILL46_2153 VDD VSS sg13g2_FILL1
XSTDFILL47_0 VDD VSS sg13g2_FILL8
XSTDFILL47_8 VDD VSS sg13g2_FILL8
XSTDFILL47_16 VDD VSS sg13g2_FILL8
XSTDFILL47_24 VDD VSS sg13g2_FILL8
XSTDFILL47_32 VDD VSS sg13g2_FILL8
XSTDFILL47_40 VDD VSS sg13g2_FILL8
XSTDFILL47_48 VDD VSS sg13g2_FILL8
XSTDFILL47_56 VDD VSS sg13g2_FILL8
XSTDFILL47_64 VDD VSS sg13g2_FILL8
XSTDFILL47_72 VDD VSS sg13g2_FILL8
XSTDFILL47_80 VDD VSS sg13g2_FILL8
XSTDFILL47_88 VDD VSS sg13g2_FILL8
XSTDFILL47_96 VDD VSS sg13g2_FILL8
XSTDFILL47_104 VDD VSS sg13g2_FILL8
XSTDFILL47_112 VDD VSS sg13g2_FILL8
XSTDFILL47_120 VDD VSS sg13g2_FILL8
XSTDFILL47_128 VDD VSS sg13g2_FILL4
XSTDFILL47_1835 VDD VSS sg13g2_FILL8
XSTDFILL47_1843 VDD VSS sg13g2_FILL8
XSTDFILL47_1851 VDD VSS sg13g2_FILL8
XSTDFILL47_1859 VDD VSS sg13g2_FILL8
XSTDFILL47_1867 VDD VSS sg13g2_FILL8
XSTDFILL47_1875 VDD VSS sg13g2_FILL8
XSTDFILL47_1883 VDD VSS sg13g2_FILL8
XSTDFILL47_1891 VDD VSS sg13g2_FILL8
XSTDFILL47_1899 VDD VSS sg13g2_FILL8
XSTDFILL47_1907 VDD VSS sg13g2_FILL8
XSTDFILL47_1915 VDD VSS sg13g2_FILL8
XSTDFILL47_1923 VDD VSS sg13g2_FILL8
XSTDFILL47_1931 VDD VSS sg13g2_FILL8
XSTDFILL47_1939 VDD VSS sg13g2_FILL8
XSTDFILL47_1947 VDD VSS sg13g2_FILL8
XSTDFILL47_1955 VDD VSS sg13g2_FILL8
XSTDFILL47_1963 VDD VSS sg13g2_FILL8
XSTDFILL47_1971 VDD VSS sg13g2_FILL8
XSTDFILL47_1979 VDD VSS sg13g2_FILL8
XSTDFILL47_1987 VDD VSS sg13g2_FILL8
XSTDFILL47_1995 VDD VSS sg13g2_FILL8
XSTDFILL47_2003 VDD VSS sg13g2_FILL8
XSTDFILL47_2011 VDD VSS sg13g2_FILL8
XSTDFILL47_2019 VDD VSS sg13g2_FILL8
XSTDFILL47_2027 VDD VSS sg13g2_FILL8
XSTDFILL47_2035 VDD VSS sg13g2_FILL8
XSTDFILL47_2043 VDD VSS sg13g2_FILL8
XSTDFILL47_2051 VDD VSS sg13g2_FILL8
XSTDFILL47_2059 VDD VSS sg13g2_FILL8
XSTDFILL47_2067 VDD VSS sg13g2_FILL8
XSTDFILL47_2075 VDD VSS sg13g2_FILL8
XSTDFILL47_2083 VDD VSS sg13g2_FILL8
XSTDFILL47_2091 VDD VSS sg13g2_FILL8
XSTDFILL47_2099 VDD VSS sg13g2_FILL8
XSTDFILL47_2107 VDD VSS sg13g2_FILL8
XSTDFILL47_2115 VDD VSS sg13g2_FILL8
XSTDFILL47_2123 VDD VSS sg13g2_FILL8
XSTDFILL47_2131 VDD VSS sg13g2_FILL8
XSTDFILL47_2139 VDD VSS sg13g2_FILL8
XSTDFILL47_2147 VDD VSS sg13g2_FILL4
XSTDFILL47_2151 VDD VSS sg13g2_FILL2
XSTDFILL47_2153 VDD VSS sg13g2_FILL1
XSTDFILL48_0 VDD VSS sg13g2_FILL8
XSTDFILL48_8 VDD VSS sg13g2_FILL8
XSTDFILL48_16 VDD VSS sg13g2_FILL8
XSTDFILL48_24 VDD VSS sg13g2_FILL8
XSTDFILL48_32 VDD VSS sg13g2_FILL8
XSTDFILL48_40 VDD VSS sg13g2_FILL8
XSTDFILL48_48 VDD VSS sg13g2_FILL8
XSTDFILL48_56 VDD VSS sg13g2_FILL8
XSTDFILL48_64 VDD VSS sg13g2_FILL8
XSTDFILL48_72 VDD VSS sg13g2_FILL8
XSTDFILL48_80 VDD VSS sg13g2_FILL8
XSTDFILL48_88 VDD VSS sg13g2_FILL8
XSTDFILL48_96 VDD VSS sg13g2_FILL8
XSTDFILL48_104 VDD VSS sg13g2_FILL8
XSTDFILL48_112 VDD VSS sg13g2_FILL8
XSTDFILL48_120 VDD VSS sg13g2_FILL8
XSTDFILL48_128 VDD VSS sg13g2_FILL4
XSTDFILL48_1835 VDD VSS sg13g2_FILL8
XSTDFILL48_1843 VDD VSS sg13g2_FILL8
XSTDFILL48_1851 VDD VSS sg13g2_FILL8
XSTDFILL48_1859 VDD VSS sg13g2_FILL8
XSTDFILL48_1867 VDD VSS sg13g2_FILL8
XSTDFILL48_1875 VDD VSS sg13g2_FILL8
XSTDFILL48_1883 VDD VSS sg13g2_FILL8
XSTDFILL48_1891 VDD VSS sg13g2_FILL8
XSTDFILL48_1899 VDD VSS sg13g2_FILL8
XSTDFILL48_1907 VDD VSS sg13g2_FILL8
XSTDFILL48_1915 VDD VSS sg13g2_FILL8
XSTDFILL48_1923 VDD VSS sg13g2_FILL8
XSTDFILL48_1931 VDD VSS sg13g2_FILL8
XSTDFILL48_1939 VDD VSS sg13g2_FILL8
XSTDFILL48_1947 VDD VSS sg13g2_FILL8
XSTDFILL48_1955 VDD VSS sg13g2_FILL8
XSTDFILL48_1963 VDD VSS sg13g2_FILL8
XSTDFILL48_1971 VDD VSS sg13g2_FILL8
XSTDFILL48_1979 VDD VSS sg13g2_FILL8
XSTDFILL48_1987 VDD VSS sg13g2_FILL8
XSTDFILL48_1995 VDD VSS sg13g2_FILL8
XSTDFILL48_2003 VDD VSS sg13g2_FILL8
XSTDFILL48_2011 VDD VSS sg13g2_FILL8
XSTDFILL48_2019 VDD VSS sg13g2_FILL8
XSTDFILL48_2027 VDD VSS sg13g2_FILL8
XSTDFILL48_2035 VDD VSS sg13g2_FILL8
XSTDFILL48_2043 VDD VSS sg13g2_FILL8
XSTDFILL48_2051 VDD VSS sg13g2_FILL8
XSTDFILL48_2059 VDD VSS sg13g2_FILL8
XSTDFILL48_2067 VDD VSS sg13g2_FILL8
XSTDFILL48_2075 VDD VSS sg13g2_FILL8
XSTDFILL48_2083 VDD VSS sg13g2_FILL8
XSTDFILL48_2091 VDD VSS sg13g2_FILL8
XSTDFILL48_2099 VDD VSS sg13g2_FILL8
XSTDFILL48_2107 VDD VSS sg13g2_FILL8
XSTDFILL48_2115 VDD VSS sg13g2_FILL8
XSTDFILL48_2123 VDD VSS sg13g2_FILL8
XSTDFILL48_2131 VDD VSS sg13g2_FILL8
XSTDFILL48_2139 VDD VSS sg13g2_FILL8
XSTDFILL48_2147 VDD VSS sg13g2_FILL4
XSTDFILL48_2151 VDD VSS sg13g2_FILL2
XSTDFILL48_2153 VDD VSS sg13g2_FILL1
XSTDFILL49_0 VDD VSS sg13g2_FILL8
XSTDFILL49_8 VDD VSS sg13g2_FILL8
XSTDFILL49_16 VDD VSS sg13g2_FILL8
XSTDFILL49_24 VDD VSS sg13g2_FILL8
XSTDFILL49_32 VDD VSS sg13g2_FILL8
XSTDFILL49_40 VDD VSS sg13g2_FILL8
XSTDFILL49_48 VDD VSS sg13g2_FILL8
XSTDFILL49_56 VDD VSS sg13g2_FILL8
XSTDFILL49_64 VDD VSS sg13g2_FILL8
XSTDFILL49_72 VDD VSS sg13g2_FILL8
XSTDFILL49_80 VDD VSS sg13g2_FILL8
XSTDFILL49_88 VDD VSS sg13g2_FILL8
XSTDFILL49_96 VDD VSS sg13g2_FILL8
XSTDFILL49_104 VDD VSS sg13g2_FILL8
XSTDFILL49_112 VDD VSS sg13g2_FILL8
XSTDFILL49_120 VDD VSS sg13g2_FILL8
XSTDFILL49_128 VDD VSS sg13g2_FILL4
XSTDFILL49_1835 VDD VSS sg13g2_FILL8
XSTDFILL49_1843 VDD VSS sg13g2_FILL8
XSTDFILL49_1851 VDD VSS sg13g2_FILL8
XSTDFILL49_1859 VDD VSS sg13g2_FILL8
XSTDFILL49_1867 VDD VSS sg13g2_FILL8
XSTDFILL49_1875 VDD VSS sg13g2_FILL8
XSTDFILL49_1883 VDD VSS sg13g2_FILL8
XSTDFILL49_1891 VDD VSS sg13g2_FILL8
XSTDFILL49_1899 VDD VSS sg13g2_FILL8
XSTDFILL49_1907 VDD VSS sg13g2_FILL8
XSTDFILL49_1915 VDD VSS sg13g2_FILL8
XSTDFILL49_1923 VDD VSS sg13g2_FILL8
XSTDFILL49_1931 VDD VSS sg13g2_FILL8
XSTDFILL49_1939 VDD VSS sg13g2_FILL8
XSTDFILL49_1947 VDD VSS sg13g2_FILL8
XSTDFILL49_1955 VDD VSS sg13g2_FILL8
XSTDFILL49_1963 VDD VSS sg13g2_FILL8
XSTDFILL49_1971 VDD VSS sg13g2_FILL8
XSTDFILL49_1979 VDD VSS sg13g2_FILL8
XSTDFILL49_1987 VDD VSS sg13g2_FILL8
XSTDFILL49_1995 VDD VSS sg13g2_FILL8
XSTDFILL49_2003 VDD VSS sg13g2_FILL8
XSTDFILL49_2011 VDD VSS sg13g2_FILL8
XSTDFILL49_2019 VDD VSS sg13g2_FILL8
XSTDFILL49_2027 VDD VSS sg13g2_FILL8
XSTDFILL49_2035 VDD VSS sg13g2_FILL8
XSTDFILL49_2043 VDD VSS sg13g2_FILL8
XSTDFILL49_2051 VDD VSS sg13g2_FILL8
XSTDFILL49_2059 VDD VSS sg13g2_FILL8
XSTDFILL49_2067 VDD VSS sg13g2_FILL8
XSTDFILL49_2075 VDD VSS sg13g2_FILL8
XSTDFILL49_2083 VDD VSS sg13g2_FILL8
XSTDFILL49_2091 VDD VSS sg13g2_FILL8
XSTDFILL49_2099 VDD VSS sg13g2_FILL8
XSTDFILL49_2107 VDD VSS sg13g2_FILL8
XSTDFILL49_2115 VDD VSS sg13g2_FILL8
XSTDFILL49_2123 VDD VSS sg13g2_FILL8
XSTDFILL49_2131 VDD VSS sg13g2_FILL8
XSTDFILL49_2139 VDD VSS sg13g2_FILL8
XSTDFILL49_2147 VDD VSS sg13g2_FILL4
XSTDFILL49_2151 VDD VSS sg13g2_FILL2
XSTDFILL49_2153 VDD VSS sg13g2_FILL1
XSTDFILL50_0 VDD VSS sg13g2_FILL8
XSTDFILL50_8 VDD VSS sg13g2_FILL8
XSTDFILL50_16 VDD VSS sg13g2_FILL8
XSTDFILL50_24 VDD VSS sg13g2_FILL8
XSTDFILL50_32 VDD VSS sg13g2_FILL8
XSTDFILL50_40 VDD VSS sg13g2_FILL8
XSTDFILL50_48 VDD VSS sg13g2_FILL8
XSTDFILL50_56 VDD VSS sg13g2_FILL8
XSTDFILL50_64 VDD VSS sg13g2_FILL8
XSTDFILL50_72 VDD VSS sg13g2_FILL8
XSTDFILL50_80 VDD VSS sg13g2_FILL8
XSTDFILL50_88 VDD VSS sg13g2_FILL8
XSTDFILL50_96 VDD VSS sg13g2_FILL8
XSTDFILL50_104 VDD VSS sg13g2_FILL8
XSTDFILL50_112 VDD VSS sg13g2_FILL8
XSTDFILL50_120 VDD VSS sg13g2_FILL8
XSTDFILL50_128 VDD VSS sg13g2_FILL4
XSTDFILL50_1835 VDD VSS sg13g2_FILL8
XSTDFILL50_1843 VDD VSS sg13g2_FILL8
XSTDFILL50_1851 VDD VSS sg13g2_FILL8
XSTDFILL50_1859 VDD VSS sg13g2_FILL8
XSTDFILL50_1867 VDD VSS sg13g2_FILL8
XSTDFILL50_1875 VDD VSS sg13g2_FILL8
XSTDFILL50_1883 VDD VSS sg13g2_FILL8
XSTDFILL50_1891 VDD VSS sg13g2_FILL8
XSTDFILL50_1899 VDD VSS sg13g2_FILL8
XSTDFILL50_1907 VDD VSS sg13g2_FILL8
XSTDFILL50_1915 VDD VSS sg13g2_FILL8
XSTDFILL50_1923 VDD VSS sg13g2_FILL8
XSTDFILL50_1931 VDD VSS sg13g2_FILL8
XSTDFILL50_1939 VDD VSS sg13g2_FILL8
XSTDFILL50_1947 VDD VSS sg13g2_FILL8
XSTDFILL50_1955 VDD VSS sg13g2_FILL8
XSTDFILL50_1963 VDD VSS sg13g2_FILL8
XSTDFILL50_1971 VDD VSS sg13g2_FILL8
XSTDFILL50_1979 VDD VSS sg13g2_FILL8
XSTDFILL50_1987 VDD VSS sg13g2_FILL8
XSTDFILL50_1995 VDD VSS sg13g2_FILL8
XSTDFILL50_2003 VDD VSS sg13g2_FILL8
XSTDFILL50_2011 VDD VSS sg13g2_FILL8
XSTDFILL50_2019 VDD VSS sg13g2_FILL8
XSTDFILL50_2027 VDD VSS sg13g2_FILL8
XSTDFILL50_2035 VDD VSS sg13g2_FILL8
XSTDFILL50_2043 VDD VSS sg13g2_FILL8
XSTDFILL50_2051 VDD VSS sg13g2_FILL8
XSTDFILL50_2059 VDD VSS sg13g2_FILL8
XSTDFILL50_2067 VDD VSS sg13g2_FILL8
XSTDFILL50_2075 VDD VSS sg13g2_FILL8
XSTDFILL50_2083 VDD VSS sg13g2_FILL8
XSTDFILL50_2091 VDD VSS sg13g2_FILL8
XSTDFILL50_2099 VDD VSS sg13g2_FILL8
XSTDFILL50_2107 VDD VSS sg13g2_FILL8
XSTDFILL50_2115 VDD VSS sg13g2_FILL8
XSTDFILL50_2123 VDD VSS sg13g2_FILL8
XSTDFILL50_2131 VDD VSS sg13g2_FILL8
XSTDFILL50_2139 VDD VSS sg13g2_FILL8
XSTDFILL50_2147 VDD VSS sg13g2_FILL4
XSTDFILL50_2151 VDD VSS sg13g2_FILL2
XSTDFILL50_2153 VDD VSS sg13g2_FILL1
XSTDFILL51_0 VDD VSS sg13g2_FILL8
XSTDFILL51_8 VDD VSS sg13g2_FILL8
XSTDFILL51_16 VDD VSS sg13g2_FILL8
XSTDFILL51_24 VDD VSS sg13g2_FILL8
XSTDFILL51_32 VDD VSS sg13g2_FILL8
XSTDFILL51_40 VDD VSS sg13g2_FILL8
XSTDFILL51_48 VDD VSS sg13g2_FILL8
XSTDFILL51_56 VDD VSS sg13g2_FILL8
XSTDFILL51_64 VDD VSS sg13g2_FILL8
XSTDFILL51_72 VDD VSS sg13g2_FILL8
XSTDFILL51_80 VDD VSS sg13g2_FILL8
XSTDFILL51_88 VDD VSS sg13g2_FILL8
XSTDFILL51_96 VDD VSS sg13g2_FILL8
XSTDFILL51_104 VDD VSS sg13g2_FILL8
XSTDFILL51_112 VDD VSS sg13g2_FILL8
XSTDFILL51_120 VDD VSS sg13g2_FILL8
XSTDFILL51_128 VDD VSS sg13g2_FILL4
XSTDFILL51_1835 VDD VSS sg13g2_FILL8
XSTDFILL51_1843 VDD VSS sg13g2_FILL8
XSTDFILL51_1851 VDD VSS sg13g2_FILL8
XSTDFILL51_1859 VDD VSS sg13g2_FILL8
XSTDFILL51_1867 VDD VSS sg13g2_FILL8
XSTDFILL51_1875 VDD VSS sg13g2_FILL8
XSTDFILL51_1883 VDD VSS sg13g2_FILL8
XSTDFILL51_1891 VDD VSS sg13g2_FILL8
XSTDFILL51_1899 VDD VSS sg13g2_FILL8
XSTDFILL51_1907 VDD VSS sg13g2_FILL8
XSTDFILL51_1915 VDD VSS sg13g2_FILL8
XSTDFILL51_1923 VDD VSS sg13g2_FILL8
XSTDFILL51_1931 VDD VSS sg13g2_FILL8
XSTDFILL51_1939 VDD VSS sg13g2_FILL8
XSTDFILL51_1947 VDD VSS sg13g2_FILL8
XSTDFILL51_1955 VDD VSS sg13g2_FILL8
XSTDFILL51_1963 VDD VSS sg13g2_FILL8
XSTDFILL51_1971 VDD VSS sg13g2_FILL8
XSTDFILL51_1979 VDD VSS sg13g2_FILL8
XSTDFILL51_1987 VDD VSS sg13g2_FILL8
XSTDFILL51_1995 VDD VSS sg13g2_FILL8
XSTDFILL51_2003 VDD VSS sg13g2_FILL8
XSTDFILL51_2011 VDD VSS sg13g2_FILL8
XSTDFILL51_2019 VDD VSS sg13g2_FILL8
XSTDFILL51_2027 VDD VSS sg13g2_FILL8
XSTDFILL51_2035 VDD VSS sg13g2_FILL8
XSTDFILL51_2043 VDD VSS sg13g2_FILL8
XSTDFILL51_2051 VDD VSS sg13g2_FILL8
XSTDFILL51_2059 VDD VSS sg13g2_FILL8
XSTDFILL51_2067 VDD VSS sg13g2_FILL8
XSTDFILL51_2075 VDD VSS sg13g2_FILL8
XSTDFILL51_2083 VDD VSS sg13g2_FILL8
XSTDFILL51_2091 VDD VSS sg13g2_FILL8
XSTDFILL51_2099 VDD VSS sg13g2_FILL8
XSTDFILL51_2107 VDD VSS sg13g2_FILL8
XSTDFILL51_2115 VDD VSS sg13g2_FILL8
XSTDFILL51_2123 VDD VSS sg13g2_FILL8
XSTDFILL51_2131 VDD VSS sg13g2_FILL8
XSTDFILL51_2139 VDD VSS sg13g2_FILL8
XSTDFILL51_2147 VDD VSS sg13g2_FILL4
XSTDFILL51_2151 VDD VSS sg13g2_FILL2
XSTDFILL51_2153 VDD VSS sg13g2_FILL1
XSTDFILL52_0 VDD VSS sg13g2_FILL8
XSTDFILL52_8 VDD VSS sg13g2_FILL8
XSTDFILL52_16 VDD VSS sg13g2_FILL8
XSTDFILL52_24 VDD VSS sg13g2_FILL8
XSTDFILL52_32 VDD VSS sg13g2_FILL8
XSTDFILL52_40 VDD VSS sg13g2_FILL8
XSTDFILL52_48 VDD VSS sg13g2_FILL8
XSTDFILL52_56 VDD VSS sg13g2_FILL8
XSTDFILL52_64 VDD VSS sg13g2_FILL8
XSTDFILL52_72 VDD VSS sg13g2_FILL8
XSTDFILL52_80 VDD VSS sg13g2_FILL8
XSTDFILL52_88 VDD VSS sg13g2_FILL8
XSTDFILL52_96 VDD VSS sg13g2_FILL8
XSTDFILL52_104 VDD VSS sg13g2_FILL8
XSTDFILL52_112 VDD VSS sg13g2_FILL8
XSTDFILL52_120 VDD VSS sg13g2_FILL8
XSTDFILL52_128 VDD VSS sg13g2_FILL4
XSTDFILL52_1835 VDD VSS sg13g2_FILL8
XSTDFILL52_1843 VDD VSS sg13g2_FILL8
XSTDFILL52_1851 VDD VSS sg13g2_FILL8
XSTDFILL52_1859 VDD VSS sg13g2_FILL8
XSTDFILL52_1867 VDD VSS sg13g2_FILL8
XSTDFILL52_1875 VDD VSS sg13g2_FILL8
XSTDFILL52_1883 VDD VSS sg13g2_FILL8
XSTDFILL52_1891 VDD VSS sg13g2_FILL8
XSTDFILL52_1899 VDD VSS sg13g2_FILL8
XSTDFILL52_1907 VDD VSS sg13g2_FILL8
XSTDFILL52_1915 VDD VSS sg13g2_FILL8
XSTDFILL52_1923 VDD VSS sg13g2_FILL8
XSTDFILL52_1931 VDD VSS sg13g2_FILL8
XSTDFILL52_1939 VDD VSS sg13g2_FILL8
XSTDFILL52_1947 VDD VSS sg13g2_FILL8
XSTDFILL52_1955 VDD VSS sg13g2_FILL8
XSTDFILL52_1963 VDD VSS sg13g2_FILL8
XSTDFILL52_1971 VDD VSS sg13g2_FILL8
XSTDFILL52_1979 VDD VSS sg13g2_FILL8
XSTDFILL52_1987 VDD VSS sg13g2_FILL8
XSTDFILL52_1995 VDD VSS sg13g2_FILL8
XSTDFILL52_2003 VDD VSS sg13g2_FILL8
XSTDFILL52_2011 VDD VSS sg13g2_FILL8
XSTDFILL52_2019 VDD VSS sg13g2_FILL8
XSTDFILL52_2027 VDD VSS sg13g2_FILL8
XSTDFILL52_2035 VDD VSS sg13g2_FILL8
XSTDFILL52_2043 VDD VSS sg13g2_FILL8
XSTDFILL52_2051 VDD VSS sg13g2_FILL8
XSTDFILL52_2059 VDD VSS sg13g2_FILL8
XSTDFILL52_2067 VDD VSS sg13g2_FILL8
XSTDFILL52_2075 VDD VSS sg13g2_FILL8
XSTDFILL52_2083 VDD VSS sg13g2_FILL8
XSTDFILL52_2091 VDD VSS sg13g2_FILL8
XSTDFILL52_2099 VDD VSS sg13g2_FILL8
XSTDFILL52_2107 VDD VSS sg13g2_FILL8
XSTDFILL52_2115 VDD VSS sg13g2_FILL8
XSTDFILL52_2123 VDD VSS sg13g2_FILL8
XSTDFILL52_2131 VDD VSS sg13g2_FILL8
XSTDFILL52_2139 VDD VSS sg13g2_FILL8
XSTDFILL52_2147 VDD VSS sg13g2_FILL4
XSTDFILL52_2151 VDD VSS sg13g2_FILL2
XSTDFILL52_2153 VDD VSS sg13g2_FILL1
XSTDFILL53_0 VDD VSS sg13g2_FILL8
XSTDFILL53_8 VDD VSS sg13g2_FILL8
XSTDFILL53_16 VDD VSS sg13g2_FILL8
XSTDFILL53_24 VDD VSS sg13g2_FILL8
XSTDFILL53_32 VDD VSS sg13g2_FILL8
XSTDFILL53_40 VDD VSS sg13g2_FILL8
XSTDFILL53_48 VDD VSS sg13g2_FILL8
XSTDFILL53_56 VDD VSS sg13g2_FILL8
XSTDFILL53_64 VDD VSS sg13g2_FILL8
XSTDFILL53_72 VDD VSS sg13g2_FILL8
XSTDFILL53_80 VDD VSS sg13g2_FILL8
XSTDFILL53_88 VDD VSS sg13g2_FILL8
XSTDFILL53_96 VDD VSS sg13g2_FILL8
XSTDFILL53_104 VDD VSS sg13g2_FILL8
XSTDFILL53_112 VDD VSS sg13g2_FILL8
XSTDFILL53_120 VDD VSS sg13g2_FILL8
XSTDFILL53_128 VDD VSS sg13g2_FILL4
XSTDFILL53_1835 VDD VSS sg13g2_FILL8
XSTDFILL53_1843 VDD VSS sg13g2_FILL8
XSTDFILL53_1851 VDD VSS sg13g2_FILL8
XSTDFILL53_1859 VDD VSS sg13g2_FILL8
XSTDFILL53_1867 VDD VSS sg13g2_FILL8
XSTDFILL53_1875 VDD VSS sg13g2_FILL8
XSTDFILL53_1883 VDD VSS sg13g2_FILL8
XSTDFILL53_1891 VDD VSS sg13g2_FILL8
XSTDFILL53_1899 VDD VSS sg13g2_FILL8
XSTDFILL53_1907 VDD VSS sg13g2_FILL8
XSTDFILL53_1915 VDD VSS sg13g2_FILL8
XSTDFILL53_1923 VDD VSS sg13g2_FILL8
XSTDFILL53_1931 VDD VSS sg13g2_FILL8
XSTDFILL53_1939 VDD VSS sg13g2_FILL8
XSTDFILL53_1947 VDD VSS sg13g2_FILL8
XSTDFILL53_1955 VDD VSS sg13g2_FILL8
XSTDFILL53_1963 VDD VSS sg13g2_FILL8
XSTDFILL53_1971 VDD VSS sg13g2_FILL8
XSTDFILL53_1979 VDD VSS sg13g2_FILL8
XSTDFILL53_1987 VDD VSS sg13g2_FILL8
XSTDFILL53_1995 VDD VSS sg13g2_FILL8
XSTDFILL53_2003 VDD VSS sg13g2_FILL8
XSTDFILL53_2011 VDD VSS sg13g2_FILL8
XSTDFILL53_2019 VDD VSS sg13g2_FILL8
XSTDFILL53_2027 VDD VSS sg13g2_FILL8
XSTDFILL53_2035 VDD VSS sg13g2_FILL8
XSTDFILL53_2043 VDD VSS sg13g2_FILL8
XSTDFILL53_2051 VDD VSS sg13g2_FILL8
XSTDFILL53_2059 VDD VSS sg13g2_FILL8
XSTDFILL53_2067 VDD VSS sg13g2_FILL8
XSTDFILL53_2075 VDD VSS sg13g2_FILL8
XSTDFILL53_2083 VDD VSS sg13g2_FILL8
XSTDFILL53_2091 VDD VSS sg13g2_FILL8
XSTDFILL53_2099 VDD VSS sg13g2_FILL8
XSTDFILL53_2107 VDD VSS sg13g2_FILL8
XSTDFILL53_2115 VDD VSS sg13g2_FILL8
XSTDFILL53_2123 VDD VSS sg13g2_FILL8
XSTDFILL53_2131 VDD VSS sg13g2_FILL8
XSTDFILL53_2139 VDD VSS sg13g2_FILL8
XSTDFILL53_2147 VDD VSS sg13g2_FILL4
XSTDFILL53_2151 VDD VSS sg13g2_FILL2
XSTDFILL53_2153 VDD VSS sg13g2_FILL1
XSTDFILL54_0 VDD VSS sg13g2_FILL8
XSTDFILL54_8 VDD VSS sg13g2_FILL8
XSTDFILL54_16 VDD VSS sg13g2_FILL8
XSTDFILL54_24 VDD VSS sg13g2_FILL8
XSTDFILL54_32 VDD VSS sg13g2_FILL8
XSTDFILL54_40 VDD VSS sg13g2_FILL8
XSTDFILL54_48 VDD VSS sg13g2_FILL8
XSTDFILL54_56 VDD VSS sg13g2_FILL8
XSTDFILL54_64 VDD VSS sg13g2_FILL8
XSTDFILL54_72 VDD VSS sg13g2_FILL8
XSTDFILL54_80 VDD VSS sg13g2_FILL8
XSTDFILL54_88 VDD VSS sg13g2_FILL8
XSTDFILL54_96 VDD VSS sg13g2_FILL8
XSTDFILL54_104 VDD VSS sg13g2_FILL8
XSTDFILL54_112 VDD VSS sg13g2_FILL8
XSTDFILL54_120 VDD VSS sg13g2_FILL8
XSTDFILL54_128 VDD VSS sg13g2_FILL4
XSTDFILL54_1835 VDD VSS sg13g2_FILL8
XSTDFILL54_1843 VDD VSS sg13g2_FILL8
XSTDFILL54_1851 VDD VSS sg13g2_FILL8
XSTDFILL54_1859 VDD VSS sg13g2_FILL8
XSTDFILL54_1867 VDD VSS sg13g2_FILL8
XSTDFILL54_1875 VDD VSS sg13g2_FILL8
XSTDFILL54_1883 VDD VSS sg13g2_FILL8
XSTDFILL54_1891 VDD VSS sg13g2_FILL8
XSTDFILL54_1899 VDD VSS sg13g2_FILL8
XSTDFILL54_1907 VDD VSS sg13g2_FILL8
XSTDFILL54_1915 VDD VSS sg13g2_FILL8
XSTDFILL54_1923 VDD VSS sg13g2_FILL8
XSTDFILL54_1931 VDD VSS sg13g2_FILL8
XSTDFILL54_1939 VDD VSS sg13g2_FILL8
XSTDFILL54_1947 VDD VSS sg13g2_FILL8
XSTDFILL54_1955 VDD VSS sg13g2_FILL8
XSTDFILL54_1963 VDD VSS sg13g2_FILL8
XSTDFILL54_1971 VDD VSS sg13g2_FILL8
XSTDFILL54_1979 VDD VSS sg13g2_FILL8
XSTDFILL54_1987 VDD VSS sg13g2_FILL8
XSTDFILL54_1995 VDD VSS sg13g2_FILL8
XSTDFILL54_2003 VDD VSS sg13g2_FILL8
XSTDFILL54_2011 VDD VSS sg13g2_FILL8
XSTDFILL54_2019 VDD VSS sg13g2_FILL8
XSTDFILL54_2027 VDD VSS sg13g2_FILL8
XSTDFILL54_2035 VDD VSS sg13g2_FILL8
XSTDFILL54_2043 VDD VSS sg13g2_FILL8
XSTDFILL54_2051 VDD VSS sg13g2_FILL8
XSTDFILL54_2059 VDD VSS sg13g2_FILL8
XSTDFILL54_2067 VDD VSS sg13g2_FILL8
XSTDFILL54_2075 VDD VSS sg13g2_FILL8
XSTDFILL54_2083 VDD VSS sg13g2_FILL8
XSTDFILL54_2091 VDD VSS sg13g2_FILL8
XSTDFILL54_2099 VDD VSS sg13g2_FILL8
XSTDFILL54_2107 VDD VSS sg13g2_FILL8
XSTDFILL54_2115 VDD VSS sg13g2_FILL8
XSTDFILL54_2123 VDD VSS sg13g2_FILL8
XSTDFILL54_2131 VDD VSS sg13g2_FILL8
XSTDFILL54_2139 VDD VSS sg13g2_FILL8
XSTDFILL54_2147 VDD VSS sg13g2_FILL4
XSTDFILL54_2151 VDD VSS sg13g2_FILL2
XSTDFILL54_2153 VDD VSS sg13g2_FILL1
XSTDFILL55_0 VDD VSS sg13g2_FILL8
XSTDFILL55_8 VDD VSS sg13g2_FILL8
XSTDFILL55_16 VDD VSS sg13g2_FILL8
XSTDFILL55_24 VDD VSS sg13g2_FILL8
XSTDFILL55_32 VDD VSS sg13g2_FILL8
XSTDFILL55_40 VDD VSS sg13g2_FILL8
XSTDFILL55_48 VDD VSS sg13g2_FILL8
XSTDFILL55_56 VDD VSS sg13g2_FILL8
XSTDFILL55_64 VDD VSS sg13g2_FILL8
XSTDFILL55_72 VDD VSS sg13g2_FILL8
XSTDFILL55_80 VDD VSS sg13g2_FILL8
XSTDFILL55_88 VDD VSS sg13g2_FILL8
XSTDFILL55_96 VDD VSS sg13g2_FILL8
XSTDFILL55_104 VDD VSS sg13g2_FILL8
XSTDFILL55_112 VDD VSS sg13g2_FILL8
XSTDFILL55_120 VDD VSS sg13g2_FILL8
XSTDFILL55_128 VDD VSS sg13g2_FILL4
XSTDFILL55_1835 VDD VSS sg13g2_FILL8
XSTDFILL55_1843 VDD VSS sg13g2_FILL8
XSTDFILL55_1851 VDD VSS sg13g2_FILL8
XSTDFILL55_1859 VDD VSS sg13g2_FILL8
XSTDFILL55_1867 VDD VSS sg13g2_FILL8
XSTDFILL55_1875 VDD VSS sg13g2_FILL8
XSTDFILL55_1883 VDD VSS sg13g2_FILL8
XSTDFILL55_1891 VDD VSS sg13g2_FILL8
XSTDFILL55_1899 VDD VSS sg13g2_FILL8
XSTDFILL55_1907 VDD VSS sg13g2_FILL8
XSTDFILL55_1915 VDD VSS sg13g2_FILL8
XSTDFILL55_1923 VDD VSS sg13g2_FILL8
XSTDFILL55_1931 VDD VSS sg13g2_FILL8
XSTDFILL55_1939 VDD VSS sg13g2_FILL8
XSTDFILL55_1947 VDD VSS sg13g2_FILL8
XSTDFILL55_1955 VDD VSS sg13g2_FILL8
XSTDFILL55_1963 VDD VSS sg13g2_FILL8
XSTDFILL55_1971 VDD VSS sg13g2_FILL8
XSTDFILL55_1979 VDD VSS sg13g2_FILL8
XSTDFILL55_1987 VDD VSS sg13g2_FILL8
XSTDFILL55_1995 VDD VSS sg13g2_FILL8
XSTDFILL55_2003 VDD VSS sg13g2_FILL8
XSTDFILL55_2011 VDD VSS sg13g2_FILL8
XSTDFILL55_2019 VDD VSS sg13g2_FILL8
XSTDFILL55_2027 VDD VSS sg13g2_FILL8
XSTDFILL55_2035 VDD VSS sg13g2_FILL8
XSTDFILL55_2043 VDD VSS sg13g2_FILL8
XSTDFILL55_2051 VDD VSS sg13g2_FILL8
XSTDFILL55_2059 VDD VSS sg13g2_FILL8
XSTDFILL55_2067 VDD VSS sg13g2_FILL8
XSTDFILL55_2075 VDD VSS sg13g2_FILL8
XSTDFILL55_2083 VDD VSS sg13g2_FILL8
XSTDFILL55_2091 VDD VSS sg13g2_FILL8
XSTDFILL55_2099 VDD VSS sg13g2_FILL8
XSTDFILL55_2107 VDD VSS sg13g2_FILL8
XSTDFILL55_2115 VDD VSS sg13g2_FILL8
XSTDFILL55_2123 VDD VSS sg13g2_FILL8
XSTDFILL55_2131 VDD VSS sg13g2_FILL8
XSTDFILL55_2139 VDD VSS sg13g2_FILL8
XSTDFILL55_2147 VDD VSS sg13g2_FILL4
XSTDFILL55_2151 VDD VSS sg13g2_FILL2
XSTDFILL55_2153 VDD VSS sg13g2_FILL1
XSTDFILL56_0 VDD VSS sg13g2_FILL8
XSTDFILL56_8 VDD VSS sg13g2_FILL8
XSTDFILL56_16 VDD VSS sg13g2_FILL8
XSTDFILL56_24 VDD VSS sg13g2_FILL8
XSTDFILL56_32 VDD VSS sg13g2_FILL8
XSTDFILL56_40 VDD VSS sg13g2_FILL8
XSTDFILL56_48 VDD VSS sg13g2_FILL8
XSTDFILL56_56 VDD VSS sg13g2_FILL8
XSTDFILL56_64 VDD VSS sg13g2_FILL8
XSTDFILL56_72 VDD VSS sg13g2_FILL8
XSTDFILL56_80 VDD VSS sg13g2_FILL8
XSTDFILL56_88 VDD VSS sg13g2_FILL8
XSTDFILL56_96 VDD VSS sg13g2_FILL8
XSTDFILL56_104 VDD VSS sg13g2_FILL8
XSTDFILL56_112 VDD VSS sg13g2_FILL8
XSTDFILL56_120 VDD VSS sg13g2_FILL8
XSTDFILL56_128 VDD VSS sg13g2_FILL4
XSTDFILL56_1835 VDD VSS sg13g2_FILL8
XSTDFILL56_1843 VDD VSS sg13g2_FILL8
XSTDFILL56_1851 VDD VSS sg13g2_FILL8
XSTDFILL56_1859 VDD VSS sg13g2_FILL8
XSTDFILL56_1867 VDD VSS sg13g2_FILL8
XSTDFILL56_1875 VDD VSS sg13g2_FILL8
XSTDFILL56_1883 VDD VSS sg13g2_FILL8
XSTDFILL56_1891 VDD VSS sg13g2_FILL8
XSTDFILL56_1899 VDD VSS sg13g2_FILL8
XSTDFILL56_1907 VDD VSS sg13g2_FILL8
XSTDFILL56_1915 VDD VSS sg13g2_FILL8
XSTDFILL56_1923 VDD VSS sg13g2_FILL8
XSTDFILL56_1931 VDD VSS sg13g2_FILL8
XSTDFILL56_1939 VDD VSS sg13g2_FILL8
XSTDFILL56_1947 VDD VSS sg13g2_FILL8
XSTDFILL56_1955 VDD VSS sg13g2_FILL8
XSTDFILL56_1963 VDD VSS sg13g2_FILL8
XSTDFILL56_1971 VDD VSS sg13g2_FILL8
XSTDFILL56_1979 VDD VSS sg13g2_FILL8
XSTDFILL56_1987 VDD VSS sg13g2_FILL8
XSTDFILL56_1995 VDD VSS sg13g2_FILL8
XSTDFILL56_2003 VDD VSS sg13g2_FILL8
XSTDFILL56_2011 VDD VSS sg13g2_FILL8
XSTDFILL56_2019 VDD VSS sg13g2_FILL8
XSTDFILL56_2027 VDD VSS sg13g2_FILL8
XSTDFILL56_2035 VDD VSS sg13g2_FILL8
XSTDFILL56_2043 VDD VSS sg13g2_FILL8
XSTDFILL56_2051 VDD VSS sg13g2_FILL8
XSTDFILL56_2059 VDD VSS sg13g2_FILL8
XSTDFILL56_2067 VDD VSS sg13g2_FILL8
XSTDFILL56_2075 VDD VSS sg13g2_FILL8
XSTDFILL56_2083 VDD VSS sg13g2_FILL8
XSTDFILL56_2091 VDD VSS sg13g2_FILL8
XSTDFILL56_2099 VDD VSS sg13g2_FILL8
XSTDFILL56_2107 VDD VSS sg13g2_FILL8
XSTDFILL56_2115 VDD VSS sg13g2_FILL8
XSTDFILL56_2123 VDD VSS sg13g2_FILL8
XSTDFILL56_2131 VDD VSS sg13g2_FILL8
XSTDFILL56_2139 VDD VSS sg13g2_FILL8
XSTDFILL56_2147 VDD VSS sg13g2_FILL4
XSTDFILL56_2151 VDD VSS sg13g2_FILL2
XSTDFILL56_2153 VDD VSS sg13g2_FILL1
XSTDFILL57_0 VDD VSS sg13g2_FILL8
XSTDFILL57_8 VDD VSS sg13g2_FILL8
XSTDFILL57_16 VDD VSS sg13g2_FILL8
XSTDFILL57_24 VDD VSS sg13g2_FILL8
XSTDFILL57_32 VDD VSS sg13g2_FILL8
XSTDFILL57_40 VDD VSS sg13g2_FILL8
XSTDFILL57_48 VDD VSS sg13g2_FILL8
XSTDFILL57_56 VDD VSS sg13g2_FILL8
XSTDFILL57_64 VDD VSS sg13g2_FILL8
XSTDFILL57_72 VDD VSS sg13g2_FILL8
XSTDFILL57_80 VDD VSS sg13g2_FILL8
XSTDFILL57_88 VDD VSS sg13g2_FILL8
XSTDFILL57_96 VDD VSS sg13g2_FILL8
XSTDFILL57_104 VDD VSS sg13g2_FILL8
XSTDFILL57_112 VDD VSS sg13g2_FILL8
XSTDFILL57_120 VDD VSS sg13g2_FILL8
XSTDFILL57_128 VDD VSS sg13g2_FILL4
XSTDFILL57_1835 VDD VSS sg13g2_FILL8
XSTDFILL57_1843 VDD VSS sg13g2_FILL8
XSTDFILL57_1851 VDD VSS sg13g2_FILL8
XSTDFILL57_1859 VDD VSS sg13g2_FILL8
XSTDFILL57_1867 VDD VSS sg13g2_FILL8
XSTDFILL57_1875 VDD VSS sg13g2_FILL8
XSTDFILL57_1883 VDD VSS sg13g2_FILL8
XSTDFILL57_1891 VDD VSS sg13g2_FILL8
XSTDFILL57_1899 VDD VSS sg13g2_FILL8
XSTDFILL57_1907 VDD VSS sg13g2_FILL8
XSTDFILL57_1915 VDD VSS sg13g2_FILL8
XSTDFILL57_1923 VDD VSS sg13g2_FILL8
XSTDFILL57_1931 VDD VSS sg13g2_FILL8
XSTDFILL57_1939 VDD VSS sg13g2_FILL8
XSTDFILL57_1947 VDD VSS sg13g2_FILL8
XSTDFILL57_1955 VDD VSS sg13g2_FILL8
XSTDFILL57_1963 VDD VSS sg13g2_FILL8
XSTDFILL57_1971 VDD VSS sg13g2_FILL8
XSTDFILL57_1979 VDD VSS sg13g2_FILL8
XSTDFILL57_1987 VDD VSS sg13g2_FILL8
XSTDFILL57_1995 VDD VSS sg13g2_FILL8
XSTDFILL57_2003 VDD VSS sg13g2_FILL8
XSTDFILL57_2011 VDD VSS sg13g2_FILL8
XSTDFILL57_2019 VDD VSS sg13g2_FILL8
XSTDFILL57_2027 VDD VSS sg13g2_FILL8
XSTDFILL57_2035 VDD VSS sg13g2_FILL8
XSTDFILL57_2043 VDD VSS sg13g2_FILL8
XSTDFILL57_2051 VDD VSS sg13g2_FILL8
XSTDFILL57_2059 VDD VSS sg13g2_FILL8
XSTDFILL57_2067 VDD VSS sg13g2_FILL8
XSTDFILL57_2075 VDD VSS sg13g2_FILL8
XSTDFILL57_2083 VDD VSS sg13g2_FILL8
XSTDFILL57_2091 VDD VSS sg13g2_FILL8
XSTDFILL57_2099 VDD VSS sg13g2_FILL8
XSTDFILL57_2107 VDD VSS sg13g2_FILL8
XSTDFILL57_2115 VDD VSS sg13g2_FILL8
XSTDFILL57_2123 VDD VSS sg13g2_FILL8
XSTDFILL57_2131 VDD VSS sg13g2_FILL8
XSTDFILL57_2139 VDD VSS sg13g2_FILL8
XSTDFILL57_2147 VDD VSS sg13g2_FILL4
XSTDFILL57_2151 VDD VSS sg13g2_FILL2
XSTDFILL57_2153 VDD VSS sg13g2_FILL1
XSTDFILL58_0 VDD VSS sg13g2_FILL8
XSTDFILL58_8 VDD VSS sg13g2_FILL8
XSTDFILL58_16 VDD VSS sg13g2_FILL8
XSTDFILL58_24 VDD VSS sg13g2_FILL8
XSTDFILL58_32 VDD VSS sg13g2_FILL8
XSTDFILL58_40 VDD VSS sg13g2_FILL8
XSTDFILL58_48 VDD VSS sg13g2_FILL8
XSTDFILL58_56 VDD VSS sg13g2_FILL8
XSTDFILL58_64 VDD VSS sg13g2_FILL8
XSTDFILL58_72 VDD VSS sg13g2_FILL8
XSTDFILL58_80 VDD VSS sg13g2_FILL8
XSTDFILL58_88 VDD VSS sg13g2_FILL8
XSTDFILL58_96 VDD VSS sg13g2_FILL8
XSTDFILL58_104 VDD VSS sg13g2_FILL8
XSTDFILL58_112 VDD VSS sg13g2_FILL8
XSTDFILL58_120 VDD VSS sg13g2_FILL8
XSTDFILL58_128 VDD VSS sg13g2_FILL4
XSTDFILL58_1835 VDD VSS sg13g2_FILL8
XSTDFILL58_1843 VDD VSS sg13g2_FILL8
XSTDFILL58_1851 VDD VSS sg13g2_FILL8
XSTDFILL58_1859 VDD VSS sg13g2_FILL8
XSTDFILL58_1867 VDD VSS sg13g2_FILL8
XSTDFILL58_1875 VDD VSS sg13g2_FILL8
XSTDFILL58_1883 VDD VSS sg13g2_FILL8
XSTDFILL58_1891 VDD VSS sg13g2_FILL8
XSTDFILL58_1899 VDD VSS sg13g2_FILL8
XSTDFILL58_1907 VDD VSS sg13g2_FILL8
XSTDFILL58_1915 VDD VSS sg13g2_FILL8
XSTDFILL58_1923 VDD VSS sg13g2_FILL8
XSTDFILL58_1931 VDD VSS sg13g2_FILL8
XSTDFILL58_1939 VDD VSS sg13g2_FILL8
XSTDFILL58_1947 VDD VSS sg13g2_FILL8
XSTDFILL58_1955 VDD VSS sg13g2_FILL8
XSTDFILL58_1963 VDD VSS sg13g2_FILL8
XSTDFILL58_1971 VDD VSS sg13g2_FILL8
XSTDFILL58_1979 VDD VSS sg13g2_FILL8
XSTDFILL58_1987 VDD VSS sg13g2_FILL8
XSTDFILL58_1995 VDD VSS sg13g2_FILL8
XSTDFILL58_2003 VDD VSS sg13g2_FILL8
XSTDFILL58_2011 VDD VSS sg13g2_FILL8
XSTDFILL58_2019 VDD VSS sg13g2_FILL8
XSTDFILL58_2027 VDD VSS sg13g2_FILL8
XSTDFILL58_2035 VDD VSS sg13g2_FILL8
XSTDFILL58_2043 VDD VSS sg13g2_FILL8
XSTDFILL58_2051 VDD VSS sg13g2_FILL8
XSTDFILL58_2059 VDD VSS sg13g2_FILL8
XSTDFILL58_2067 VDD VSS sg13g2_FILL8
XSTDFILL58_2075 VDD VSS sg13g2_FILL8
XSTDFILL58_2083 VDD VSS sg13g2_FILL8
XSTDFILL58_2091 VDD VSS sg13g2_FILL8
XSTDFILL58_2099 VDD VSS sg13g2_FILL8
XSTDFILL58_2107 VDD VSS sg13g2_FILL8
XSTDFILL58_2115 VDD VSS sg13g2_FILL8
XSTDFILL58_2123 VDD VSS sg13g2_FILL8
XSTDFILL58_2131 VDD VSS sg13g2_FILL8
XSTDFILL58_2139 VDD VSS sg13g2_FILL8
XSTDFILL58_2147 VDD VSS sg13g2_FILL4
XSTDFILL58_2151 VDD VSS sg13g2_FILL2
XSTDFILL58_2153 VDD VSS sg13g2_FILL1
XSTDFILL59_0 VDD VSS sg13g2_FILL8
XSTDFILL59_8 VDD VSS sg13g2_FILL8
XSTDFILL59_16 VDD VSS sg13g2_FILL8
XSTDFILL59_24 VDD VSS sg13g2_FILL8
XSTDFILL59_32 VDD VSS sg13g2_FILL8
XSTDFILL59_40 VDD VSS sg13g2_FILL8
XSTDFILL59_48 VDD VSS sg13g2_FILL8
XSTDFILL59_56 VDD VSS sg13g2_FILL8
XSTDFILL59_64 VDD VSS sg13g2_FILL8
XSTDFILL59_72 VDD VSS sg13g2_FILL8
XSTDFILL59_80 VDD VSS sg13g2_FILL8
XSTDFILL59_88 VDD VSS sg13g2_FILL8
XSTDFILL59_96 VDD VSS sg13g2_FILL8
XSTDFILL59_104 VDD VSS sg13g2_FILL8
XSTDFILL59_112 VDD VSS sg13g2_FILL8
XSTDFILL59_120 VDD VSS sg13g2_FILL8
XSTDFILL59_128 VDD VSS sg13g2_FILL4
XSTDFILL59_1835 VDD VSS sg13g2_FILL8
XSTDFILL59_1843 VDD VSS sg13g2_FILL8
XSTDFILL59_1851 VDD VSS sg13g2_FILL8
XSTDFILL59_1859 VDD VSS sg13g2_FILL8
XSTDFILL59_1867 VDD VSS sg13g2_FILL8
XSTDFILL59_1875 VDD VSS sg13g2_FILL8
XSTDFILL59_1883 VDD VSS sg13g2_FILL8
XSTDFILL59_1891 VDD VSS sg13g2_FILL8
XSTDFILL59_1899 VDD VSS sg13g2_FILL8
XSTDFILL59_1907 VDD VSS sg13g2_FILL8
XSTDFILL59_1915 VDD VSS sg13g2_FILL8
XSTDFILL59_1923 VDD VSS sg13g2_FILL8
XSTDFILL59_1931 VDD VSS sg13g2_FILL8
XSTDFILL59_1939 VDD VSS sg13g2_FILL8
XSTDFILL59_1947 VDD VSS sg13g2_FILL8
XSTDFILL59_1955 VDD VSS sg13g2_FILL8
XSTDFILL59_1963 VDD VSS sg13g2_FILL8
XSTDFILL59_1971 VDD VSS sg13g2_FILL8
XSTDFILL59_1979 VDD VSS sg13g2_FILL8
XSTDFILL59_1987 VDD VSS sg13g2_FILL8
XSTDFILL59_1995 VDD VSS sg13g2_FILL8
XSTDFILL59_2003 VDD VSS sg13g2_FILL8
XSTDFILL59_2011 VDD VSS sg13g2_FILL8
XSTDFILL59_2019 VDD VSS sg13g2_FILL8
XSTDFILL59_2027 VDD VSS sg13g2_FILL8
XSTDFILL59_2035 VDD VSS sg13g2_FILL8
XSTDFILL59_2043 VDD VSS sg13g2_FILL8
XSTDFILL59_2051 VDD VSS sg13g2_FILL8
XSTDFILL59_2059 VDD VSS sg13g2_FILL8
XSTDFILL59_2067 VDD VSS sg13g2_FILL8
XSTDFILL59_2075 VDD VSS sg13g2_FILL8
XSTDFILL59_2083 VDD VSS sg13g2_FILL8
XSTDFILL59_2091 VDD VSS sg13g2_FILL8
XSTDFILL59_2099 VDD VSS sg13g2_FILL8
XSTDFILL59_2107 VDD VSS sg13g2_FILL8
XSTDFILL59_2115 VDD VSS sg13g2_FILL8
XSTDFILL59_2123 VDD VSS sg13g2_FILL8
XSTDFILL59_2131 VDD VSS sg13g2_FILL8
XSTDFILL59_2139 VDD VSS sg13g2_FILL8
XSTDFILL59_2147 VDD VSS sg13g2_FILL4
XSTDFILL59_2151 VDD VSS sg13g2_FILL2
XSTDFILL59_2153 VDD VSS sg13g2_FILL1
XSTDFILL60_0 VDD VSS sg13g2_FILL8
XSTDFILL60_8 VDD VSS sg13g2_FILL8
XSTDFILL60_16 VDD VSS sg13g2_FILL8
XSTDFILL60_24 VDD VSS sg13g2_FILL8
XSTDFILL60_32 VDD VSS sg13g2_FILL8
XSTDFILL60_40 VDD VSS sg13g2_FILL8
XSTDFILL60_48 VDD VSS sg13g2_FILL8
XSTDFILL60_56 VDD VSS sg13g2_FILL8
XSTDFILL60_64 VDD VSS sg13g2_FILL8
XSTDFILL60_72 VDD VSS sg13g2_FILL8
XSTDFILL60_80 VDD VSS sg13g2_FILL8
XSTDFILL60_88 VDD VSS sg13g2_FILL8
XSTDFILL60_96 VDD VSS sg13g2_FILL8
XSTDFILL60_104 VDD VSS sg13g2_FILL8
XSTDFILL60_112 VDD VSS sg13g2_FILL8
XSTDFILL60_120 VDD VSS sg13g2_FILL8
XSTDFILL60_128 VDD VSS sg13g2_FILL4
XSTDFILL60_1835 VDD VSS sg13g2_FILL8
XSTDFILL60_1843 VDD VSS sg13g2_FILL8
XSTDFILL60_1851 VDD VSS sg13g2_FILL8
XSTDFILL60_1859 VDD VSS sg13g2_FILL8
XSTDFILL60_1867 VDD VSS sg13g2_FILL8
XSTDFILL60_1875 VDD VSS sg13g2_FILL8
XSTDFILL60_1883 VDD VSS sg13g2_FILL8
XSTDFILL60_1891 VDD VSS sg13g2_FILL8
XSTDFILL60_1899 VDD VSS sg13g2_FILL8
XSTDFILL60_1907 VDD VSS sg13g2_FILL8
XSTDFILL60_1915 VDD VSS sg13g2_FILL8
XSTDFILL60_1923 VDD VSS sg13g2_FILL8
XSTDFILL60_1931 VDD VSS sg13g2_FILL8
XSTDFILL60_1939 VDD VSS sg13g2_FILL8
XSTDFILL60_1947 VDD VSS sg13g2_FILL8
XSTDFILL60_1955 VDD VSS sg13g2_FILL8
XSTDFILL60_1963 VDD VSS sg13g2_FILL8
XSTDFILL60_1971 VDD VSS sg13g2_FILL8
XSTDFILL60_1979 VDD VSS sg13g2_FILL8
XSTDFILL60_1987 VDD VSS sg13g2_FILL8
XSTDFILL60_1995 VDD VSS sg13g2_FILL8
XSTDFILL60_2003 VDD VSS sg13g2_FILL8
XSTDFILL60_2011 VDD VSS sg13g2_FILL8
XSTDFILL60_2019 VDD VSS sg13g2_FILL8
XSTDFILL60_2027 VDD VSS sg13g2_FILL8
XSTDFILL60_2035 VDD VSS sg13g2_FILL8
XSTDFILL60_2043 VDD VSS sg13g2_FILL8
XSTDFILL60_2051 VDD VSS sg13g2_FILL8
XSTDFILL60_2059 VDD VSS sg13g2_FILL8
XSTDFILL60_2067 VDD VSS sg13g2_FILL8
XSTDFILL60_2075 VDD VSS sg13g2_FILL8
XSTDFILL60_2083 VDD VSS sg13g2_FILL8
XSTDFILL60_2091 VDD VSS sg13g2_FILL8
XSTDFILL60_2099 VDD VSS sg13g2_FILL8
XSTDFILL60_2107 VDD VSS sg13g2_FILL8
XSTDFILL60_2115 VDD VSS sg13g2_FILL8
XSTDFILL60_2123 VDD VSS sg13g2_FILL8
XSTDFILL60_2131 VDD VSS sg13g2_FILL8
XSTDFILL60_2139 VDD VSS sg13g2_FILL8
XSTDFILL60_2147 VDD VSS sg13g2_FILL4
XSTDFILL60_2151 VDD VSS sg13g2_FILL2
XSTDFILL60_2153 VDD VSS sg13g2_FILL1
XSTDFILL61_0 VDD VSS sg13g2_FILL8
XSTDFILL61_8 VDD VSS sg13g2_FILL8
XSTDFILL61_16 VDD VSS sg13g2_FILL8
XSTDFILL61_24 VDD VSS sg13g2_FILL8
XSTDFILL61_32 VDD VSS sg13g2_FILL8
XSTDFILL61_40 VDD VSS sg13g2_FILL8
XSTDFILL61_48 VDD VSS sg13g2_FILL8
XSTDFILL61_56 VDD VSS sg13g2_FILL8
XSTDFILL61_64 VDD VSS sg13g2_FILL8
XSTDFILL61_72 VDD VSS sg13g2_FILL8
XSTDFILL61_80 VDD VSS sg13g2_FILL8
XSTDFILL61_88 VDD VSS sg13g2_FILL8
XSTDFILL61_96 VDD VSS sg13g2_FILL8
XSTDFILL61_104 VDD VSS sg13g2_FILL8
XSTDFILL61_112 VDD VSS sg13g2_FILL8
XSTDFILL61_120 VDD VSS sg13g2_FILL8
XSTDFILL61_128 VDD VSS sg13g2_FILL8
XSTDFILL61_136 VDD VSS sg13g2_FILL8
XSTDFILL61_144 VDD VSS sg13g2_FILL8
XSTDFILL61_152 VDD VSS sg13g2_FILL8
XSTDFILL61_160 VDD VSS sg13g2_FILL8
XSTDFILL61_168 VDD VSS sg13g2_FILL8
XSTDFILL61_176 VDD VSS sg13g2_FILL8
XSTDFILL61_184 VDD VSS sg13g2_FILL8
XSTDFILL61_192 VDD VSS sg13g2_FILL8
XSTDFILL61_200 VDD VSS sg13g2_FILL8
XSTDFILL61_208 VDD VSS sg13g2_FILL8
XSTDFILL61_216 VDD VSS sg13g2_FILL8
XSTDFILL61_224 VDD VSS sg13g2_FILL8
XSTDFILL61_232 VDD VSS sg13g2_FILL8
XSTDFILL61_240 VDD VSS sg13g2_FILL8
XSTDFILL61_248 VDD VSS sg13g2_FILL8
XSTDFILL61_256 VDD VSS sg13g2_FILL8
XSTDFILL61_264 VDD VSS sg13g2_FILL8
XSTDFILL61_272 VDD VSS sg13g2_FILL8
XSTDFILL61_280 VDD VSS sg13g2_FILL8
XSTDFILL61_288 VDD VSS sg13g2_FILL8
XSTDFILL61_296 VDD VSS sg13g2_FILL8
XSTDFILL61_304 VDD VSS sg13g2_FILL8
XSTDFILL61_312 VDD VSS sg13g2_FILL8
XSTDFILL61_320 VDD VSS sg13g2_FILL8
XSTDFILL61_328 VDD VSS sg13g2_FILL8
XSTDFILL61_336 VDD VSS sg13g2_FILL8
XSTDFILL61_344 VDD VSS sg13g2_FILL8
XSTDFILL61_352 VDD VSS sg13g2_FILL8
XSTDFILL61_360 VDD VSS sg13g2_FILL8
XSTDFILL61_368 VDD VSS sg13g2_FILL8
XSTDFILL61_376 VDD VSS sg13g2_FILL8
XSTDFILL61_384 VDD VSS sg13g2_FILL8
XSTDFILL61_392 VDD VSS sg13g2_FILL8
XSTDFILL61_400 VDD VSS sg13g2_FILL8
XSTDFILL61_408 VDD VSS sg13g2_FILL8
XSTDFILL61_416 VDD VSS sg13g2_FILL8
XSTDFILL61_424 VDD VSS sg13g2_FILL8
XSTDFILL61_432 VDD VSS sg13g2_FILL8
XSTDFILL61_440 VDD VSS sg13g2_FILL8
XSTDFILL61_448 VDD VSS sg13g2_FILL8
XSTDFILL61_456 VDD VSS sg13g2_FILL8
XSTDFILL61_464 VDD VSS sg13g2_FILL8
XSTDFILL61_472 VDD VSS sg13g2_FILL8
XSTDFILL61_480 VDD VSS sg13g2_FILL8
XSTDFILL61_488 VDD VSS sg13g2_FILL8
XSTDFILL61_496 VDD VSS sg13g2_FILL8
XSTDFILL61_504 VDD VSS sg13g2_FILL8
XSTDFILL61_512 VDD VSS sg13g2_FILL8
XSTDFILL61_520 VDD VSS sg13g2_FILL8
XSTDFILL61_528 VDD VSS sg13g2_FILL8
XSTDFILL61_536 VDD VSS sg13g2_FILL8
XSTDFILL61_544 VDD VSS sg13g2_FILL8
XSTDFILL61_552 VDD VSS sg13g2_FILL8
XSTDFILL61_560 VDD VSS sg13g2_FILL8
XSTDFILL61_568 VDD VSS sg13g2_FILL8
XSTDFILL61_576 VDD VSS sg13g2_FILL8
XSTDFILL61_584 VDD VSS sg13g2_FILL8
XSTDFILL61_592 VDD VSS sg13g2_FILL8
XSTDFILL61_600 VDD VSS sg13g2_FILL8
XSTDFILL61_608 VDD VSS sg13g2_FILL8
XSTDFILL61_616 VDD VSS sg13g2_FILL8
XSTDFILL61_624 VDD VSS sg13g2_FILL8
XSTDFILL61_632 VDD VSS sg13g2_FILL8
XSTDFILL61_640 VDD VSS sg13g2_FILL8
XSTDFILL61_648 VDD VSS sg13g2_FILL8
XSTDFILL61_656 VDD VSS sg13g2_FILL8
XSTDFILL61_664 VDD VSS sg13g2_FILL8
XSTDFILL61_672 VDD VSS sg13g2_FILL8
XSTDFILL61_680 VDD VSS sg13g2_FILL8
XSTDFILL61_688 VDD VSS sg13g2_FILL8
XSTDFILL61_696 VDD VSS sg13g2_FILL8
XSTDFILL61_704 VDD VSS sg13g2_FILL8
XSTDFILL61_712 VDD VSS sg13g2_FILL8
XSTDFILL61_720 VDD VSS sg13g2_FILL8
XSTDFILL61_728 VDD VSS sg13g2_FILL8
XSTDFILL61_736 VDD VSS sg13g2_FILL8
XSTDFILL61_744 VDD VSS sg13g2_FILL8
XSTDFILL61_752 VDD VSS sg13g2_FILL8
XSTDFILL61_760 VDD VSS sg13g2_FILL8
XSTDFILL61_768 VDD VSS sg13g2_FILL8
XSTDFILL61_776 VDD VSS sg13g2_FILL8
XSTDFILL61_784 VDD VSS sg13g2_FILL8
XSTDFILL61_792 VDD VSS sg13g2_FILL8
XSTDFILL61_800 VDD VSS sg13g2_FILL8
XSTDFILL61_808 VDD VSS sg13g2_FILL8
XSTDFILL61_816 VDD VSS sg13g2_FILL8
XSTDFILL61_824 VDD VSS sg13g2_FILL8
XSTDFILL61_832 VDD VSS sg13g2_FILL8
XSTDFILL61_840 VDD VSS sg13g2_FILL8
XSTDFILL61_848 VDD VSS sg13g2_FILL8
XSTDFILL61_856 VDD VSS sg13g2_FILL8
XSTDFILL61_864 VDD VSS sg13g2_FILL8
XSTDFILL61_872 VDD VSS sg13g2_FILL8
XSTDFILL61_880 VDD VSS sg13g2_FILL8
XSTDFILL61_888 VDD VSS sg13g2_FILL8
XSTDFILL61_896 VDD VSS sg13g2_FILL8
XSTDFILL61_904 VDD VSS sg13g2_FILL8
XSTDFILL61_912 VDD VSS sg13g2_FILL8
XSTDFILL61_920 VDD VSS sg13g2_FILL8
XSTDFILL61_928 VDD VSS sg13g2_FILL8
XSTDFILL61_936 VDD VSS sg13g2_FILL8
XSTDFILL61_944 VDD VSS sg13g2_FILL8
XSTDFILL61_952 VDD VSS sg13g2_FILL8
XSTDFILL61_960 VDD VSS sg13g2_FILL8
XSTDFILL61_968 VDD VSS sg13g2_FILL8
XSTDFILL61_976 VDD VSS sg13g2_FILL8
XSTDFILL61_984 VDD VSS sg13g2_FILL8
XSTDFILL61_992 VDD VSS sg13g2_FILL8
XSTDFILL61_1000 VDD VSS sg13g2_FILL8
XSTDFILL61_1008 VDD VSS sg13g2_FILL8
XSTDFILL61_1016 VDD VSS sg13g2_FILL8
XSTDFILL61_1024 VDD VSS sg13g2_FILL8
XSTDFILL61_1032 VDD VSS sg13g2_FILL8
XSTDFILL61_1040 VDD VSS sg13g2_FILL8
XSTDFILL61_1048 VDD VSS sg13g2_FILL8
XSTDFILL61_1056 VDD VSS sg13g2_FILL8
XSTDFILL61_1064 VDD VSS sg13g2_FILL8
XSTDFILL61_1072 VDD VSS sg13g2_FILL8
XSTDFILL61_1080 VDD VSS sg13g2_FILL8
XSTDFILL61_1088 VDD VSS sg13g2_FILL8
XSTDFILL61_1096 VDD VSS sg13g2_FILL8
XSTDFILL61_1104 VDD VSS sg13g2_FILL8
XSTDFILL61_1112 VDD VSS sg13g2_FILL8
XSTDFILL61_1120 VDD VSS sg13g2_FILL8
XSTDFILL61_1128 VDD VSS sg13g2_FILL8
XSTDFILL61_1136 VDD VSS sg13g2_FILL8
XSTDFILL61_1144 VDD VSS sg13g2_FILL8
XSTDFILL61_1152 VDD VSS sg13g2_FILL8
XSTDFILL61_1160 VDD VSS sg13g2_FILL8
XSTDFILL61_1168 VDD VSS sg13g2_FILL8
XSTDFILL61_1176 VDD VSS sg13g2_FILL8
XSTDFILL61_1192 VDD VSS sg13g2_FILL8
XSTDFILL61_1200 VDD VSS sg13g2_FILL8
XSTDFILL61_1208 VDD VSS sg13g2_FILL8
XSTDFILL61_1216 VDD VSS sg13g2_FILL8
XSTDFILL61_1224 VDD VSS sg13g2_FILL8
XSTDFILL61_1232 VDD VSS sg13g2_FILL8
XSTDFILL61_1240 VDD VSS sg13g2_FILL8
XSTDFILL61_1248 VDD VSS sg13g2_FILL8
XSTDFILL61_1256 VDD VSS sg13g2_FILL8
XSTDFILL61_1264 VDD VSS sg13g2_FILL8
XSTDFILL61_1272 VDD VSS sg13g2_FILL8
XSTDFILL61_1280 VDD VSS sg13g2_FILL8
XSTDFILL61_1288 VDD VSS sg13g2_FILL8
XSTDFILL61_1296 VDD VSS sg13g2_FILL8
XSTDFILL61_1304 VDD VSS sg13g2_FILL8
XSTDFILL61_1312 VDD VSS sg13g2_FILL4
XSTDFILL61_1316 VDD VSS sg13g2_FILL2
XSTDFILL61_1340 VDD VSS sg13g2_FILL8
XSTDFILL61_1348 VDD VSS sg13g2_FILL8
XSTDFILL61_1356 VDD VSS sg13g2_FILL8
XSTDFILL61_1364 VDD VSS sg13g2_FILL8
XSTDFILL61_1372 VDD VSS sg13g2_FILL8
XSTDFILL61_1380 VDD VSS sg13g2_FILL8
XSTDFILL61_1388 VDD VSS sg13g2_FILL8
XSTDFILL61_1396 VDD VSS sg13g2_FILL8
XSTDFILL61_1404 VDD VSS sg13g2_FILL8
XSTDFILL61_1412 VDD VSS sg13g2_FILL8
XSTDFILL61_1420 VDD VSS sg13g2_FILL8
XSTDFILL61_1428 VDD VSS sg13g2_FILL8
XSTDFILL61_1436 VDD VSS sg13g2_FILL8
XSTDFILL61_1444 VDD VSS sg13g2_FILL8
XSTDFILL61_1452 VDD VSS sg13g2_FILL8
XSTDFILL61_1460 VDD VSS sg13g2_FILL8
XSTDFILL61_1468 VDD VSS sg13g2_FILL8
XSTDFILL61_1476 VDD VSS sg13g2_FILL8
XSTDFILL61_1484 VDD VSS sg13g2_FILL8
XSTDFILL61_1492 VDD VSS sg13g2_FILL8
XSTDFILL61_1500 VDD VSS sg13g2_FILL8
XSTDFILL61_1508 VDD VSS sg13g2_FILL8
XSTDFILL61_1516 VDD VSS sg13g2_FILL8
XSTDFILL61_1524 VDD VSS sg13g2_FILL8
XSTDFILL61_1532 VDD VSS sg13g2_FILL8
XSTDFILL61_1540 VDD VSS sg13g2_FILL8
XSTDFILL61_1548 VDD VSS sg13g2_FILL8
XSTDFILL61_1556 VDD VSS sg13g2_FILL8
XSTDFILL61_1564 VDD VSS sg13g2_FILL8
XSTDFILL61_1572 VDD VSS sg13g2_FILL8
XSTDFILL61_1580 VDD VSS sg13g2_FILL8
XSTDFILL61_1588 VDD VSS sg13g2_FILL8
XSTDFILL61_1596 VDD VSS sg13g2_FILL8
XSTDFILL61_1604 VDD VSS sg13g2_FILL8
XSTDFILL61_1612 VDD VSS sg13g2_FILL8
XSTDFILL61_1620 VDD VSS sg13g2_FILL8
XSTDFILL61_1628 VDD VSS sg13g2_FILL8
XSTDFILL61_1636 VDD VSS sg13g2_FILL8
XSTDFILL61_1644 VDD VSS sg13g2_FILL8
XSTDFILL61_1652 VDD VSS sg13g2_FILL8
XSTDFILL61_1660 VDD VSS sg13g2_FILL8
XSTDFILL61_1668 VDD VSS sg13g2_FILL8
XSTDFILL61_1676 VDD VSS sg13g2_FILL8
XSTDFILL61_1684 VDD VSS sg13g2_FILL8
XSTDFILL61_1692 VDD VSS sg13g2_FILL8
XSTDFILL61_1700 VDD VSS sg13g2_FILL8
XSTDFILL61_1708 VDD VSS sg13g2_FILL8
XSTDFILL61_1716 VDD VSS sg13g2_FILL8
XSTDFILL61_1724 VDD VSS sg13g2_FILL8
XSTDFILL61_1732 VDD VSS sg13g2_FILL8
XSTDFILL61_1740 VDD VSS sg13g2_FILL8
XSTDFILL61_1748 VDD VSS sg13g2_FILL8
XSTDFILL61_1756 VDD VSS sg13g2_FILL8
XSTDFILL61_1764 VDD VSS sg13g2_FILL8
XSTDFILL61_1772 VDD VSS sg13g2_FILL8
XSTDFILL61_1780 VDD VSS sg13g2_FILL8
XSTDFILL61_1788 VDD VSS sg13g2_FILL8
XSTDFILL61_1796 VDD VSS sg13g2_FILL8
XSTDFILL61_1804 VDD VSS sg13g2_FILL8
XSTDFILL61_1812 VDD VSS sg13g2_FILL8
XSTDFILL61_1820 VDD VSS sg13g2_FILL8
XSTDFILL61_1828 VDD VSS sg13g2_FILL8
XSTDFILL61_1836 VDD VSS sg13g2_FILL8
XSTDFILL61_1844 VDD VSS sg13g2_FILL8
XSTDFILL61_1852 VDD VSS sg13g2_FILL8
XSTDFILL61_1860 VDD VSS sg13g2_FILL8
XSTDFILL61_1868 VDD VSS sg13g2_FILL8
XSTDFILL61_1876 VDD VSS sg13g2_FILL8
XSTDFILL61_1884 VDD VSS sg13g2_FILL8
XSTDFILL61_1892 VDD VSS sg13g2_FILL8
XSTDFILL61_1900 VDD VSS sg13g2_FILL8
XSTDFILL61_1908 VDD VSS sg13g2_FILL8
XSTDFILL61_1916 VDD VSS sg13g2_FILL8
XSTDFILL61_1924 VDD VSS sg13g2_FILL8
XSTDFILL61_1932 VDD VSS sg13g2_FILL8
XSTDFILL61_1940 VDD VSS sg13g2_FILL8
XSTDFILL61_1948 VDD VSS sg13g2_FILL8
XSTDFILL61_1956 VDD VSS sg13g2_FILL8
XSTDFILL61_1964 VDD VSS sg13g2_FILL8
XSTDFILL61_1972 VDD VSS sg13g2_FILL8
XSTDFILL61_1980 VDD VSS sg13g2_FILL8
XSTDFILL61_1988 VDD VSS sg13g2_FILL8
XSTDFILL61_1996 VDD VSS sg13g2_FILL8
XSTDFILL61_2004 VDD VSS sg13g2_FILL8
XSTDFILL61_2012 VDD VSS sg13g2_FILL8
XSTDFILL61_2020 VDD VSS sg13g2_FILL8
XSTDFILL61_2028 VDD VSS sg13g2_FILL8
XSTDFILL61_2036 VDD VSS sg13g2_FILL8
XSTDFILL61_2044 VDD VSS sg13g2_FILL8
XSTDFILL61_2052 VDD VSS sg13g2_FILL8
XSTDFILL61_2060 VDD VSS sg13g2_FILL8
XSTDFILL61_2068 VDD VSS sg13g2_FILL8
XSTDFILL61_2076 VDD VSS sg13g2_FILL8
XSTDFILL61_2084 VDD VSS sg13g2_FILL8
XSTDFILL61_2092 VDD VSS sg13g2_FILL8
XSTDFILL61_2100 VDD VSS sg13g2_FILL8
XSTDFILL61_2108 VDD VSS sg13g2_FILL8
XSTDFILL61_2116 VDD VSS sg13g2_FILL8
XSTDFILL61_2124 VDD VSS sg13g2_FILL8
XSTDFILL61_2132 VDD VSS sg13g2_FILL8
XSTDFILL61_2140 VDD VSS sg13g2_FILL8
XSTDFILL61_2148 VDD VSS sg13g2_FILL4
XSTDFILL61_2152 VDD VSS sg13g2_FILL2
XSTDFILL62_0 VDD VSS sg13g2_FILL8
XSTDFILL62_8 VDD VSS sg13g2_FILL8
XSTDFILL62_16 VDD VSS sg13g2_FILL8
XSTDFILL62_24 VDD VSS sg13g2_FILL8
XSTDFILL62_32 VDD VSS sg13g2_FILL8
XSTDFILL62_40 VDD VSS sg13g2_FILL8
XSTDFILL62_48 VDD VSS sg13g2_FILL8
XSTDFILL62_56 VDD VSS sg13g2_FILL8
XSTDFILL62_64 VDD VSS sg13g2_FILL8
XSTDFILL62_72 VDD VSS sg13g2_FILL8
XSTDFILL62_80 VDD VSS sg13g2_FILL8
XSTDFILL62_88 VDD VSS sg13g2_FILL8
XSTDFILL62_96 VDD VSS sg13g2_FILL8
XSTDFILL62_104 VDD VSS sg13g2_FILL8
XSTDFILL62_112 VDD VSS sg13g2_FILL8
XSTDFILL62_120 VDD VSS sg13g2_FILL8
XSTDFILL62_128 VDD VSS sg13g2_FILL8
XSTDFILL62_136 VDD VSS sg13g2_FILL8
XSTDFILL62_144 VDD VSS sg13g2_FILL8
XSTDFILL62_152 VDD VSS sg13g2_FILL8
XSTDFILL62_160 VDD VSS sg13g2_FILL8
XSTDFILL62_168 VDD VSS sg13g2_FILL8
XSTDFILL62_176 VDD VSS sg13g2_FILL8
XSTDFILL62_184 VDD VSS sg13g2_FILL8
XSTDFILL62_192 VDD VSS sg13g2_FILL8
XSTDFILL62_200 VDD VSS sg13g2_FILL8
XSTDFILL62_208 VDD VSS sg13g2_FILL8
XSTDFILL62_216 VDD VSS sg13g2_FILL8
XSTDFILL62_224 VDD VSS sg13g2_FILL8
XSTDFILL62_232 VDD VSS sg13g2_FILL8
XSTDFILL62_240 VDD VSS sg13g2_FILL8
XSTDFILL62_248 VDD VSS sg13g2_FILL8
XSTDFILL62_256 VDD VSS sg13g2_FILL8
XSTDFILL62_264 VDD VSS sg13g2_FILL8
XSTDFILL62_272 VDD VSS sg13g2_FILL8
XSTDFILL62_280 VDD VSS sg13g2_FILL8
XSTDFILL62_288 VDD VSS sg13g2_FILL8
XSTDFILL62_296 VDD VSS sg13g2_FILL8
XSTDFILL62_304 VDD VSS sg13g2_FILL8
XSTDFILL62_312 VDD VSS sg13g2_FILL8
XSTDFILL62_320 VDD VSS sg13g2_FILL8
XSTDFILL62_328 VDD VSS sg13g2_FILL8
XSTDFILL62_336 VDD VSS sg13g2_FILL8
XSTDFILL62_344 VDD VSS sg13g2_FILL8
XSTDFILL62_352 VDD VSS sg13g2_FILL8
XSTDFILL62_360 VDD VSS sg13g2_FILL8
XSTDFILL62_368 VDD VSS sg13g2_FILL8
XSTDFILL62_376 VDD VSS sg13g2_FILL8
XSTDFILL62_384 VDD VSS sg13g2_FILL8
XSTDFILL62_392 VDD VSS sg13g2_FILL8
XSTDFILL62_400 VDD VSS sg13g2_FILL8
XSTDFILL62_408 VDD VSS sg13g2_FILL8
XSTDFILL62_416 VDD VSS sg13g2_FILL8
XSTDFILL62_424 VDD VSS sg13g2_FILL8
XSTDFILL62_432 VDD VSS sg13g2_FILL8
XSTDFILL62_440 VDD VSS sg13g2_FILL8
XSTDFILL62_448 VDD VSS sg13g2_FILL8
XSTDFILL62_456 VDD VSS sg13g2_FILL8
XSTDFILL62_464 VDD VSS sg13g2_FILL8
XSTDFILL62_472 VDD VSS sg13g2_FILL8
XSTDFILL62_480 VDD VSS sg13g2_FILL8
XSTDFILL62_488 VDD VSS sg13g2_FILL8
XSTDFILL62_496 VDD VSS sg13g2_FILL8
XSTDFILL62_504 VDD VSS sg13g2_FILL8
XSTDFILL62_512 VDD VSS sg13g2_FILL8
XSTDFILL62_520 VDD VSS sg13g2_FILL8
XSTDFILL62_528 VDD VSS sg13g2_FILL8
XSTDFILL62_536 VDD VSS sg13g2_FILL8
XSTDFILL62_544 VDD VSS sg13g2_FILL8
XSTDFILL62_552 VDD VSS sg13g2_FILL8
XSTDFILL62_560 VDD VSS sg13g2_FILL8
XSTDFILL62_568 VDD VSS sg13g2_FILL8
XSTDFILL62_576 VDD VSS sg13g2_FILL8
XSTDFILL62_584 VDD VSS sg13g2_FILL8
XSTDFILL62_592 VDD VSS sg13g2_FILL8
XSTDFILL62_600 VDD VSS sg13g2_FILL8
XSTDFILL62_608 VDD VSS sg13g2_FILL8
XSTDFILL62_616 VDD VSS sg13g2_FILL8
XSTDFILL62_624 VDD VSS sg13g2_FILL8
XSTDFILL62_632 VDD VSS sg13g2_FILL8
XSTDFILL62_640 VDD VSS sg13g2_FILL8
XSTDFILL62_648 VDD VSS sg13g2_FILL8
XSTDFILL62_656 VDD VSS sg13g2_FILL8
XSTDFILL62_664 VDD VSS sg13g2_FILL8
XSTDFILL62_672 VDD VSS sg13g2_FILL8
XSTDFILL62_680 VDD VSS sg13g2_FILL8
XSTDFILL62_688 VDD VSS sg13g2_FILL8
XSTDFILL62_696 VDD VSS sg13g2_FILL8
XSTDFILL62_704 VDD VSS sg13g2_FILL8
XSTDFILL62_712 VDD VSS sg13g2_FILL8
XSTDFILL62_720 VDD VSS sg13g2_FILL8
XSTDFILL62_728 VDD VSS sg13g2_FILL8
XSTDFILL62_736 VDD VSS sg13g2_FILL8
XSTDFILL62_744 VDD VSS sg13g2_FILL8
XSTDFILL62_752 VDD VSS sg13g2_FILL8
XSTDFILL62_760 VDD VSS sg13g2_FILL8
XSTDFILL62_768 VDD VSS sg13g2_FILL8
XSTDFILL62_776 VDD VSS sg13g2_FILL8
XSTDFILL62_784 VDD VSS sg13g2_FILL8
XSTDFILL62_792 VDD VSS sg13g2_FILL8
XSTDFILL62_800 VDD VSS sg13g2_FILL8
XSTDFILL62_808 VDD VSS sg13g2_FILL8
XSTDFILL62_816 VDD VSS sg13g2_FILL8
XSTDFILL62_824 VDD VSS sg13g2_FILL8
XSTDFILL62_832 VDD VSS sg13g2_FILL8
XSTDFILL62_840 VDD VSS sg13g2_FILL8
XSTDFILL62_848 VDD VSS sg13g2_FILL8
XSTDFILL62_856 VDD VSS sg13g2_FILL8
XSTDFILL62_864 VDD VSS sg13g2_FILL8
XSTDFILL62_872 VDD VSS sg13g2_FILL8
XSTDFILL62_880 VDD VSS sg13g2_FILL8
XSTDFILL62_888 VDD VSS sg13g2_FILL8
XSTDFILL62_896 VDD VSS sg13g2_FILL8
XSTDFILL62_904 VDD VSS sg13g2_FILL8
XSTDFILL62_912 VDD VSS sg13g2_FILL8
XSTDFILL62_920 VDD VSS sg13g2_FILL8
XSTDFILL62_928 VDD VSS sg13g2_FILL8
XSTDFILL62_936 VDD VSS sg13g2_FILL8
XSTDFILL62_944 VDD VSS sg13g2_FILL8
XSTDFILL62_952 VDD VSS sg13g2_FILL8
XSTDFILL62_960 VDD VSS sg13g2_FILL8
XSTDFILL62_968 VDD VSS sg13g2_FILL8
XSTDFILL62_976 VDD VSS sg13g2_FILL8
XSTDFILL62_984 VDD VSS sg13g2_FILL8
XSTDFILL62_992 VDD VSS sg13g2_FILL8
XSTDFILL62_1000 VDD VSS sg13g2_FILL8
XSTDFILL62_1008 VDD VSS sg13g2_FILL8
XSTDFILL62_1016 VDD VSS sg13g2_FILL8
XSTDFILL62_1024 VDD VSS sg13g2_FILL8
XSTDFILL62_1032 VDD VSS sg13g2_FILL8
XSTDFILL62_1040 VDD VSS sg13g2_FILL8
XSTDFILL62_1048 VDD VSS sg13g2_FILL8
XSTDFILL62_1056 VDD VSS sg13g2_FILL8
XSTDFILL62_1064 VDD VSS sg13g2_FILL8
XSTDFILL62_1072 VDD VSS sg13g2_FILL8
XSTDFILL62_1080 VDD VSS sg13g2_FILL8
XSTDFILL62_1088 VDD VSS sg13g2_FILL8
XSTDFILL62_1096 VDD VSS sg13g2_FILL8
XSTDFILL62_1104 VDD VSS sg13g2_FILL8
XSTDFILL62_1112 VDD VSS sg13g2_FILL8
XSTDFILL62_1120 VDD VSS sg13g2_FILL8
XSTDFILL62_1128 VDD VSS sg13g2_FILL8
XSTDFILL62_1136 VDD VSS sg13g2_FILL8
XSTDFILL62_1144 VDD VSS sg13g2_FILL8
XSTDFILL62_1152 VDD VSS sg13g2_FILL8
XSTDFILL62_1160 VDD VSS sg13g2_FILL8
XSTDFILL62_1168 VDD VSS sg13g2_FILL8
XSTDFILL62_1176 VDD VSS sg13g2_FILL8
XSTDFILL62_1184 VDD VSS sg13g2_FILL8
XSTDFILL62_1192 VDD VSS sg13g2_FILL8
XSTDFILL62_1200 VDD VSS sg13g2_FILL8
XSTDFILL62_1208 VDD VSS sg13g2_FILL8
XSTDFILL62_1216 VDD VSS sg13g2_FILL8
XSTDFILL62_1224 VDD VSS sg13g2_FILL8
XSTDFILL62_1232 VDD VSS sg13g2_FILL8
XSTDFILL62_1240 VDD VSS sg13g2_FILL8
XSTDFILL62_1248 VDD VSS sg13g2_FILL8
XSTDFILL62_1256 VDD VSS sg13g2_FILL8
XSTDFILL62_1264 VDD VSS sg13g2_FILL8
XSTDFILL62_1272 VDD VSS sg13g2_FILL8
XSTDFILL62_1280 VDD VSS sg13g2_FILL8
XSTDFILL62_1288 VDD VSS sg13g2_FILL8
XSTDFILL62_1296 VDD VSS sg13g2_FILL8
XSTDFILL62_1304 VDD VSS sg13g2_FILL8
XSTDFILL62_1312 VDD VSS sg13g2_FILL8
XSTDFILL62_1320 VDD VSS sg13g2_FILL8
XSTDFILL62_1328 VDD VSS sg13g2_FILL8
XSTDFILL62_1336 VDD VSS sg13g2_FILL8
XSTDFILL62_1344 VDD VSS sg13g2_FILL8
XSTDFILL62_1352 VDD VSS sg13g2_FILL8
XSTDFILL62_1360 VDD VSS sg13g2_FILL8
XSTDFILL62_1368 VDD VSS sg13g2_FILL8
XSTDFILL62_1376 VDD VSS sg13g2_FILL8
XSTDFILL62_1384 VDD VSS sg13g2_FILL8
XSTDFILL62_1392 VDD VSS sg13g2_FILL8
XSTDFILL62_1400 VDD VSS sg13g2_FILL8
XSTDFILL62_1408 VDD VSS sg13g2_FILL8
XSTDFILL62_1416 VDD VSS sg13g2_FILL8
XSTDFILL62_1424 VDD VSS sg13g2_FILL8
XSTDFILL62_1432 VDD VSS sg13g2_FILL8
XSTDFILL62_1440 VDD VSS sg13g2_FILL8
XSTDFILL62_1448 VDD VSS sg13g2_FILL8
XSTDFILL62_1456 VDD VSS sg13g2_FILL8
XSTDFILL62_1464 VDD VSS sg13g2_FILL8
XSTDFILL62_1472 VDD VSS sg13g2_FILL8
XSTDFILL62_1480 VDD VSS sg13g2_FILL8
XSTDFILL62_1488 VDD VSS sg13g2_FILL8
XSTDFILL62_1496 VDD VSS sg13g2_FILL8
XSTDFILL62_1504 VDD VSS sg13g2_FILL8
XSTDFILL62_1512 VDD VSS sg13g2_FILL8
XSTDFILL62_1520 VDD VSS sg13g2_FILL8
XSTDFILL62_1528 VDD VSS sg13g2_FILL8
XSTDFILL62_1536 VDD VSS sg13g2_FILL8
XSTDFILL62_1544 VDD VSS sg13g2_FILL8
XSTDFILL62_1552 VDD VSS sg13g2_FILL8
XSTDFILL62_1560 VDD VSS sg13g2_FILL8
XSTDFILL62_1568 VDD VSS sg13g2_FILL8
XSTDFILL62_1576 VDD VSS sg13g2_FILL8
XSTDFILL62_1584 VDD VSS sg13g2_FILL8
XSTDFILL62_1592 VDD VSS sg13g2_FILL8
XSTDFILL62_1600 VDD VSS sg13g2_FILL8
XSTDFILL62_1608 VDD VSS sg13g2_FILL8
XSTDFILL62_1616 VDD VSS sg13g2_FILL8
XSTDFILL62_1624 VDD VSS sg13g2_FILL8
XSTDFILL62_1632 VDD VSS sg13g2_FILL8
XSTDFILL62_1640 VDD VSS sg13g2_FILL8
XSTDFILL62_1648 VDD VSS sg13g2_FILL8
XSTDFILL62_1656 VDD VSS sg13g2_FILL8
XSTDFILL62_1664 VDD VSS sg13g2_FILL8
XSTDFILL62_1672 VDD VSS sg13g2_FILL8
XSTDFILL62_1680 VDD VSS sg13g2_FILL8
XSTDFILL62_1688 VDD VSS sg13g2_FILL8
XSTDFILL62_1696 VDD VSS sg13g2_FILL8
XSTDFILL62_1704 VDD VSS sg13g2_FILL8
XSTDFILL62_1712 VDD VSS sg13g2_FILL8
XSTDFILL62_1720 VDD VSS sg13g2_FILL8
XSTDFILL62_1728 VDD VSS sg13g2_FILL8
XSTDFILL62_1736 VDD VSS sg13g2_FILL8
XSTDFILL62_1744 VDD VSS sg13g2_FILL8
XSTDFILL62_1752 VDD VSS sg13g2_FILL8
XSTDFILL62_1760 VDD VSS sg13g2_FILL8
XSTDFILL62_1768 VDD VSS sg13g2_FILL8
XSTDFILL62_1776 VDD VSS sg13g2_FILL8
XSTDFILL62_1784 VDD VSS sg13g2_FILL8
XSTDFILL62_1792 VDD VSS sg13g2_FILL8
XSTDFILL62_1800 VDD VSS sg13g2_FILL8
XSTDFILL62_1808 VDD VSS sg13g2_FILL8
XSTDFILL62_1816 VDD VSS sg13g2_FILL8
XSTDFILL62_1824 VDD VSS sg13g2_FILL8
XSTDFILL62_1832 VDD VSS sg13g2_FILL8
XSTDFILL62_1840 VDD VSS sg13g2_FILL8
XSTDFILL62_1848 VDD VSS sg13g2_FILL8
XSTDFILL62_1856 VDD VSS sg13g2_FILL8
XSTDFILL62_1864 VDD VSS sg13g2_FILL8
XSTDFILL62_1872 VDD VSS sg13g2_FILL8
XSTDFILL62_1880 VDD VSS sg13g2_FILL8
XSTDFILL62_1888 VDD VSS sg13g2_FILL8
XSTDFILL62_1896 VDD VSS sg13g2_FILL8
XSTDFILL62_1904 VDD VSS sg13g2_FILL8
XSTDFILL62_1912 VDD VSS sg13g2_FILL8
XSTDFILL62_1920 VDD VSS sg13g2_FILL8
XSTDFILL62_1928 VDD VSS sg13g2_FILL8
XSTDFILL62_1936 VDD VSS sg13g2_FILL8
XSTDFILL62_1944 VDD VSS sg13g2_FILL8
XSTDFILL62_1952 VDD VSS sg13g2_FILL8
XSTDFILL62_1960 VDD VSS sg13g2_FILL8
XSTDFILL62_1968 VDD VSS sg13g2_FILL8
XSTDFILL62_1976 VDD VSS sg13g2_FILL8
XSTDFILL62_1984 VDD VSS sg13g2_FILL8
XSTDFILL62_1992 VDD VSS sg13g2_FILL8
XSTDFILL62_2000 VDD VSS sg13g2_FILL8
XSTDFILL62_2008 VDD VSS sg13g2_FILL8
XSTDFILL62_2016 VDD VSS sg13g2_FILL8
XSTDFILL62_2024 VDD VSS sg13g2_FILL8
XSTDFILL62_2032 VDD VSS sg13g2_FILL8
XSTDFILL62_2040 VDD VSS sg13g2_FILL8
XSTDFILL62_2048 VDD VSS sg13g2_FILL8
XSTDFILL62_2056 VDD VSS sg13g2_FILL8
XSTDFILL62_2064 VDD VSS sg13g2_FILL8
XSTDFILL62_2072 VDD VSS sg13g2_FILL8
XSTDFILL62_2080 VDD VSS sg13g2_FILL8
XSTDFILL62_2088 VDD VSS sg13g2_FILL8
XSTDFILL62_2096 VDD VSS sg13g2_FILL8
XSTDFILL62_2104 VDD VSS sg13g2_FILL8
XSTDFILL62_2112 VDD VSS sg13g2_FILL8
XSTDFILL62_2120 VDD VSS sg13g2_FILL8
XSTDFILL62_2128 VDD VSS sg13g2_FILL8
XSTDFILL62_2136 VDD VSS sg13g2_FILL8
XSTDFILL62_2144 VDD VSS sg13g2_FILL8
XSTDFILL62_2152 VDD VSS sg13g2_FILL2
XSTDFILL63_0 VDD VSS sg13g2_FILL8
XSTDFILL63_8 VDD VSS sg13g2_FILL8
XSTDFILL63_16 VDD VSS sg13g2_FILL8
XSTDFILL63_24 VDD VSS sg13g2_FILL8
XSTDFILL63_32 VDD VSS sg13g2_FILL8
XSTDFILL63_40 VDD VSS sg13g2_FILL8
XSTDFILL63_48 VDD VSS sg13g2_FILL8
XSTDFILL63_56 VDD VSS sg13g2_FILL8
XSTDFILL63_64 VDD VSS sg13g2_FILL8
XSTDFILL63_72 VDD VSS sg13g2_FILL8
XSTDFILL63_80 VDD VSS sg13g2_FILL8
XSTDFILL63_88 VDD VSS sg13g2_FILL8
XSTDFILL63_96 VDD VSS sg13g2_FILL8
XSTDFILL63_104 VDD VSS sg13g2_FILL8
XSTDFILL63_112 VDD VSS sg13g2_FILL8
XSTDFILL63_120 VDD VSS sg13g2_FILL8
XSTDFILL63_128 VDD VSS sg13g2_FILL8
XSTDFILL63_136 VDD VSS sg13g2_FILL8
XSTDFILL63_144 VDD VSS sg13g2_FILL8
XSTDFILL63_152 VDD VSS sg13g2_FILL8
XSTDFILL63_160 VDD VSS sg13g2_FILL8
XSTDFILL63_168 VDD VSS sg13g2_FILL8
XSTDFILL63_176 VDD VSS sg13g2_FILL8
XSTDFILL63_184 VDD VSS sg13g2_FILL8
XSTDFILL63_192 VDD VSS sg13g2_FILL8
XSTDFILL63_200 VDD VSS sg13g2_FILL8
XSTDFILL63_208 VDD VSS sg13g2_FILL8
XSTDFILL63_216 VDD VSS sg13g2_FILL8
XSTDFILL63_224 VDD VSS sg13g2_FILL8
XSTDFILL63_232 VDD VSS sg13g2_FILL8
XSTDFILL63_240 VDD VSS sg13g2_FILL8
XSTDFILL63_248 VDD VSS sg13g2_FILL8
XSTDFILL63_256 VDD VSS sg13g2_FILL8
XSTDFILL63_264 VDD VSS sg13g2_FILL8
XSTDFILL63_272 VDD VSS sg13g2_FILL8
XSTDFILL63_280 VDD VSS sg13g2_FILL8
XSTDFILL63_288 VDD VSS sg13g2_FILL8
XSTDFILL63_296 VDD VSS sg13g2_FILL8
XSTDFILL63_304 VDD VSS sg13g2_FILL8
XSTDFILL63_312 VDD VSS sg13g2_FILL8
XSTDFILL63_320 VDD VSS sg13g2_FILL8
XSTDFILL63_328 VDD VSS sg13g2_FILL8
XSTDFILL63_336 VDD VSS sg13g2_FILL8
XSTDFILL63_344 VDD VSS sg13g2_FILL8
XSTDFILL63_352 VDD VSS sg13g2_FILL8
XSTDFILL63_360 VDD VSS sg13g2_FILL8
XSTDFILL63_368 VDD VSS sg13g2_FILL8
XSTDFILL63_376 VDD VSS sg13g2_FILL8
XSTDFILL63_384 VDD VSS sg13g2_FILL8
XSTDFILL63_392 VDD VSS sg13g2_FILL8
XSTDFILL63_400 VDD VSS sg13g2_FILL8
XSTDFILL63_408 VDD VSS sg13g2_FILL8
XSTDFILL63_416 VDD VSS sg13g2_FILL8
XSTDFILL63_424 VDD VSS sg13g2_FILL8
XSTDFILL63_432 VDD VSS sg13g2_FILL8
XSTDFILL63_440 VDD VSS sg13g2_FILL8
XSTDFILL63_448 VDD VSS sg13g2_FILL8
XSTDFILL63_456 VDD VSS sg13g2_FILL8
XSTDFILL63_464 VDD VSS sg13g2_FILL8
XSTDFILL63_472 VDD VSS sg13g2_FILL8
XSTDFILL63_480 VDD VSS sg13g2_FILL8
XSTDFILL63_488 VDD VSS sg13g2_FILL8
XSTDFILL63_496 VDD VSS sg13g2_FILL8
XSTDFILL63_504 VDD VSS sg13g2_FILL8
XSTDFILL63_512 VDD VSS sg13g2_FILL8
XSTDFILL63_520 VDD VSS sg13g2_FILL8
XSTDFILL63_528 VDD VSS sg13g2_FILL8
XSTDFILL63_536 VDD VSS sg13g2_FILL8
XSTDFILL63_544 VDD VSS sg13g2_FILL8
XSTDFILL63_552 VDD VSS sg13g2_FILL8
XSTDFILL63_560 VDD VSS sg13g2_FILL8
XSTDFILL63_568 VDD VSS sg13g2_FILL8
XSTDFILL63_576 VDD VSS sg13g2_FILL8
XSTDFILL63_584 VDD VSS sg13g2_FILL8
XSTDFILL63_592 VDD VSS sg13g2_FILL8
XSTDFILL63_600 VDD VSS sg13g2_FILL8
XSTDFILL63_608 VDD VSS sg13g2_FILL8
XSTDFILL63_616 VDD VSS sg13g2_FILL8
XSTDFILL63_624 VDD VSS sg13g2_FILL8
XSTDFILL63_632 VDD VSS sg13g2_FILL8
XSTDFILL63_640 VDD VSS sg13g2_FILL8
XSTDFILL63_648 VDD VSS sg13g2_FILL8
XSTDFILL63_656 VDD VSS sg13g2_FILL8
XSTDFILL63_664 VDD VSS sg13g2_FILL8
XSTDFILL63_672 VDD VSS sg13g2_FILL8
XSTDFILL63_680 VDD VSS sg13g2_FILL8
XSTDFILL63_688 VDD VSS sg13g2_FILL8
XSTDFILL63_696 VDD VSS sg13g2_FILL8
XSTDFILL63_704 VDD VSS sg13g2_FILL8
XSTDFILL63_712 VDD VSS sg13g2_FILL8
XSTDFILL63_720 VDD VSS sg13g2_FILL8
XSTDFILL63_728 VDD VSS sg13g2_FILL8
XSTDFILL63_736 VDD VSS sg13g2_FILL8
XSTDFILL63_744 VDD VSS sg13g2_FILL8
XSTDFILL63_752 VDD VSS sg13g2_FILL8
XSTDFILL63_760 VDD VSS sg13g2_FILL8
XSTDFILL63_768 VDD VSS sg13g2_FILL8
XSTDFILL63_776 VDD VSS sg13g2_FILL8
XSTDFILL63_784 VDD VSS sg13g2_FILL8
XSTDFILL63_792 VDD VSS sg13g2_FILL8
XSTDFILL63_800 VDD VSS sg13g2_FILL8
XSTDFILL63_808 VDD VSS sg13g2_FILL8
XSTDFILL63_816 VDD VSS sg13g2_FILL8
XSTDFILL63_824 VDD VSS sg13g2_FILL8
XSTDFILL63_832 VDD VSS sg13g2_FILL8
XSTDFILL63_840 VDD VSS sg13g2_FILL8
XSTDFILL63_848 VDD VSS sg13g2_FILL8
XSTDFILL63_856 VDD VSS sg13g2_FILL8
XSTDFILL63_864 VDD VSS sg13g2_FILL8
XSTDFILL63_872 VDD VSS sg13g2_FILL8
XSTDFILL63_880 VDD VSS sg13g2_FILL8
XSTDFILL63_888 VDD VSS sg13g2_FILL8
XSTDFILL63_896 VDD VSS sg13g2_FILL8
XSTDFILL63_904 VDD VSS sg13g2_FILL8
XSTDFILL63_912 VDD VSS sg13g2_FILL8
XSTDFILL63_920 VDD VSS sg13g2_FILL8
XSTDFILL63_928 VDD VSS sg13g2_FILL8
XSTDFILL63_936 VDD VSS sg13g2_FILL8
XSTDFILL63_944 VDD VSS sg13g2_FILL8
XSTDFILL63_952 VDD VSS sg13g2_FILL8
XSTDFILL63_960 VDD VSS sg13g2_FILL8
XSTDFILL63_968 VDD VSS sg13g2_FILL8
XSTDFILL63_976 VDD VSS sg13g2_FILL8
XSTDFILL63_984 VDD VSS sg13g2_FILL8
XSTDFILL63_992 VDD VSS sg13g2_FILL8
XSTDFILL63_1000 VDD VSS sg13g2_FILL8
XSTDFILL63_1008 VDD VSS sg13g2_FILL8
XSTDFILL63_1016 VDD VSS sg13g2_FILL8
XSTDFILL63_1024 VDD VSS sg13g2_FILL8
XSTDFILL63_1032 VDD VSS sg13g2_FILL8
XSTDFILL63_1040 VDD VSS sg13g2_FILL8
XSTDFILL63_1048 VDD VSS sg13g2_FILL8
XSTDFILL63_1056 VDD VSS sg13g2_FILL8
XSTDFILL63_1064 VDD VSS sg13g2_FILL8
XSTDFILL63_1072 VDD VSS sg13g2_FILL8
XSTDFILL63_1080 VDD VSS sg13g2_FILL8
XSTDFILL63_1088 VDD VSS sg13g2_FILL8
XSTDFILL63_1096 VDD VSS sg13g2_FILL8
XSTDFILL63_1104 VDD VSS sg13g2_FILL8
XSTDFILL63_1112 VDD VSS sg13g2_FILL8
XSTDFILL63_1120 VDD VSS sg13g2_FILL8
XSTDFILL63_1128 VDD VSS sg13g2_FILL8
XSTDFILL63_1136 VDD VSS sg13g2_FILL8
XSTDFILL63_1144 VDD VSS sg13g2_FILL8
XSTDFILL63_1152 VDD VSS sg13g2_FILL8
XSTDFILL63_1160 VDD VSS sg13g2_FILL8
XSTDFILL63_1168 VDD VSS sg13g2_FILL8
XSTDFILL63_1176 VDD VSS sg13g2_FILL8
XSTDFILL63_1184 VDD VSS sg13g2_FILL8
XSTDFILL63_1192 VDD VSS sg13g2_FILL8
XSTDFILL63_1200 VDD VSS sg13g2_FILL8
XSTDFILL63_1208 VDD VSS sg13g2_FILL8
XSTDFILL63_1216 VDD VSS sg13g2_FILL8
XSTDFILL63_1224 VDD VSS sg13g2_FILL8
XSTDFILL63_1232 VDD VSS sg13g2_FILL8
XSTDFILL63_1240 VDD VSS sg13g2_FILL8
XSTDFILL63_1248 VDD VSS sg13g2_FILL8
XSTDFILL63_1256 VDD VSS sg13g2_FILL8
XSTDFILL63_1264 VDD VSS sg13g2_FILL8
XSTDFILL63_1272 VDD VSS sg13g2_FILL8
XSTDFILL63_1280 VDD VSS sg13g2_FILL8
XSTDFILL63_1288 VDD VSS sg13g2_FILL8
XSTDFILL63_1296 VDD VSS sg13g2_FILL8
XSTDFILL63_1304 VDD VSS sg13g2_FILL8
XSTDFILL63_1312 VDD VSS sg13g2_FILL8
XSTDFILL63_1320 VDD VSS sg13g2_FILL8
XSTDFILL63_1328 VDD VSS sg13g2_FILL8
XSTDFILL63_1336 VDD VSS sg13g2_FILL8
XSTDFILL63_1344 VDD VSS sg13g2_FILL8
XSTDFILL63_1352 VDD VSS sg13g2_FILL8
XSTDFILL63_1360 VDD VSS sg13g2_FILL8
XSTDFILL63_1368 VDD VSS sg13g2_FILL8
XSTDFILL63_1376 VDD VSS sg13g2_FILL8
XSTDFILL63_1384 VDD VSS sg13g2_FILL8
XSTDFILL63_1392 VDD VSS sg13g2_FILL8
XSTDFILL63_1400 VDD VSS sg13g2_FILL8
XSTDFILL63_1408 VDD VSS sg13g2_FILL8
XSTDFILL63_1416 VDD VSS sg13g2_FILL8
XSTDFILL63_1424 VDD VSS sg13g2_FILL8
XSTDFILL63_1432 VDD VSS sg13g2_FILL8
XSTDFILL63_1440 VDD VSS sg13g2_FILL8
XSTDFILL63_1448 VDD VSS sg13g2_FILL8
XSTDFILL63_1456 VDD VSS sg13g2_FILL8
XSTDFILL63_1464 VDD VSS sg13g2_FILL8
XSTDFILL63_1472 VDD VSS sg13g2_FILL8
XSTDFILL63_1480 VDD VSS sg13g2_FILL8
XSTDFILL63_1488 VDD VSS sg13g2_FILL8
XSTDFILL63_1496 VDD VSS sg13g2_FILL8
XSTDFILL63_1504 VDD VSS sg13g2_FILL8
XSTDFILL63_1512 VDD VSS sg13g2_FILL8
XSTDFILL63_1520 VDD VSS sg13g2_FILL8
XSTDFILL63_1528 VDD VSS sg13g2_FILL8
XSTDFILL63_1536 VDD VSS sg13g2_FILL8
XSTDFILL63_1544 VDD VSS sg13g2_FILL8
XSTDFILL63_1552 VDD VSS sg13g2_FILL8
XSTDFILL63_1560 VDD VSS sg13g2_FILL8
XSTDFILL63_1568 VDD VSS sg13g2_FILL8
XSTDFILL63_1576 VDD VSS sg13g2_FILL8
XSTDFILL63_1584 VDD VSS sg13g2_FILL8
XSTDFILL63_1592 VDD VSS sg13g2_FILL8
XSTDFILL63_1600 VDD VSS sg13g2_FILL8
XSTDFILL63_1608 VDD VSS sg13g2_FILL8
XSTDFILL63_1616 VDD VSS sg13g2_FILL8
XSTDFILL63_1624 VDD VSS sg13g2_FILL8
XSTDFILL63_1632 VDD VSS sg13g2_FILL8
XSTDFILL63_1640 VDD VSS sg13g2_FILL8
XSTDFILL63_1648 VDD VSS sg13g2_FILL8
XSTDFILL63_1656 VDD VSS sg13g2_FILL8
XSTDFILL63_1664 VDD VSS sg13g2_FILL8
XSTDFILL63_1672 VDD VSS sg13g2_FILL8
XSTDFILL63_1680 VDD VSS sg13g2_FILL8
XSTDFILL63_1688 VDD VSS sg13g2_FILL8
XSTDFILL63_1696 VDD VSS sg13g2_FILL8
XSTDFILL63_1704 VDD VSS sg13g2_FILL8
XSTDFILL63_1712 VDD VSS sg13g2_FILL8
XSTDFILL63_1720 VDD VSS sg13g2_FILL8
XSTDFILL63_1728 VDD VSS sg13g2_FILL8
XSTDFILL63_1736 VDD VSS sg13g2_FILL8
XSTDFILL63_1744 VDD VSS sg13g2_FILL8
XSTDFILL63_1752 VDD VSS sg13g2_FILL8
XSTDFILL63_1760 VDD VSS sg13g2_FILL8
XSTDFILL63_1768 VDD VSS sg13g2_FILL8
XSTDFILL63_1776 VDD VSS sg13g2_FILL8
XSTDFILL63_1784 VDD VSS sg13g2_FILL8
XSTDFILL63_1792 VDD VSS sg13g2_FILL8
XSTDFILL63_1800 VDD VSS sg13g2_FILL8
XSTDFILL63_1808 VDD VSS sg13g2_FILL8
XSTDFILL63_1816 VDD VSS sg13g2_FILL8
XSTDFILL63_1824 VDD VSS sg13g2_FILL8
XSTDFILL63_1832 VDD VSS sg13g2_FILL8
XSTDFILL63_1840 VDD VSS sg13g2_FILL8
XSTDFILL63_1848 VDD VSS sg13g2_FILL8
XSTDFILL63_1856 VDD VSS sg13g2_FILL8
XSTDFILL63_1864 VDD VSS sg13g2_FILL8
XSTDFILL63_1872 VDD VSS sg13g2_FILL8
XSTDFILL63_1880 VDD VSS sg13g2_FILL8
XSTDFILL63_1888 VDD VSS sg13g2_FILL8
XSTDFILL63_1896 VDD VSS sg13g2_FILL8
XSTDFILL63_1904 VDD VSS sg13g2_FILL8
XSTDFILL63_1912 VDD VSS sg13g2_FILL8
XSTDFILL63_1920 VDD VSS sg13g2_FILL8
XSTDFILL63_1928 VDD VSS sg13g2_FILL8
XSTDFILL63_1936 VDD VSS sg13g2_FILL8
XSTDFILL63_1944 VDD VSS sg13g2_FILL8
XSTDFILL63_1952 VDD VSS sg13g2_FILL8
XSTDFILL63_1960 VDD VSS sg13g2_FILL8
XSTDFILL63_1968 VDD VSS sg13g2_FILL8
XSTDFILL63_1976 VDD VSS sg13g2_FILL8
XSTDFILL63_1984 VDD VSS sg13g2_FILL8
XSTDFILL63_1992 VDD VSS sg13g2_FILL8
XSTDFILL63_2000 VDD VSS sg13g2_FILL8
XSTDFILL63_2008 VDD VSS sg13g2_FILL8
XSTDFILL63_2016 VDD VSS sg13g2_FILL8
XSTDFILL63_2024 VDD VSS sg13g2_FILL8
XSTDFILL63_2032 VDD VSS sg13g2_FILL8
XSTDFILL63_2040 VDD VSS sg13g2_FILL8
XSTDFILL63_2048 VDD VSS sg13g2_FILL8
XSTDFILL63_2056 VDD VSS sg13g2_FILL8
XSTDFILL63_2064 VDD VSS sg13g2_FILL8
XSTDFILL63_2072 VDD VSS sg13g2_FILL8
XSTDFILL63_2080 VDD VSS sg13g2_FILL8
XSTDFILL63_2088 VDD VSS sg13g2_FILL8
XSTDFILL63_2096 VDD VSS sg13g2_FILL8
XSTDFILL63_2104 VDD VSS sg13g2_FILL8
XSTDFILL63_2112 VDD VSS sg13g2_FILL8
XSTDFILL63_2120 VDD VSS sg13g2_FILL8
XSTDFILL63_2128 VDD VSS sg13g2_FILL8
XSTDFILL63_2136 VDD VSS sg13g2_FILL8
XSTDFILL63_2144 VDD VSS sg13g2_FILL8
XSTDFILL63_2152 VDD VSS sg13g2_FILL2
XSTDFILL64_0 VDD VSS sg13g2_FILL8
XSTDFILL64_8 VDD VSS sg13g2_FILL8
XSTDFILL64_16 VDD VSS sg13g2_FILL8
XSTDFILL64_24 VDD VSS sg13g2_FILL8
XSTDFILL64_32 VDD VSS sg13g2_FILL8
XSTDFILL64_40 VDD VSS sg13g2_FILL8
XSTDFILL64_48 VDD VSS sg13g2_FILL8
XSTDFILL64_56 VDD VSS sg13g2_FILL8
XSTDFILL64_64 VDD VSS sg13g2_FILL8
XSTDFILL64_72 VDD VSS sg13g2_FILL8
XSTDFILL64_80 VDD VSS sg13g2_FILL8
XSTDFILL64_88 VDD VSS sg13g2_FILL8
XSTDFILL64_96 VDD VSS sg13g2_FILL8
XSTDFILL64_104 VDD VSS sg13g2_FILL8
XSTDFILL64_112 VDD VSS sg13g2_FILL8
XSTDFILL64_120 VDD VSS sg13g2_FILL8
XSTDFILL64_128 VDD VSS sg13g2_FILL8
XSTDFILL64_136 VDD VSS sg13g2_FILL8
XSTDFILL64_144 VDD VSS sg13g2_FILL8
XSTDFILL64_152 VDD VSS sg13g2_FILL8
XSTDFILL64_160 VDD VSS sg13g2_FILL8
XSTDFILL64_168 VDD VSS sg13g2_FILL8
XSTDFILL64_176 VDD VSS sg13g2_FILL8
XSTDFILL64_184 VDD VSS sg13g2_FILL8
XSTDFILL64_192 VDD VSS sg13g2_FILL8
XSTDFILL64_200 VDD VSS sg13g2_FILL8
XSTDFILL64_208 VDD VSS sg13g2_FILL8
XSTDFILL64_216 VDD VSS sg13g2_FILL8
XSTDFILL64_224 VDD VSS sg13g2_FILL8
XSTDFILL64_232 VDD VSS sg13g2_FILL8
XSTDFILL64_240 VDD VSS sg13g2_FILL8
XSTDFILL64_248 VDD VSS sg13g2_FILL8
XSTDFILL64_256 VDD VSS sg13g2_FILL8
XSTDFILL64_264 VDD VSS sg13g2_FILL8
XSTDFILL64_272 VDD VSS sg13g2_FILL8
XSTDFILL64_280 VDD VSS sg13g2_FILL8
XSTDFILL64_288 VDD VSS sg13g2_FILL8
XSTDFILL64_296 VDD VSS sg13g2_FILL8
XSTDFILL64_304 VDD VSS sg13g2_FILL8
XSTDFILL64_312 VDD VSS sg13g2_FILL8
XSTDFILL64_320 VDD VSS sg13g2_FILL8
XSTDFILL64_328 VDD VSS sg13g2_FILL8
XSTDFILL64_336 VDD VSS sg13g2_FILL8
XSTDFILL64_344 VDD VSS sg13g2_FILL8
XSTDFILL64_352 VDD VSS sg13g2_FILL8
XSTDFILL64_360 VDD VSS sg13g2_FILL8
XSTDFILL64_368 VDD VSS sg13g2_FILL8
XSTDFILL64_376 VDD VSS sg13g2_FILL8
XSTDFILL64_384 VDD VSS sg13g2_FILL8
XSTDFILL64_392 VDD VSS sg13g2_FILL8
XSTDFILL64_400 VDD VSS sg13g2_FILL8
XSTDFILL64_408 VDD VSS sg13g2_FILL8
XSTDFILL64_416 VDD VSS sg13g2_FILL8
XSTDFILL64_424 VDD VSS sg13g2_FILL8
XSTDFILL64_432 VDD VSS sg13g2_FILL8
XSTDFILL64_440 VDD VSS sg13g2_FILL8
XSTDFILL64_448 VDD VSS sg13g2_FILL8
XSTDFILL64_456 VDD VSS sg13g2_FILL8
XSTDFILL64_464 VDD VSS sg13g2_FILL8
XSTDFILL64_472 VDD VSS sg13g2_FILL8
XSTDFILL64_480 VDD VSS sg13g2_FILL8
XSTDFILL64_488 VDD VSS sg13g2_FILL8
XSTDFILL64_496 VDD VSS sg13g2_FILL8
XSTDFILL64_504 VDD VSS sg13g2_FILL8
XSTDFILL64_512 VDD VSS sg13g2_FILL8
XSTDFILL64_520 VDD VSS sg13g2_FILL8
XSTDFILL64_528 VDD VSS sg13g2_FILL8
XSTDFILL64_536 VDD VSS sg13g2_FILL8
XSTDFILL64_544 VDD VSS sg13g2_FILL8
XSTDFILL64_552 VDD VSS sg13g2_FILL8
XSTDFILL64_560 VDD VSS sg13g2_FILL8
XSTDFILL64_568 VDD VSS sg13g2_FILL8
XSTDFILL64_576 VDD VSS sg13g2_FILL8
XSTDFILL64_584 VDD VSS sg13g2_FILL8
XSTDFILL64_592 VDD VSS sg13g2_FILL8
XSTDFILL64_600 VDD VSS sg13g2_FILL8
XSTDFILL64_608 VDD VSS sg13g2_FILL8
XSTDFILL64_616 VDD VSS sg13g2_FILL8
XSTDFILL64_624 VDD VSS sg13g2_FILL8
XSTDFILL64_632 VDD VSS sg13g2_FILL8
XSTDFILL64_640 VDD VSS sg13g2_FILL8
XSTDFILL64_648 VDD VSS sg13g2_FILL8
XSTDFILL64_656 VDD VSS sg13g2_FILL8
XSTDFILL64_664 VDD VSS sg13g2_FILL8
XSTDFILL64_672 VDD VSS sg13g2_FILL8
XSTDFILL64_680 VDD VSS sg13g2_FILL8
XSTDFILL64_688 VDD VSS sg13g2_FILL8
XSTDFILL64_696 VDD VSS sg13g2_FILL8
XSTDFILL64_704 VDD VSS sg13g2_FILL8
XSTDFILL64_712 VDD VSS sg13g2_FILL8
XSTDFILL64_720 VDD VSS sg13g2_FILL8
XSTDFILL64_728 VDD VSS sg13g2_FILL8
XSTDFILL64_736 VDD VSS sg13g2_FILL8
XSTDFILL64_744 VDD VSS sg13g2_FILL8
XSTDFILL64_752 VDD VSS sg13g2_FILL8
XSTDFILL64_760 VDD VSS sg13g2_FILL8
XSTDFILL64_768 VDD VSS sg13g2_FILL8
XSTDFILL64_776 VDD VSS sg13g2_FILL8
XSTDFILL64_784 VDD VSS sg13g2_FILL8
XSTDFILL64_792 VDD VSS sg13g2_FILL8
XSTDFILL64_800 VDD VSS sg13g2_FILL8
XSTDFILL64_808 VDD VSS sg13g2_FILL8
XSTDFILL64_816 VDD VSS sg13g2_FILL8
XSTDFILL64_824 VDD VSS sg13g2_FILL8
XSTDFILL64_832 VDD VSS sg13g2_FILL8
XSTDFILL64_840 VDD VSS sg13g2_FILL8
XSTDFILL64_848 VDD VSS sg13g2_FILL8
XSTDFILL64_856 VDD VSS sg13g2_FILL8
XSTDFILL64_864 VDD VSS sg13g2_FILL8
XSTDFILL64_872 VDD VSS sg13g2_FILL8
XSTDFILL64_880 VDD VSS sg13g2_FILL8
XSTDFILL64_888 VDD VSS sg13g2_FILL8
XSTDFILL64_896 VDD VSS sg13g2_FILL8
XSTDFILL64_904 VDD VSS sg13g2_FILL8
XSTDFILL64_912 VDD VSS sg13g2_FILL8
XSTDFILL64_920 VDD VSS sg13g2_FILL8
XSTDFILL64_928 VDD VSS sg13g2_FILL8
XSTDFILL64_936 VDD VSS sg13g2_FILL8
XSTDFILL64_944 VDD VSS sg13g2_FILL8
XSTDFILL64_952 VDD VSS sg13g2_FILL8
XSTDFILL64_960 VDD VSS sg13g2_FILL8
XSTDFILL64_968 VDD VSS sg13g2_FILL8
XSTDFILL64_976 VDD VSS sg13g2_FILL8
XSTDFILL64_984 VDD VSS sg13g2_FILL8
XSTDFILL64_992 VDD VSS sg13g2_FILL8
XSTDFILL64_1000 VDD VSS sg13g2_FILL8
XSTDFILL64_1008 VDD VSS sg13g2_FILL8
XSTDFILL64_1016 VDD VSS sg13g2_FILL8
XSTDFILL64_1024 VDD VSS sg13g2_FILL8
XSTDFILL64_1032 VDD VSS sg13g2_FILL8
XSTDFILL64_1040 VDD VSS sg13g2_FILL8
XSTDFILL64_1048 VDD VSS sg13g2_FILL8
XSTDFILL64_1056 VDD VSS sg13g2_FILL8
XSTDFILL64_1064 VDD VSS sg13g2_FILL8
XSTDFILL64_1072 VDD VSS sg13g2_FILL8
XSTDFILL64_1080 VDD VSS sg13g2_FILL8
XSTDFILL64_1088 VDD VSS sg13g2_FILL8
XSTDFILL64_1096 VDD VSS sg13g2_FILL8
XSTDFILL64_1104 VDD VSS sg13g2_FILL8
XSTDFILL64_1112 VDD VSS sg13g2_FILL8
XSTDFILL64_1120 VDD VSS sg13g2_FILL8
XSTDFILL64_1128 VDD VSS sg13g2_FILL8
XSTDFILL64_1136 VDD VSS sg13g2_FILL8
XSTDFILL64_1144 VDD VSS sg13g2_FILL8
XSTDFILL64_1152 VDD VSS sg13g2_FILL8
XSTDFILL64_1160 VDD VSS sg13g2_FILL8
XSTDFILL64_1168 VDD VSS sg13g2_FILL8
XSTDFILL64_1176 VDD VSS sg13g2_FILL8
XSTDFILL64_1184 VDD VSS sg13g2_FILL8
XSTDFILL64_1192 VDD VSS sg13g2_FILL8
XSTDFILL64_1200 VDD VSS sg13g2_FILL8
XSTDFILL64_1208 VDD VSS sg13g2_FILL8
XSTDFILL64_1216 VDD VSS sg13g2_FILL8
XSTDFILL64_1224 VDD VSS sg13g2_FILL8
XSTDFILL64_1232 VDD VSS sg13g2_FILL8
XSTDFILL64_1240 VDD VSS sg13g2_FILL8
XSTDFILL64_1248 VDD VSS sg13g2_FILL8
XSTDFILL64_1256 VDD VSS sg13g2_FILL8
XSTDFILL64_1264 VDD VSS sg13g2_FILL8
XSTDFILL64_1272 VDD VSS sg13g2_FILL8
XSTDFILL64_1280 VDD VSS sg13g2_FILL8
XSTDFILL64_1288 VDD VSS sg13g2_FILL8
XSTDFILL64_1296 VDD VSS sg13g2_FILL8
XSTDFILL64_1304 VDD VSS sg13g2_FILL8
XSTDFILL64_1312 VDD VSS sg13g2_FILL8
XSTDFILL64_1320 VDD VSS sg13g2_FILL8
XSTDFILL64_1328 VDD VSS sg13g2_FILL8
XSTDFILL64_1336 VDD VSS sg13g2_FILL8
XSTDFILL64_1344 VDD VSS sg13g2_FILL8
XSTDFILL64_1352 VDD VSS sg13g2_FILL8
XSTDFILL64_1360 VDD VSS sg13g2_FILL8
XSTDFILL64_1368 VDD VSS sg13g2_FILL8
XSTDFILL64_1376 VDD VSS sg13g2_FILL8
XSTDFILL64_1384 VDD VSS sg13g2_FILL8
XSTDFILL64_1392 VDD VSS sg13g2_FILL8
XSTDFILL64_1400 VDD VSS sg13g2_FILL8
XSTDFILL64_1408 VDD VSS sg13g2_FILL8
XSTDFILL64_1416 VDD VSS sg13g2_FILL8
XSTDFILL64_1424 VDD VSS sg13g2_FILL8
XSTDFILL64_1432 VDD VSS sg13g2_FILL8
XSTDFILL64_1440 VDD VSS sg13g2_FILL8
XSTDFILL64_1448 VDD VSS sg13g2_FILL8
XSTDFILL64_1456 VDD VSS sg13g2_FILL8
XSTDFILL64_1464 VDD VSS sg13g2_FILL8
XSTDFILL64_1472 VDD VSS sg13g2_FILL8
XSTDFILL64_1480 VDD VSS sg13g2_FILL8
XSTDFILL64_1488 VDD VSS sg13g2_FILL8
XSTDFILL64_1496 VDD VSS sg13g2_FILL8
XSTDFILL64_1504 VDD VSS sg13g2_FILL8
XSTDFILL64_1512 VDD VSS sg13g2_FILL8
XSTDFILL64_1520 VDD VSS sg13g2_FILL8
XSTDFILL64_1528 VDD VSS sg13g2_FILL8
XSTDFILL64_1536 VDD VSS sg13g2_FILL8
XSTDFILL64_1544 VDD VSS sg13g2_FILL8
XSTDFILL64_1552 VDD VSS sg13g2_FILL8
XSTDFILL64_1560 VDD VSS sg13g2_FILL8
XSTDFILL64_1568 VDD VSS sg13g2_FILL8
XSTDFILL64_1576 VDD VSS sg13g2_FILL8
XSTDFILL64_1584 VDD VSS sg13g2_FILL8
XSTDFILL64_1592 VDD VSS sg13g2_FILL8
XSTDFILL64_1600 VDD VSS sg13g2_FILL8
XSTDFILL64_1608 VDD VSS sg13g2_FILL8
XSTDFILL64_1616 VDD VSS sg13g2_FILL8
XSTDFILL64_1624 VDD VSS sg13g2_FILL8
XSTDFILL64_1632 VDD VSS sg13g2_FILL8
XSTDFILL64_1640 VDD VSS sg13g2_FILL8
XSTDFILL64_1648 VDD VSS sg13g2_FILL8
XSTDFILL64_1656 VDD VSS sg13g2_FILL8
XSTDFILL64_1664 VDD VSS sg13g2_FILL8
XSTDFILL64_1672 VDD VSS sg13g2_FILL8
XSTDFILL64_1680 VDD VSS sg13g2_FILL8
XSTDFILL64_1688 VDD VSS sg13g2_FILL8
XSTDFILL64_1696 VDD VSS sg13g2_FILL8
XSTDFILL64_1704 VDD VSS sg13g2_FILL8
XSTDFILL64_1712 VDD VSS sg13g2_FILL8
XSTDFILL64_1720 VDD VSS sg13g2_FILL8
XSTDFILL64_1728 VDD VSS sg13g2_FILL8
XSTDFILL64_1736 VDD VSS sg13g2_FILL8
XSTDFILL64_1744 VDD VSS sg13g2_FILL8
XSTDFILL64_1752 VDD VSS sg13g2_FILL8
XSTDFILL64_1760 VDD VSS sg13g2_FILL8
XSTDFILL64_1768 VDD VSS sg13g2_FILL8
XSTDFILL64_1776 VDD VSS sg13g2_FILL8
XSTDFILL64_1784 VDD VSS sg13g2_FILL8
XSTDFILL64_1792 VDD VSS sg13g2_FILL8
XSTDFILL64_1800 VDD VSS sg13g2_FILL8
XSTDFILL64_1808 VDD VSS sg13g2_FILL8
XSTDFILL64_1816 VDD VSS sg13g2_FILL8
XSTDFILL64_1824 VDD VSS sg13g2_FILL8
XSTDFILL64_1832 VDD VSS sg13g2_FILL8
XSTDFILL64_1840 VDD VSS sg13g2_FILL8
XSTDFILL64_1848 VDD VSS sg13g2_FILL8
XSTDFILL64_1856 VDD VSS sg13g2_FILL8
XSTDFILL64_1864 VDD VSS sg13g2_FILL8
XSTDFILL64_1872 VDD VSS sg13g2_FILL8
XSTDFILL64_1880 VDD VSS sg13g2_FILL8
XSTDFILL64_1888 VDD VSS sg13g2_FILL8
XSTDFILL64_1896 VDD VSS sg13g2_FILL8
XSTDFILL64_1904 VDD VSS sg13g2_FILL8
XSTDFILL64_1912 VDD VSS sg13g2_FILL8
XSTDFILL64_1920 VDD VSS sg13g2_FILL8
XSTDFILL64_1928 VDD VSS sg13g2_FILL8
XSTDFILL64_1936 VDD VSS sg13g2_FILL8
XSTDFILL64_1944 VDD VSS sg13g2_FILL8
XSTDFILL64_1952 VDD VSS sg13g2_FILL8
XSTDFILL64_1960 VDD VSS sg13g2_FILL8
XSTDFILL64_1968 VDD VSS sg13g2_FILL8
XSTDFILL64_1976 VDD VSS sg13g2_FILL8
XSTDFILL64_1984 VDD VSS sg13g2_FILL8
XSTDFILL64_1992 VDD VSS sg13g2_FILL8
XSTDFILL64_2000 VDD VSS sg13g2_FILL8
XSTDFILL64_2008 VDD VSS sg13g2_FILL8
XSTDFILL64_2016 VDD VSS sg13g2_FILL8
XSTDFILL64_2024 VDD VSS sg13g2_FILL8
XSTDFILL64_2032 VDD VSS sg13g2_FILL8
XSTDFILL64_2040 VDD VSS sg13g2_FILL8
XSTDFILL64_2048 VDD VSS sg13g2_FILL8
XSTDFILL64_2056 VDD VSS sg13g2_FILL8
XSTDFILL64_2064 VDD VSS sg13g2_FILL8
XSTDFILL64_2072 VDD VSS sg13g2_FILL8
XSTDFILL64_2080 VDD VSS sg13g2_FILL8
XSTDFILL64_2088 VDD VSS sg13g2_FILL8
XSTDFILL64_2096 VDD VSS sg13g2_FILL8
XSTDFILL64_2104 VDD VSS sg13g2_FILL8
XSTDFILL64_2112 VDD VSS sg13g2_FILL8
XSTDFILL64_2120 VDD VSS sg13g2_FILL8
XSTDFILL64_2128 VDD VSS sg13g2_FILL8
XSTDFILL64_2136 VDD VSS sg13g2_FILL8
XSTDFILL64_2144 VDD VSS sg13g2_FILL8
XSTDFILL64_2152 VDD VSS sg13g2_FILL2
XSTDFILL65_0 VDD VSS sg13g2_FILL8
XSTDFILL65_8 VDD VSS sg13g2_FILL8
XSTDFILL65_16 VDD VSS sg13g2_FILL8
XSTDFILL65_24 VDD VSS sg13g2_FILL8
XSTDFILL65_32 VDD VSS sg13g2_FILL8
XSTDFILL65_40 VDD VSS sg13g2_FILL8
XSTDFILL65_48 VDD VSS sg13g2_FILL8
XSTDFILL65_56 VDD VSS sg13g2_FILL8
XSTDFILL65_64 VDD VSS sg13g2_FILL8
XSTDFILL65_72 VDD VSS sg13g2_FILL8
XSTDFILL65_80 VDD VSS sg13g2_FILL8
XSTDFILL65_88 VDD VSS sg13g2_FILL8
XSTDFILL65_96 VDD VSS sg13g2_FILL8
XSTDFILL65_104 VDD VSS sg13g2_FILL8
XSTDFILL65_112 VDD VSS sg13g2_FILL8
XSTDFILL65_120 VDD VSS sg13g2_FILL8
XSTDFILL65_128 VDD VSS sg13g2_FILL8
XSTDFILL65_136 VDD VSS sg13g2_FILL8
XSTDFILL65_144 VDD VSS sg13g2_FILL8
XSTDFILL65_152 VDD VSS sg13g2_FILL8
XSTDFILL65_160 VDD VSS sg13g2_FILL8
XSTDFILL65_168 VDD VSS sg13g2_FILL8
XSTDFILL65_176 VDD VSS sg13g2_FILL8
XSTDFILL65_184 VDD VSS sg13g2_FILL8
XSTDFILL65_192 VDD VSS sg13g2_FILL8
XSTDFILL65_200 VDD VSS sg13g2_FILL8
XSTDFILL65_208 VDD VSS sg13g2_FILL8
XSTDFILL65_216 VDD VSS sg13g2_FILL8
XSTDFILL65_224 VDD VSS sg13g2_FILL8
XSTDFILL65_232 VDD VSS sg13g2_FILL8
XSTDFILL65_240 VDD VSS sg13g2_FILL8
XSTDFILL65_248 VDD VSS sg13g2_FILL8
XSTDFILL65_256 VDD VSS sg13g2_FILL8
XSTDFILL65_264 VDD VSS sg13g2_FILL8
XSTDFILL65_272 VDD VSS sg13g2_FILL8
XSTDFILL65_280 VDD VSS sg13g2_FILL8
XSTDFILL65_288 VDD VSS sg13g2_FILL8
XSTDFILL65_296 VDD VSS sg13g2_FILL8
XSTDFILL65_304 VDD VSS sg13g2_FILL8
XSTDFILL65_312 VDD VSS sg13g2_FILL8
XSTDFILL65_320 VDD VSS sg13g2_FILL8
XSTDFILL65_328 VDD VSS sg13g2_FILL8
XSTDFILL65_336 VDD VSS sg13g2_FILL8
XSTDFILL65_344 VDD VSS sg13g2_FILL8
XSTDFILL65_352 VDD VSS sg13g2_FILL8
XSTDFILL65_360 VDD VSS sg13g2_FILL8
XSTDFILL65_368 VDD VSS sg13g2_FILL8
XSTDFILL65_376 VDD VSS sg13g2_FILL8
XSTDFILL65_384 VDD VSS sg13g2_FILL8
XSTDFILL65_392 VDD VSS sg13g2_FILL8
XSTDFILL65_400 VDD VSS sg13g2_FILL8
XSTDFILL65_408 VDD VSS sg13g2_FILL8
XSTDFILL65_416 VDD VSS sg13g2_FILL8
XSTDFILL65_424 VDD VSS sg13g2_FILL8
XSTDFILL65_432 VDD VSS sg13g2_FILL8
XSTDFILL65_440 VDD VSS sg13g2_FILL8
XSTDFILL65_448 VDD VSS sg13g2_FILL8
XSTDFILL65_456 VDD VSS sg13g2_FILL8
XSTDFILL65_464 VDD VSS sg13g2_FILL8
XSTDFILL65_472 VDD VSS sg13g2_FILL8
XSTDFILL65_480 VDD VSS sg13g2_FILL8
XSTDFILL65_488 VDD VSS sg13g2_FILL8
XSTDFILL65_496 VDD VSS sg13g2_FILL8
XSTDFILL65_504 VDD VSS sg13g2_FILL8
XSTDFILL65_512 VDD VSS sg13g2_FILL8
XSTDFILL65_520 VDD VSS sg13g2_FILL8
XSTDFILL65_528 VDD VSS sg13g2_FILL8
XSTDFILL65_536 VDD VSS sg13g2_FILL8
XSTDFILL65_544 VDD VSS sg13g2_FILL8
XSTDFILL65_552 VDD VSS sg13g2_FILL8
XSTDFILL65_560 VDD VSS sg13g2_FILL8
XSTDFILL65_568 VDD VSS sg13g2_FILL8
XSTDFILL65_576 VDD VSS sg13g2_FILL8
XSTDFILL65_584 VDD VSS sg13g2_FILL8
XSTDFILL65_592 VDD VSS sg13g2_FILL8
XSTDFILL65_600 VDD VSS sg13g2_FILL8
XSTDFILL65_608 VDD VSS sg13g2_FILL8
XSTDFILL65_616 VDD VSS sg13g2_FILL8
XSTDFILL65_624 VDD VSS sg13g2_FILL8
XSTDFILL65_632 VDD VSS sg13g2_FILL8
XSTDFILL65_640 VDD VSS sg13g2_FILL8
XSTDFILL65_648 VDD VSS sg13g2_FILL8
XSTDFILL65_656 VDD VSS sg13g2_FILL8
XSTDFILL65_664 VDD VSS sg13g2_FILL8
XSTDFILL65_672 VDD VSS sg13g2_FILL8
XSTDFILL65_680 VDD VSS sg13g2_FILL8
XSTDFILL65_688 VDD VSS sg13g2_FILL8
XSTDFILL65_696 VDD VSS sg13g2_FILL8
XSTDFILL65_704 VDD VSS sg13g2_FILL8
XSTDFILL65_712 VDD VSS sg13g2_FILL8
XSTDFILL65_720 VDD VSS sg13g2_FILL8
XSTDFILL65_728 VDD VSS sg13g2_FILL8
XSTDFILL65_736 VDD VSS sg13g2_FILL8
XSTDFILL65_744 VDD VSS sg13g2_FILL8
XSTDFILL65_752 VDD VSS sg13g2_FILL8
XSTDFILL65_760 VDD VSS sg13g2_FILL8
XSTDFILL65_768 VDD VSS sg13g2_FILL8
XSTDFILL65_776 VDD VSS sg13g2_FILL8
XSTDFILL65_784 VDD VSS sg13g2_FILL8
XSTDFILL65_792 VDD VSS sg13g2_FILL8
XSTDFILL65_800 VDD VSS sg13g2_FILL8
XSTDFILL65_808 VDD VSS sg13g2_FILL8
XSTDFILL65_816 VDD VSS sg13g2_FILL8
XSTDFILL65_824 VDD VSS sg13g2_FILL8
XSTDFILL65_832 VDD VSS sg13g2_FILL8
XSTDFILL65_840 VDD VSS sg13g2_FILL8
XSTDFILL65_848 VDD VSS sg13g2_FILL8
XSTDFILL65_856 VDD VSS sg13g2_FILL8
XSTDFILL65_864 VDD VSS sg13g2_FILL8
XSTDFILL65_872 VDD VSS sg13g2_FILL8
XSTDFILL65_880 VDD VSS sg13g2_FILL8
XSTDFILL65_888 VDD VSS sg13g2_FILL8
XSTDFILL65_896 VDD VSS sg13g2_FILL8
XSTDFILL65_904 VDD VSS sg13g2_FILL8
XSTDFILL65_912 VDD VSS sg13g2_FILL8
XSTDFILL65_920 VDD VSS sg13g2_FILL8
XSTDFILL65_928 VDD VSS sg13g2_FILL8
XSTDFILL65_936 VDD VSS sg13g2_FILL8
XSTDFILL65_944 VDD VSS sg13g2_FILL8
XSTDFILL65_952 VDD VSS sg13g2_FILL8
XSTDFILL65_960 VDD VSS sg13g2_FILL8
XSTDFILL65_968 VDD VSS sg13g2_FILL8
XSTDFILL65_976 VDD VSS sg13g2_FILL8
XSTDFILL65_984 VDD VSS sg13g2_FILL8
XSTDFILL65_992 VDD VSS sg13g2_FILL8
XSTDFILL65_1000 VDD VSS sg13g2_FILL8
XSTDFILL65_1008 VDD VSS sg13g2_FILL8
XSTDFILL65_1016 VDD VSS sg13g2_FILL8
XSTDFILL65_1024 VDD VSS sg13g2_FILL8
XSTDFILL65_1032 VDD VSS sg13g2_FILL8
XSTDFILL65_1040 VDD VSS sg13g2_FILL8
XSTDFILL65_1048 VDD VSS sg13g2_FILL8
XSTDFILL65_1056 VDD VSS sg13g2_FILL8
XSTDFILL65_1064 VDD VSS sg13g2_FILL8
XSTDFILL65_1072 VDD VSS sg13g2_FILL8
XSTDFILL65_1080 VDD VSS sg13g2_FILL8
XSTDFILL65_1088 VDD VSS sg13g2_FILL8
XSTDFILL65_1096 VDD VSS sg13g2_FILL8
XSTDFILL65_1104 VDD VSS sg13g2_FILL8
XSTDFILL65_1112 VDD VSS sg13g2_FILL8
XSTDFILL65_1120 VDD VSS sg13g2_FILL8
XSTDFILL65_1128 VDD VSS sg13g2_FILL8
XSTDFILL65_1136 VDD VSS sg13g2_FILL8
XSTDFILL65_1144 VDD VSS sg13g2_FILL8
XSTDFILL65_1152 VDD VSS sg13g2_FILL8
XSTDFILL65_1160 VDD VSS sg13g2_FILL8
XSTDFILL65_1168 VDD VSS sg13g2_FILL8
XSTDFILL65_1176 VDD VSS sg13g2_FILL8
XSTDFILL65_1184 VDD VSS sg13g2_FILL8
XSTDFILL65_1192 VDD VSS sg13g2_FILL8
XSTDFILL65_1200 VDD VSS sg13g2_FILL8
XSTDFILL65_1208 VDD VSS sg13g2_FILL8
XSTDFILL65_1216 VDD VSS sg13g2_FILL8
XSTDFILL65_1224 VDD VSS sg13g2_FILL8
XSTDFILL65_1232 VDD VSS sg13g2_FILL8
XSTDFILL65_1240 VDD VSS sg13g2_FILL8
XSTDFILL65_1248 VDD VSS sg13g2_FILL8
XSTDFILL65_1256 VDD VSS sg13g2_FILL8
XSTDFILL65_1264 VDD VSS sg13g2_FILL8
XSTDFILL65_1272 VDD VSS sg13g2_FILL8
XSTDFILL65_1280 VDD VSS sg13g2_FILL8
XSTDFILL65_1288 VDD VSS sg13g2_FILL8
XSTDFILL65_1296 VDD VSS sg13g2_FILL8
XSTDFILL65_1304 VDD VSS sg13g2_FILL8
XSTDFILL65_1312 VDD VSS sg13g2_FILL8
XSTDFILL65_1320 VDD VSS sg13g2_FILL8
XSTDFILL65_1328 VDD VSS sg13g2_FILL8
XSTDFILL65_1336 VDD VSS sg13g2_FILL8
XSTDFILL65_1344 VDD VSS sg13g2_FILL8
XSTDFILL65_1352 VDD VSS sg13g2_FILL8
XSTDFILL65_1360 VDD VSS sg13g2_FILL8
XSTDFILL65_1368 VDD VSS sg13g2_FILL8
XSTDFILL65_1376 VDD VSS sg13g2_FILL8
XSTDFILL65_1384 VDD VSS sg13g2_FILL8
XSTDFILL65_1392 VDD VSS sg13g2_FILL8
XSTDFILL65_1400 VDD VSS sg13g2_FILL8
XSTDFILL65_1408 VDD VSS sg13g2_FILL8
XSTDFILL65_1416 VDD VSS sg13g2_FILL8
XSTDFILL65_1424 VDD VSS sg13g2_FILL8
XSTDFILL65_1432 VDD VSS sg13g2_FILL8
XSTDFILL65_1440 VDD VSS sg13g2_FILL8
XSTDFILL65_1448 VDD VSS sg13g2_FILL8
XSTDFILL65_1456 VDD VSS sg13g2_FILL8
XSTDFILL65_1464 VDD VSS sg13g2_FILL8
XSTDFILL65_1472 VDD VSS sg13g2_FILL8
XSTDFILL65_1480 VDD VSS sg13g2_FILL8
XSTDFILL65_1488 VDD VSS sg13g2_FILL8
XSTDFILL65_1496 VDD VSS sg13g2_FILL8
XSTDFILL65_1504 VDD VSS sg13g2_FILL8
XSTDFILL65_1512 VDD VSS sg13g2_FILL8
XSTDFILL65_1520 VDD VSS sg13g2_FILL8
XSTDFILL65_1528 VDD VSS sg13g2_FILL8
XSTDFILL65_1536 VDD VSS sg13g2_FILL8
XSTDFILL65_1544 VDD VSS sg13g2_FILL8
XSTDFILL65_1552 VDD VSS sg13g2_FILL8
XSTDFILL65_1560 VDD VSS sg13g2_FILL8
XSTDFILL65_1568 VDD VSS sg13g2_FILL8
XSTDFILL65_1576 VDD VSS sg13g2_FILL8
XSTDFILL65_1584 VDD VSS sg13g2_FILL8
XSTDFILL65_1592 VDD VSS sg13g2_FILL8
XSTDFILL65_1600 VDD VSS sg13g2_FILL8
XSTDFILL65_1608 VDD VSS sg13g2_FILL8
XSTDFILL65_1616 VDD VSS sg13g2_FILL8
XSTDFILL65_1624 VDD VSS sg13g2_FILL8
XSTDFILL65_1632 VDD VSS sg13g2_FILL8
XSTDFILL65_1640 VDD VSS sg13g2_FILL8
XSTDFILL65_1648 VDD VSS sg13g2_FILL8
XSTDFILL65_1656 VDD VSS sg13g2_FILL8
XSTDFILL65_1664 VDD VSS sg13g2_FILL8
XSTDFILL65_1672 VDD VSS sg13g2_FILL8
XSTDFILL65_1680 VDD VSS sg13g2_FILL8
XSTDFILL65_1688 VDD VSS sg13g2_FILL8
XSTDFILL65_1696 VDD VSS sg13g2_FILL8
XSTDFILL65_1704 VDD VSS sg13g2_FILL8
XSTDFILL65_1712 VDD VSS sg13g2_FILL8
XSTDFILL65_1720 VDD VSS sg13g2_FILL8
XSTDFILL65_1728 VDD VSS sg13g2_FILL8
XSTDFILL65_1736 VDD VSS sg13g2_FILL8
XSTDFILL65_1744 VDD VSS sg13g2_FILL8
XSTDFILL65_1752 VDD VSS sg13g2_FILL8
XSTDFILL65_1760 VDD VSS sg13g2_FILL8
XSTDFILL65_1768 VDD VSS sg13g2_FILL8
XSTDFILL65_1776 VDD VSS sg13g2_FILL8
XSTDFILL65_1784 VDD VSS sg13g2_FILL8
XSTDFILL65_1792 VDD VSS sg13g2_FILL8
XSTDFILL65_1800 VDD VSS sg13g2_FILL8
XSTDFILL65_1808 VDD VSS sg13g2_FILL8
XSTDFILL65_1816 VDD VSS sg13g2_FILL8
XSTDFILL65_1824 VDD VSS sg13g2_FILL8
XSTDFILL65_1832 VDD VSS sg13g2_FILL8
XSTDFILL65_1840 VDD VSS sg13g2_FILL8
XSTDFILL65_1848 VDD VSS sg13g2_FILL8
XSTDFILL65_1856 VDD VSS sg13g2_FILL8
XSTDFILL65_1864 VDD VSS sg13g2_FILL8
XSTDFILL65_1872 VDD VSS sg13g2_FILL8
XSTDFILL65_1880 VDD VSS sg13g2_FILL8
XSTDFILL65_1888 VDD VSS sg13g2_FILL8
XSTDFILL65_1896 VDD VSS sg13g2_FILL8
XSTDFILL65_1904 VDD VSS sg13g2_FILL8
XSTDFILL65_1912 VDD VSS sg13g2_FILL8
XSTDFILL65_1920 VDD VSS sg13g2_FILL8
XSTDFILL65_1928 VDD VSS sg13g2_FILL8
XSTDFILL65_1936 VDD VSS sg13g2_FILL8
XSTDFILL65_1944 VDD VSS sg13g2_FILL8
XSTDFILL65_1952 VDD VSS sg13g2_FILL8
XSTDFILL65_1960 VDD VSS sg13g2_FILL8
XSTDFILL65_1968 VDD VSS sg13g2_FILL8
XSTDFILL65_1976 VDD VSS sg13g2_FILL8
XSTDFILL65_1984 VDD VSS sg13g2_FILL8
XSTDFILL65_1992 VDD VSS sg13g2_FILL8
XSTDFILL65_2000 VDD VSS sg13g2_FILL8
XSTDFILL65_2008 VDD VSS sg13g2_FILL8
XSTDFILL65_2016 VDD VSS sg13g2_FILL8
XSTDFILL65_2024 VDD VSS sg13g2_FILL8
XSTDFILL65_2032 VDD VSS sg13g2_FILL8
XSTDFILL65_2040 VDD VSS sg13g2_FILL8
XSTDFILL65_2048 VDD VSS sg13g2_FILL8
XSTDFILL65_2056 VDD VSS sg13g2_FILL8
XSTDFILL65_2064 VDD VSS sg13g2_FILL8
XSTDFILL65_2072 VDD VSS sg13g2_FILL8
XSTDFILL65_2080 VDD VSS sg13g2_FILL8
XSTDFILL65_2088 VDD VSS sg13g2_FILL8
XSTDFILL65_2096 VDD VSS sg13g2_FILL8
XSTDFILL65_2104 VDD VSS sg13g2_FILL8
XSTDFILL65_2112 VDD VSS sg13g2_FILL8
XSTDFILL65_2120 VDD VSS sg13g2_FILL8
XSTDFILL65_2128 VDD VSS sg13g2_FILL8
XSTDFILL65_2136 VDD VSS sg13g2_FILL8
XSTDFILL65_2144 VDD VSS sg13g2_FILL8
XSTDFILL65_2152 VDD VSS sg13g2_FILL2
XSTDFILL66_0 VDD VSS sg13g2_FILL8
XSTDFILL66_8 VDD VSS sg13g2_FILL8
XSTDFILL66_16 VDD VSS sg13g2_FILL8
XSTDFILL66_24 VDD VSS sg13g2_FILL8
XSTDFILL66_32 VDD VSS sg13g2_FILL8
XSTDFILL66_40 VDD VSS sg13g2_FILL8
XSTDFILL66_48 VDD VSS sg13g2_FILL8
XSTDFILL66_56 VDD VSS sg13g2_FILL8
XSTDFILL66_64 VDD VSS sg13g2_FILL8
XSTDFILL66_72 VDD VSS sg13g2_FILL8
XSTDFILL66_80 VDD VSS sg13g2_FILL8
XSTDFILL66_88 VDD VSS sg13g2_FILL8
XSTDFILL66_96 VDD VSS sg13g2_FILL8
XSTDFILL66_104 VDD VSS sg13g2_FILL8
XSTDFILL66_112 VDD VSS sg13g2_FILL8
XSTDFILL66_120 VDD VSS sg13g2_FILL8
XSTDFILL66_128 VDD VSS sg13g2_FILL8
XSTDFILL66_136 VDD VSS sg13g2_FILL8
XSTDFILL66_144 VDD VSS sg13g2_FILL8
XSTDFILL66_152 VDD VSS sg13g2_FILL8
XSTDFILL66_160 VDD VSS sg13g2_FILL8
XSTDFILL66_168 VDD VSS sg13g2_FILL8
XSTDFILL66_176 VDD VSS sg13g2_FILL8
XSTDFILL66_184 VDD VSS sg13g2_FILL8
XSTDFILL66_192 VDD VSS sg13g2_FILL8
XSTDFILL66_200 VDD VSS sg13g2_FILL8
XSTDFILL66_208 VDD VSS sg13g2_FILL8
XSTDFILL66_216 VDD VSS sg13g2_FILL8
XSTDFILL66_224 VDD VSS sg13g2_FILL8
XSTDFILL66_232 VDD VSS sg13g2_FILL8
XSTDFILL66_240 VDD VSS sg13g2_FILL8
XSTDFILL66_248 VDD VSS sg13g2_FILL8
XSTDFILL66_256 VDD VSS sg13g2_FILL8
XSTDFILL66_264 VDD VSS sg13g2_FILL8
XSTDFILL66_272 VDD VSS sg13g2_FILL8
XSTDFILL66_280 VDD VSS sg13g2_FILL8
XSTDFILL66_288 VDD VSS sg13g2_FILL8
XSTDFILL66_296 VDD VSS sg13g2_FILL8
XSTDFILL66_304 VDD VSS sg13g2_FILL8
XSTDFILL66_312 VDD VSS sg13g2_FILL8
XSTDFILL66_320 VDD VSS sg13g2_FILL8
XSTDFILL66_328 VDD VSS sg13g2_FILL8
XSTDFILL66_336 VDD VSS sg13g2_FILL8
XSTDFILL66_344 VDD VSS sg13g2_FILL8
XSTDFILL66_352 VDD VSS sg13g2_FILL8
XSTDFILL66_360 VDD VSS sg13g2_FILL8
XSTDFILL66_368 VDD VSS sg13g2_FILL8
XSTDFILL66_376 VDD VSS sg13g2_FILL8
XSTDFILL66_384 VDD VSS sg13g2_FILL8
XSTDFILL66_392 VDD VSS sg13g2_FILL8
XSTDFILL66_400 VDD VSS sg13g2_FILL8
XSTDFILL66_408 VDD VSS sg13g2_FILL8
XSTDFILL66_416 VDD VSS sg13g2_FILL8
XSTDFILL66_424 VDD VSS sg13g2_FILL8
XSTDFILL66_432 VDD VSS sg13g2_FILL8
XSTDFILL66_440 VDD VSS sg13g2_FILL8
XSTDFILL66_448 VDD VSS sg13g2_FILL8
XSTDFILL66_456 VDD VSS sg13g2_FILL8
XSTDFILL66_464 VDD VSS sg13g2_FILL8
XSTDFILL66_472 VDD VSS sg13g2_FILL8
XSTDFILL66_480 VDD VSS sg13g2_FILL8
XSTDFILL66_488 VDD VSS sg13g2_FILL8
XSTDFILL66_496 VDD VSS sg13g2_FILL8
XSTDFILL66_504 VDD VSS sg13g2_FILL8
XSTDFILL66_512 VDD VSS sg13g2_FILL8
XSTDFILL66_520 VDD VSS sg13g2_FILL8
XSTDFILL66_528 VDD VSS sg13g2_FILL8
XSTDFILL66_536 VDD VSS sg13g2_FILL8
XSTDFILL66_544 VDD VSS sg13g2_FILL8
XSTDFILL66_552 VDD VSS sg13g2_FILL8
XSTDFILL66_560 VDD VSS sg13g2_FILL8
XSTDFILL66_568 VDD VSS sg13g2_FILL8
XSTDFILL66_576 VDD VSS sg13g2_FILL8
XSTDFILL66_584 VDD VSS sg13g2_FILL8
XSTDFILL66_592 VDD VSS sg13g2_FILL8
XSTDFILL66_600 VDD VSS sg13g2_FILL8
XSTDFILL66_608 VDD VSS sg13g2_FILL8
XSTDFILL66_616 VDD VSS sg13g2_FILL8
XSTDFILL66_624 VDD VSS sg13g2_FILL8
XSTDFILL66_632 VDD VSS sg13g2_FILL8
XSTDFILL66_640 VDD VSS sg13g2_FILL8
XSTDFILL66_648 VDD VSS sg13g2_FILL8
XSTDFILL66_656 VDD VSS sg13g2_FILL8
XSTDFILL66_664 VDD VSS sg13g2_FILL8
XSTDFILL66_672 VDD VSS sg13g2_FILL8
XSTDFILL66_680 VDD VSS sg13g2_FILL8
XSTDFILL66_688 VDD VSS sg13g2_FILL8
XSTDFILL66_696 VDD VSS sg13g2_FILL8
XSTDFILL66_704 VDD VSS sg13g2_FILL8
XSTDFILL66_712 VDD VSS sg13g2_FILL8
XSTDFILL66_720 VDD VSS sg13g2_FILL8
XSTDFILL66_728 VDD VSS sg13g2_FILL8
XSTDFILL66_736 VDD VSS sg13g2_FILL8
XSTDFILL66_744 VDD VSS sg13g2_FILL8
XSTDFILL66_752 VDD VSS sg13g2_FILL8
XSTDFILL66_760 VDD VSS sg13g2_FILL8
XSTDFILL66_768 VDD VSS sg13g2_FILL8
XSTDFILL66_776 VDD VSS sg13g2_FILL8
XSTDFILL66_784 VDD VSS sg13g2_FILL8
XSTDFILL66_792 VDD VSS sg13g2_FILL8
XSTDFILL66_800 VDD VSS sg13g2_FILL8
XSTDFILL66_808 VDD VSS sg13g2_FILL8
XSTDFILL66_816 VDD VSS sg13g2_FILL8
XSTDFILL66_824 VDD VSS sg13g2_FILL8
XSTDFILL66_832 VDD VSS sg13g2_FILL8
XSTDFILL66_840 VDD VSS sg13g2_FILL8
XSTDFILL66_848 VDD VSS sg13g2_FILL8
XSTDFILL66_856 VDD VSS sg13g2_FILL8
XSTDFILL66_864 VDD VSS sg13g2_FILL8
XSTDFILL66_872 VDD VSS sg13g2_FILL8
XSTDFILL66_880 VDD VSS sg13g2_FILL8
XSTDFILL66_888 VDD VSS sg13g2_FILL8
XSTDFILL66_896 VDD VSS sg13g2_FILL8
XSTDFILL66_904 VDD VSS sg13g2_FILL8
XSTDFILL66_912 VDD VSS sg13g2_FILL8
XSTDFILL66_920 VDD VSS sg13g2_FILL8
XSTDFILL66_928 VDD VSS sg13g2_FILL8
XSTDFILL66_936 VDD VSS sg13g2_FILL8
XSTDFILL66_944 VDD VSS sg13g2_FILL8
XSTDFILL66_952 VDD VSS sg13g2_FILL8
XSTDFILL66_960 VDD VSS sg13g2_FILL8
XSTDFILL66_968 VDD VSS sg13g2_FILL8
XSTDFILL66_976 VDD VSS sg13g2_FILL8
XSTDFILL66_984 VDD VSS sg13g2_FILL8
XSTDFILL66_992 VDD VSS sg13g2_FILL8
XSTDFILL66_1000 VDD VSS sg13g2_FILL8
XSTDFILL66_1008 VDD VSS sg13g2_FILL8
XSTDFILL66_1016 VDD VSS sg13g2_FILL8
XSTDFILL66_1024 VDD VSS sg13g2_FILL8
XSTDFILL66_1032 VDD VSS sg13g2_FILL8
XSTDFILL66_1040 VDD VSS sg13g2_FILL8
XSTDFILL66_1048 VDD VSS sg13g2_FILL8
XSTDFILL66_1056 VDD VSS sg13g2_FILL8
XSTDFILL66_1064 VDD VSS sg13g2_FILL8
XSTDFILL66_1072 VDD VSS sg13g2_FILL8
XSTDFILL66_1080 VDD VSS sg13g2_FILL8
XSTDFILL66_1088 VDD VSS sg13g2_FILL8
XSTDFILL66_1096 VDD VSS sg13g2_FILL8
XSTDFILL66_1104 VDD VSS sg13g2_FILL8
XSTDFILL66_1112 VDD VSS sg13g2_FILL8
XSTDFILL66_1120 VDD VSS sg13g2_FILL8
XSTDFILL66_1128 VDD VSS sg13g2_FILL8
XSTDFILL66_1136 VDD VSS sg13g2_FILL8
XSTDFILL66_1144 VDD VSS sg13g2_FILL8
XSTDFILL66_1152 VDD VSS sg13g2_FILL8
XSTDFILL66_1160 VDD VSS sg13g2_FILL8
XSTDFILL66_1168 VDD VSS sg13g2_FILL8
XSTDFILL66_1176 VDD VSS sg13g2_FILL8
XSTDFILL66_1184 VDD VSS sg13g2_FILL8
XSTDFILL66_1192 VDD VSS sg13g2_FILL8
XSTDFILL66_1200 VDD VSS sg13g2_FILL8
XSTDFILL66_1208 VDD VSS sg13g2_FILL8
XSTDFILL66_1216 VDD VSS sg13g2_FILL8
XSTDFILL66_1224 VDD VSS sg13g2_FILL8
XSTDFILL66_1232 VDD VSS sg13g2_FILL8
XSTDFILL66_1240 VDD VSS sg13g2_FILL8
XSTDFILL66_1248 VDD VSS sg13g2_FILL8
XSTDFILL66_1256 VDD VSS sg13g2_FILL8
XSTDFILL66_1264 VDD VSS sg13g2_FILL8
XSTDFILL66_1272 VDD VSS sg13g2_FILL8
XSTDFILL66_1280 VDD VSS sg13g2_FILL8
XSTDFILL66_1288 VDD VSS sg13g2_FILL8
XSTDFILL66_1296 VDD VSS sg13g2_FILL8
XSTDFILL66_1304 VDD VSS sg13g2_FILL8
XSTDFILL66_1312 VDD VSS sg13g2_FILL8
XSTDFILL66_1320 VDD VSS sg13g2_FILL8
XSTDFILL66_1328 VDD VSS sg13g2_FILL8
XSTDFILL66_1336 VDD VSS sg13g2_FILL8
XSTDFILL66_1344 VDD VSS sg13g2_FILL8
XSTDFILL66_1352 VDD VSS sg13g2_FILL8
XSTDFILL66_1360 VDD VSS sg13g2_FILL8
XSTDFILL66_1368 VDD VSS sg13g2_FILL8
XSTDFILL66_1376 VDD VSS sg13g2_FILL8
XSTDFILL66_1384 VDD VSS sg13g2_FILL8
XSTDFILL66_1392 VDD VSS sg13g2_FILL8
XSTDFILL66_1400 VDD VSS sg13g2_FILL8
XSTDFILL66_1408 VDD VSS sg13g2_FILL8
XSTDFILL66_1416 VDD VSS sg13g2_FILL8
XSTDFILL66_1424 VDD VSS sg13g2_FILL8
XSTDFILL66_1432 VDD VSS sg13g2_FILL8
XSTDFILL66_1440 VDD VSS sg13g2_FILL8
XSTDFILL66_1448 VDD VSS sg13g2_FILL8
XSTDFILL66_1456 VDD VSS sg13g2_FILL8
XSTDFILL66_1464 VDD VSS sg13g2_FILL8
XSTDFILL66_1472 VDD VSS sg13g2_FILL8
XSTDFILL66_1480 VDD VSS sg13g2_FILL8
XSTDFILL66_1488 VDD VSS sg13g2_FILL8
XSTDFILL66_1496 VDD VSS sg13g2_FILL8
XSTDFILL66_1504 VDD VSS sg13g2_FILL8
XSTDFILL66_1512 VDD VSS sg13g2_FILL8
XSTDFILL66_1520 VDD VSS sg13g2_FILL8
XSTDFILL66_1528 VDD VSS sg13g2_FILL8
XSTDFILL66_1536 VDD VSS sg13g2_FILL8
XSTDFILL66_1544 VDD VSS sg13g2_FILL8
XSTDFILL66_1552 VDD VSS sg13g2_FILL8
XSTDFILL66_1560 VDD VSS sg13g2_FILL8
XSTDFILL66_1568 VDD VSS sg13g2_FILL8
XSTDFILL66_1576 VDD VSS sg13g2_FILL8
XSTDFILL66_1584 VDD VSS sg13g2_FILL8
XSTDFILL66_1592 VDD VSS sg13g2_FILL8
XSTDFILL66_1600 VDD VSS sg13g2_FILL8
XSTDFILL66_1608 VDD VSS sg13g2_FILL8
XSTDFILL66_1616 VDD VSS sg13g2_FILL8
XSTDFILL66_1624 VDD VSS sg13g2_FILL8
XSTDFILL66_1632 VDD VSS sg13g2_FILL8
XSTDFILL66_1640 VDD VSS sg13g2_FILL8
XSTDFILL66_1648 VDD VSS sg13g2_FILL8
XSTDFILL66_1656 VDD VSS sg13g2_FILL8
XSTDFILL66_1664 VDD VSS sg13g2_FILL8
XSTDFILL66_1672 VDD VSS sg13g2_FILL8
XSTDFILL66_1680 VDD VSS sg13g2_FILL8
XSTDFILL66_1688 VDD VSS sg13g2_FILL8
XSTDFILL66_1696 VDD VSS sg13g2_FILL8
XSTDFILL66_1704 VDD VSS sg13g2_FILL8
XSTDFILL66_1712 VDD VSS sg13g2_FILL8
XSTDFILL66_1720 VDD VSS sg13g2_FILL8
XSTDFILL66_1728 VDD VSS sg13g2_FILL8
XSTDFILL66_1736 VDD VSS sg13g2_FILL8
XSTDFILL66_1744 VDD VSS sg13g2_FILL8
XSTDFILL66_1752 VDD VSS sg13g2_FILL8
XSTDFILL66_1760 VDD VSS sg13g2_FILL8
XSTDFILL66_1768 VDD VSS sg13g2_FILL8
XSTDFILL66_1776 VDD VSS sg13g2_FILL8
XSTDFILL66_1784 VDD VSS sg13g2_FILL8
XSTDFILL66_1792 VDD VSS sg13g2_FILL8
XSTDFILL66_1800 VDD VSS sg13g2_FILL8
XSTDFILL66_1808 VDD VSS sg13g2_FILL8
XSTDFILL66_1816 VDD VSS sg13g2_FILL8
XSTDFILL66_1824 VDD VSS sg13g2_FILL8
XSTDFILL66_1832 VDD VSS sg13g2_FILL8
XSTDFILL66_1840 VDD VSS sg13g2_FILL8
XSTDFILL66_1848 VDD VSS sg13g2_FILL8
XSTDFILL66_1856 VDD VSS sg13g2_FILL8
XSTDFILL66_1864 VDD VSS sg13g2_FILL8
XSTDFILL66_1872 VDD VSS sg13g2_FILL8
XSTDFILL66_1880 VDD VSS sg13g2_FILL8
XSTDFILL66_1888 VDD VSS sg13g2_FILL8
XSTDFILL66_1896 VDD VSS sg13g2_FILL8
XSTDFILL66_1904 VDD VSS sg13g2_FILL8
XSTDFILL66_1912 VDD VSS sg13g2_FILL8
XSTDFILL66_1920 VDD VSS sg13g2_FILL8
XSTDFILL66_1928 VDD VSS sg13g2_FILL8
XSTDFILL66_1936 VDD VSS sg13g2_FILL8
XSTDFILL66_1944 VDD VSS sg13g2_FILL8
XSTDFILL66_1952 VDD VSS sg13g2_FILL8
XSTDFILL66_1960 VDD VSS sg13g2_FILL8
XSTDFILL66_1968 VDD VSS sg13g2_FILL8
XSTDFILL66_1976 VDD VSS sg13g2_FILL8
XSTDFILL66_1984 VDD VSS sg13g2_FILL8
XSTDFILL66_1992 VDD VSS sg13g2_FILL8
XSTDFILL66_2000 VDD VSS sg13g2_FILL8
XSTDFILL66_2008 VDD VSS sg13g2_FILL8
XSTDFILL66_2016 VDD VSS sg13g2_FILL8
XSTDFILL66_2024 VDD VSS sg13g2_FILL8
XSTDFILL66_2032 VDD VSS sg13g2_FILL8
XSTDFILL66_2040 VDD VSS sg13g2_FILL8
XSTDFILL66_2048 VDD VSS sg13g2_FILL8
XSTDFILL66_2056 VDD VSS sg13g2_FILL8
XSTDFILL66_2064 VDD VSS sg13g2_FILL8
XSTDFILL66_2072 VDD VSS sg13g2_FILL8
XSTDFILL66_2080 VDD VSS sg13g2_FILL8
XSTDFILL66_2088 VDD VSS sg13g2_FILL8
XSTDFILL66_2096 VDD VSS sg13g2_FILL8
XSTDFILL66_2104 VDD VSS sg13g2_FILL8
XSTDFILL66_2112 VDD VSS sg13g2_FILL8
XSTDFILL66_2120 VDD VSS sg13g2_FILL8
XSTDFILL66_2128 VDD VSS sg13g2_FILL8
XSTDFILL66_2136 VDD VSS sg13g2_FILL8
XSTDFILL66_2144 VDD VSS sg13g2_FILL8
XSTDFILL66_2152 VDD VSS sg13g2_FILL2
XSTDFILL67_0 VDD VSS sg13g2_FILL8
XSTDFILL67_8 VDD VSS sg13g2_FILL8
XSTDFILL67_16 VDD VSS sg13g2_FILL8
XSTDFILL67_24 VDD VSS sg13g2_FILL8
XSTDFILL67_32 VDD VSS sg13g2_FILL8
XSTDFILL67_40 VDD VSS sg13g2_FILL8
XSTDFILL67_48 VDD VSS sg13g2_FILL8
XSTDFILL67_56 VDD VSS sg13g2_FILL8
XSTDFILL67_64 VDD VSS sg13g2_FILL8
XSTDFILL67_72 VDD VSS sg13g2_FILL8
XSTDFILL67_80 VDD VSS sg13g2_FILL8
XSTDFILL67_88 VDD VSS sg13g2_FILL8
XSTDFILL67_96 VDD VSS sg13g2_FILL8
XSTDFILL67_104 VDD VSS sg13g2_FILL8
XSTDFILL67_112 VDD VSS sg13g2_FILL8
XSTDFILL67_120 VDD VSS sg13g2_FILL8
XSTDFILL67_128 VDD VSS sg13g2_FILL8
XSTDFILL67_136 VDD VSS sg13g2_FILL8
XSTDFILL67_144 VDD VSS sg13g2_FILL8
XSTDFILL67_152 VDD VSS sg13g2_FILL8
XSTDFILL67_160 VDD VSS sg13g2_FILL8
XSTDFILL67_168 VDD VSS sg13g2_FILL8
XSTDFILL67_176 VDD VSS sg13g2_FILL8
XSTDFILL67_184 VDD VSS sg13g2_FILL8
XSTDFILL67_192 VDD VSS sg13g2_FILL8
XSTDFILL67_200 VDD VSS sg13g2_FILL8
XSTDFILL67_208 VDD VSS sg13g2_FILL8
XSTDFILL67_216 VDD VSS sg13g2_FILL8
XSTDFILL67_224 VDD VSS sg13g2_FILL8
XSTDFILL67_232 VDD VSS sg13g2_FILL8
XSTDFILL67_240 VDD VSS sg13g2_FILL8
XSTDFILL67_248 VDD VSS sg13g2_FILL8
XSTDFILL67_256 VDD VSS sg13g2_FILL8
XSTDFILL67_264 VDD VSS sg13g2_FILL8
XSTDFILL67_272 VDD VSS sg13g2_FILL8
XSTDFILL67_280 VDD VSS sg13g2_FILL8
XSTDFILL67_288 VDD VSS sg13g2_FILL8
XSTDFILL67_296 VDD VSS sg13g2_FILL8
XSTDFILL67_304 VDD VSS sg13g2_FILL8
XSTDFILL67_312 VDD VSS sg13g2_FILL8
XSTDFILL67_320 VDD VSS sg13g2_FILL8
XSTDFILL67_328 VDD VSS sg13g2_FILL8
XSTDFILL67_336 VDD VSS sg13g2_FILL8
XSTDFILL67_344 VDD VSS sg13g2_FILL8
XSTDFILL67_352 VDD VSS sg13g2_FILL8
XSTDFILL67_360 VDD VSS sg13g2_FILL8
XSTDFILL67_368 VDD VSS sg13g2_FILL8
XSTDFILL67_376 VDD VSS sg13g2_FILL8
XSTDFILL67_384 VDD VSS sg13g2_FILL8
XSTDFILL67_392 VDD VSS sg13g2_FILL8
XSTDFILL67_400 VDD VSS sg13g2_FILL8
XSTDFILL67_408 VDD VSS sg13g2_FILL8
XSTDFILL67_416 VDD VSS sg13g2_FILL8
XSTDFILL67_424 VDD VSS sg13g2_FILL8
XSTDFILL67_432 VDD VSS sg13g2_FILL8
XSTDFILL67_440 VDD VSS sg13g2_FILL8
XSTDFILL67_448 VDD VSS sg13g2_FILL8
XSTDFILL67_456 VDD VSS sg13g2_FILL8
XSTDFILL67_464 VDD VSS sg13g2_FILL8
XSTDFILL67_472 VDD VSS sg13g2_FILL8
XSTDFILL67_480 VDD VSS sg13g2_FILL8
XSTDFILL67_488 VDD VSS sg13g2_FILL8
XSTDFILL67_496 VDD VSS sg13g2_FILL8
XSTDFILL67_504 VDD VSS sg13g2_FILL8
XSTDFILL67_512 VDD VSS sg13g2_FILL8
XSTDFILL67_520 VDD VSS sg13g2_FILL8
XSTDFILL67_528 VDD VSS sg13g2_FILL8
XSTDFILL67_536 VDD VSS sg13g2_FILL8
XSTDFILL67_544 VDD VSS sg13g2_FILL8
XSTDFILL67_552 VDD VSS sg13g2_FILL8
XSTDFILL67_560 VDD VSS sg13g2_FILL8
XSTDFILL67_568 VDD VSS sg13g2_FILL8
XSTDFILL67_576 VDD VSS sg13g2_FILL8
XSTDFILL67_584 VDD VSS sg13g2_FILL8
XSTDFILL67_592 VDD VSS sg13g2_FILL8
XSTDFILL67_600 VDD VSS sg13g2_FILL8
XSTDFILL67_608 VDD VSS sg13g2_FILL8
XSTDFILL67_616 VDD VSS sg13g2_FILL8
XSTDFILL67_624 VDD VSS sg13g2_FILL8
XSTDFILL67_632 VDD VSS sg13g2_FILL8
XSTDFILL67_640 VDD VSS sg13g2_FILL8
XSTDFILL67_648 VDD VSS sg13g2_FILL8
XSTDFILL67_656 VDD VSS sg13g2_FILL8
XSTDFILL67_664 VDD VSS sg13g2_FILL8
XSTDFILL67_672 VDD VSS sg13g2_FILL8
XSTDFILL67_680 VDD VSS sg13g2_FILL8
XSTDFILL67_688 VDD VSS sg13g2_FILL8
XSTDFILL67_696 VDD VSS sg13g2_FILL8
XSTDFILL67_704 VDD VSS sg13g2_FILL8
XSTDFILL67_712 VDD VSS sg13g2_FILL8
XSTDFILL67_720 VDD VSS sg13g2_FILL8
XSTDFILL67_728 VDD VSS sg13g2_FILL8
XSTDFILL67_736 VDD VSS sg13g2_FILL8
XSTDFILL67_744 VDD VSS sg13g2_FILL8
XSTDFILL67_752 VDD VSS sg13g2_FILL8
XSTDFILL67_760 VDD VSS sg13g2_FILL8
XSTDFILL67_768 VDD VSS sg13g2_FILL8
XSTDFILL67_776 VDD VSS sg13g2_FILL8
XSTDFILL67_784 VDD VSS sg13g2_FILL8
XSTDFILL67_792 VDD VSS sg13g2_FILL8
XSTDFILL67_800 VDD VSS sg13g2_FILL8
XSTDFILL67_808 VDD VSS sg13g2_FILL8
XSTDFILL67_816 VDD VSS sg13g2_FILL8
XSTDFILL67_824 VDD VSS sg13g2_FILL8
XSTDFILL67_832 VDD VSS sg13g2_FILL8
XSTDFILL67_840 VDD VSS sg13g2_FILL8
XSTDFILL67_848 VDD VSS sg13g2_FILL8
XSTDFILL67_856 VDD VSS sg13g2_FILL8
XSTDFILL67_864 VDD VSS sg13g2_FILL8
XSTDFILL67_872 VDD VSS sg13g2_FILL8
XSTDFILL67_880 VDD VSS sg13g2_FILL8
XSTDFILL67_888 VDD VSS sg13g2_FILL8
XSTDFILL67_896 VDD VSS sg13g2_FILL8
XSTDFILL67_904 VDD VSS sg13g2_FILL8
XSTDFILL67_912 VDD VSS sg13g2_FILL8
XSTDFILL67_920 VDD VSS sg13g2_FILL8
XSTDFILL67_928 VDD VSS sg13g2_FILL8
XSTDFILL67_936 VDD VSS sg13g2_FILL8
XSTDFILL67_944 VDD VSS sg13g2_FILL8
XSTDFILL67_952 VDD VSS sg13g2_FILL8
XSTDFILL67_960 VDD VSS sg13g2_FILL8
XSTDFILL67_968 VDD VSS sg13g2_FILL8
XSTDFILL67_976 VDD VSS sg13g2_FILL8
XSTDFILL67_984 VDD VSS sg13g2_FILL8
XSTDFILL67_992 VDD VSS sg13g2_FILL8
XSTDFILL67_1000 VDD VSS sg13g2_FILL8
XSTDFILL67_1008 VDD VSS sg13g2_FILL8
XSTDFILL67_1016 VDD VSS sg13g2_FILL8
XSTDFILL67_1024 VDD VSS sg13g2_FILL8
XSTDFILL67_1032 VDD VSS sg13g2_FILL8
XSTDFILL67_1040 VDD VSS sg13g2_FILL8
XSTDFILL67_1048 VDD VSS sg13g2_FILL8
XSTDFILL67_1056 VDD VSS sg13g2_FILL8
XSTDFILL67_1064 VDD VSS sg13g2_FILL8
XSTDFILL67_1072 VDD VSS sg13g2_FILL8
XSTDFILL67_1080 VDD VSS sg13g2_FILL8
XSTDFILL67_1088 VDD VSS sg13g2_FILL8
XSTDFILL67_1096 VDD VSS sg13g2_FILL8
XSTDFILL67_1104 VDD VSS sg13g2_FILL8
XSTDFILL67_1112 VDD VSS sg13g2_FILL8
XSTDFILL67_1120 VDD VSS sg13g2_FILL8
XSTDFILL67_1128 VDD VSS sg13g2_FILL8
XSTDFILL67_1136 VDD VSS sg13g2_FILL8
XSTDFILL67_1144 VDD VSS sg13g2_FILL8
XSTDFILL67_1152 VDD VSS sg13g2_FILL8
XSTDFILL67_1160 VDD VSS sg13g2_FILL8
XSTDFILL67_1168 VDD VSS sg13g2_FILL8
XSTDFILL67_1176 VDD VSS sg13g2_FILL8
XSTDFILL67_1184 VDD VSS sg13g2_FILL8
XSTDFILL67_1192 VDD VSS sg13g2_FILL8
XSTDFILL67_1200 VDD VSS sg13g2_FILL8
XSTDFILL67_1208 VDD VSS sg13g2_FILL8
XSTDFILL67_1216 VDD VSS sg13g2_FILL8
XSTDFILL67_1224 VDD VSS sg13g2_FILL8
XSTDFILL67_1232 VDD VSS sg13g2_FILL8
XSTDFILL67_1240 VDD VSS sg13g2_FILL8
XSTDFILL67_1248 VDD VSS sg13g2_FILL8
XSTDFILL67_1256 VDD VSS sg13g2_FILL8
XSTDFILL67_1264 VDD VSS sg13g2_FILL8
XSTDFILL67_1272 VDD VSS sg13g2_FILL8
XSTDFILL67_1280 VDD VSS sg13g2_FILL8
XSTDFILL67_1288 VDD VSS sg13g2_FILL8
XSTDFILL67_1296 VDD VSS sg13g2_FILL8
XSTDFILL67_1304 VDD VSS sg13g2_FILL8
XSTDFILL67_1312 VDD VSS sg13g2_FILL8
XSTDFILL67_1320 VDD VSS sg13g2_FILL8
XSTDFILL67_1328 VDD VSS sg13g2_FILL8
XSTDFILL67_1336 VDD VSS sg13g2_FILL8
XSTDFILL67_1344 VDD VSS sg13g2_FILL8
XSTDFILL67_1352 VDD VSS sg13g2_FILL8
XSTDFILL67_1360 VDD VSS sg13g2_FILL8
XSTDFILL67_1368 VDD VSS sg13g2_FILL8
XSTDFILL67_1376 VDD VSS sg13g2_FILL8
XSTDFILL67_1384 VDD VSS sg13g2_FILL8
XSTDFILL67_1392 VDD VSS sg13g2_FILL8
XSTDFILL67_1400 VDD VSS sg13g2_FILL8
XSTDFILL67_1408 VDD VSS sg13g2_FILL8
XSTDFILL67_1416 VDD VSS sg13g2_FILL8
XSTDFILL67_1424 VDD VSS sg13g2_FILL8
XSTDFILL67_1432 VDD VSS sg13g2_FILL8
XSTDFILL67_1440 VDD VSS sg13g2_FILL8
XSTDFILL67_1448 VDD VSS sg13g2_FILL8
XSTDFILL67_1456 VDD VSS sg13g2_FILL8
XSTDFILL67_1464 VDD VSS sg13g2_FILL8
XSTDFILL67_1472 VDD VSS sg13g2_FILL8
XSTDFILL67_1480 VDD VSS sg13g2_FILL8
XSTDFILL67_1488 VDD VSS sg13g2_FILL8
XSTDFILL67_1496 VDD VSS sg13g2_FILL8
XSTDFILL67_1504 VDD VSS sg13g2_FILL8
XSTDFILL67_1512 VDD VSS sg13g2_FILL8
XSTDFILL67_1520 VDD VSS sg13g2_FILL8
XSTDFILL67_1528 VDD VSS sg13g2_FILL8
XSTDFILL67_1536 VDD VSS sg13g2_FILL8
XSTDFILL67_1544 VDD VSS sg13g2_FILL8
XSTDFILL67_1552 VDD VSS sg13g2_FILL8
XSTDFILL67_1560 VDD VSS sg13g2_FILL8
XSTDFILL67_1568 VDD VSS sg13g2_FILL8
XSTDFILL67_1576 VDD VSS sg13g2_FILL8
XSTDFILL67_1584 VDD VSS sg13g2_FILL8
XSTDFILL67_1592 VDD VSS sg13g2_FILL8
XSTDFILL67_1600 VDD VSS sg13g2_FILL8
XSTDFILL67_1608 VDD VSS sg13g2_FILL8
XSTDFILL67_1616 VDD VSS sg13g2_FILL8
XSTDFILL67_1624 VDD VSS sg13g2_FILL8
XSTDFILL67_1632 VDD VSS sg13g2_FILL8
XSTDFILL67_1640 VDD VSS sg13g2_FILL8
XSTDFILL67_1648 VDD VSS sg13g2_FILL8
XSTDFILL67_1656 VDD VSS sg13g2_FILL8
XSTDFILL67_1664 VDD VSS sg13g2_FILL8
XSTDFILL67_1672 VDD VSS sg13g2_FILL8
XSTDFILL67_1680 VDD VSS sg13g2_FILL8
XSTDFILL67_1688 VDD VSS sg13g2_FILL8
XSTDFILL67_1696 VDD VSS sg13g2_FILL8
XSTDFILL67_1704 VDD VSS sg13g2_FILL8
XSTDFILL67_1712 VDD VSS sg13g2_FILL8
XSTDFILL67_1720 VDD VSS sg13g2_FILL8
XSTDFILL67_1728 VDD VSS sg13g2_FILL8
XSTDFILL67_1736 VDD VSS sg13g2_FILL8
XSTDFILL67_1744 VDD VSS sg13g2_FILL8
XSTDFILL67_1752 VDD VSS sg13g2_FILL8
XSTDFILL67_1760 VDD VSS sg13g2_FILL8
XSTDFILL67_1768 VDD VSS sg13g2_FILL8
XSTDFILL67_1776 VDD VSS sg13g2_FILL8
XSTDFILL67_1784 VDD VSS sg13g2_FILL8
XSTDFILL67_1792 VDD VSS sg13g2_FILL8
XSTDFILL67_1800 VDD VSS sg13g2_FILL8
XSTDFILL67_1808 VDD VSS sg13g2_FILL8
XSTDFILL67_1816 VDD VSS sg13g2_FILL8
XSTDFILL67_1824 VDD VSS sg13g2_FILL8
XSTDFILL67_1832 VDD VSS sg13g2_FILL8
XSTDFILL67_1840 VDD VSS sg13g2_FILL8
XSTDFILL67_1848 VDD VSS sg13g2_FILL8
XSTDFILL67_1856 VDD VSS sg13g2_FILL8
XSTDFILL67_1864 VDD VSS sg13g2_FILL8
XSTDFILL67_1872 VDD VSS sg13g2_FILL8
XSTDFILL67_1880 VDD VSS sg13g2_FILL8
XSTDFILL67_1888 VDD VSS sg13g2_FILL8
XSTDFILL67_1896 VDD VSS sg13g2_FILL8
XSTDFILL67_1904 VDD VSS sg13g2_FILL8
XSTDFILL67_1912 VDD VSS sg13g2_FILL8
XSTDFILL67_1920 VDD VSS sg13g2_FILL8
XSTDFILL67_1928 VDD VSS sg13g2_FILL8
XSTDFILL67_1936 VDD VSS sg13g2_FILL8
XSTDFILL67_1944 VDD VSS sg13g2_FILL8
XSTDFILL67_1952 VDD VSS sg13g2_FILL8
XSTDFILL67_1960 VDD VSS sg13g2_FILL8
XSTDFILL67_1968 VDD VSS sg13g2_FILL8
XSTDFILL67_1976 VDD VSS sg13g2_FILL8
XSTDFILL67_1984 VDD VSS sg13g2_FILL8
XSTDFILL67_1992 VDD VSS sg13g2_FILL8
XSTDFILL67_2000 VDD VSS sg13g2_FILL8
XSTDFILL67_2008 VDD VSS sg13g2_FILL8
XSTDFILL67_2016 VDD VSS sg13g2_FILL8
XSTDFILL67_2024 VDD VSS sg13g2_FILL8
XSTDFILL67_2032 VDD VSS sg13g2_FILL8
XSTDFILL67_2040 VDD VSS sg13g2_FILL8
XSTDFILL67_2048 VDD VSS sg13g2_FILL8
XSTDFILL67_2056 VDD VSS sg13g2_FILL8
XSTDFILL67_2064 VDD VSS sg13g2_FILL8
XSTDFILL67_2072 VDD VSS sg13g2_FILL8
XSTDFILL67_2080 VDD VSS sg13g2_FILL8
XSTDFILL67_2088 VDD VSS sg13g2_FILL8
XSTDFILL67_2096 VDD VSS sg13g2_FILL8
XSTDFILL67_2104 VDD VSS sg13g2_FILL8
XSTDFILL67_2112 VDD VSS sg13g2_FILL8
XSTDFILL67_2120 VDD VSS sg13g2_FILL8
XSTDFILL67_2128 VDD VSS sg13g2_FILL8
XSTDFILL67_2136 VDD VSS sg13g2_FILL8
XSTDFILL67_2144 VDD VSS sg13g2_FILL8
XSTDFILL67_2152 VDD VSS sg13g2_FILL2
XSTDFILL68_0 VDD VSS sg13g2_FILL8
XSTDFILL68_8 VDD VSS sg13g2_FILL8
XSTDFILL68_16 VDD VSS sg13g2_FILL8
XSTDFILL68_24 VDD VSS sg13g2_FILL8
XSTDFILL68_32 VDD VSS sg13g2_FILL8
XSTDFILL68_40 VDD VSS sg13g2_FILL8
XSTDFILL68_48 VDD VSS sg13g2_FILL8
XSTDFILL68_56 VDD VSS sg13g2_FILL8
XSTDFILL68_64 VDD VSS sg13g2_FILL8
XSTDFILL68_72 VDD VSS sg13g2_FILL8
XSTDFILL68_80 VDD VSS sg13g2_FILL8
XSTDFILL68_88 VDD VSS sg13g2_FILL8
XSTDFILL68_96 VDD VSS sg13g2_FILL8
XSTDFILL68_104 VDD VSS sg13g2_FILL8
XSTDFILL68_112 VDD VSS sg13g2_FILL8
XSTDFILL68_120 VDD VSS sg13g2_FILL8
XSTDFILL68_128 VDD VSS sg13g2_FILL8
XSTDFILL68_136 VDD VSS sg13g2_FILL8
XSTDFILL68_144 VDD VSS sg13g2_FILL8
XSTDFILL68_152 VDD VSS sg13g2_FILL8
XSTDFILL68_160 VDD VSS sg13g2_FILL8
XSTDFILL68_168 VDD VSS sg13g2_FILL8
XSTDFILL68_176 VDD VSS sg13g2_FILL8
XSTDFILL68_184 VDD VSS sg13g2_FILL8
XSTDFILL68_192 VDD VSS sg13g2_FILL8
XSTDFILL68_200 VDD VSS sg13g2_FILL8
XSTDFILL68_208 VDD VSS sg13g2_FILL8
XSTDFILL68_216 VDD VSS sg13g2_FILL8
XSTDFILL68_224 VDD VSS sg13g2_FILL8
XSTDFILL68_232 VDD VSS sg13g2_FILL8
XSTDFILL68_240 VDD VSS sg13g2_FILL8
XSTDFILL68_248 VDD VSS sg13g2_FILL8
XSTDFILL68_256 VDD VSS sg13g2_FILL8
XSTDFILL68_264 VDD VSS sg13g2_FILL8
XSTDFILL68_272 VDD VSS sg13g2_FILL8
XSTDFILL68_280 VDD VSS sg13g2_FILL8
XSTDFILL68_288 VDD VSS sg13g2_FILL8
XSTDFILL68_296 VDD VSS sg13g2_FILL8
XSTDFILL68_304 VDD VSS sg13g2_FILL8
XSTDFILL68_312 VDD VSS sg13g2_FILL8
XSTDFILL68_320 VDD VSS sg13g2_FILL8
XSTDFILL68_328 VDD VSS sg13g2_FILL8
XSTDFILL68_336 VDD VSS sg13g2_FILL8
XSTDFILL68_344 VDD VSS sg13g2_FILL8
XSTDFILL68_352 VDD VSS sg13g2_FILL8
XSTDFILL68_360 VDD VSS sg13g2_FILL8
XSTDFILL68_368 VDD VSS sg13g2_FILL8
XSTDFILL68_376 VDD VSS sg13g2_FILL8
XSTDFILL68_384 VDD VSS sg13g2_FILL8
XSTDFILL68_392 VDD VSS sg13g2_FILL8
XSTDFILL68_400 VDD VSS sg13g2_FILL8
XSTDFILL68_408 VDD VSS sg13g2_FILL8
XSTDFILL68_416 VDD VSS sg13g2_FILL8
XSTDFILL68_424 VDD VSS sg13g2_FILL8
XSTDFILL68_432 VDD VSS sg13g2_FILL8
XSTDFILL68_440 VDD VSS sg13g2_FILL8
XSTDFILL68_448 VDD VSS sg13g2_FILL8
XSTDFILL68_456 VDD VSS sg13g2_FILL8
XSTDFILL68_464 VDD VSS sg13g2_FILL8
XSTDFILL68_472 VDD VSS sg13g2_FILL8
XSTDFILL68_480 VDD VSS sg13g2_FILL8
XSTDFILL68_488 VDD VSS sg13g2_FILL8
XSTDFILL68_496 VDD VSS sg13g2_FILL8
XSTDFILL68_504 VDD VSS sg13g2_FILL8
XSTDFILL68_512 VDD VSS sg13g2_FILL8
XSTDFILL68_520 VDD VSS sg13g2_FILL8
XSTDFILL68_528 VDD VSS sg13g2_FILL8
XSTDFILL68_536 VDD VSS sg13g2_FILL8
XSTDFILL68_544 VDD VSS sg13g2_FILL8
XSTDFILL68_552 VDD VSS sg13g2_FILL8
XSTDFILL68_560 VDD VSS sg13g2_FILL8
XSTDFILL68_568 VDD VSS sg13g2_FILL8
XSTDFILL68_576 VDD VSS sg13g2_FILL8
XSTDFILL68_584 VDD VSS sg13g2_FILL8
XSTDFILL68_592 VDD VSS sg13g2_FILL8
XSTDFILL68_600 VDD VSS sg13g2_FILL8
XSTDFILL68_608 VDD VSS sg13g2_FILL8
XSTDFILL68_616 VDD VSS sg13g2_FILL8
XSTDFILL68_624 VDD VSS sg13g2_FILL8
XSTDFILL68_632 VDD VSS sg13g2_FILL8
XSTDFILL68_640 VDD VSS sg13g2_FILL8
XSTDFILL68_648 VDD VSS sg13g2_FILL8
XSTDFILL68_656 VDD VSS sg13g2_FILL8
XSTDFILL68_664 VDD VSS sg13g2_FILL8
XSTDFILL68_672 VDD VSS sg13g2_FILL8
XSTDFILL68_680 VDD VSS sg13g2_FILL8
XSTDFILL68_688 VDD VSS sg13g2_FILL8
XSTDFILL68_696 VDD VSS sg13g2_FILL8
XSTDFILL68_704 VDD VSS sg13g2_FILL8
XSTDFILL68_712 VDD VSS sg13g2_FILL8
XSTDFILL68_720 VDD VSS sg13g2_FILL8
XSTDFILL68_728 VDD VSS sg13g2_FILL8
XSTDFILL68_736 VDD VSS sg13g2_FILL8
XSTDFILL68_744 VDD VSS sg13g2_FILL8
XSTDFILL68_752 VDD VSS sg13g2_FILL8
XSTDFILL68_760 VDD VSS sg13g2_FILL8
XSTDFILL68_768 VDD VSS sg13g2_FILL8
XSTDFILL68_776 VDD VSS sg13g2_FILL8
XSTDFILL68_784 VDD VSS sg13g2_FILL8
XSTDFILL68_792 VDD VSS sg13g2_FILL8
XSTDFILL68_800 VDD VSS sg13g2_FILL8
XSTDFILL68_808 VDD VSS sg13g2_FILL8
XSTDFILL68_816 VDD VSS sg13g2_FILL8
XSTDFILL68_824 VDD VSS sg13g2_FILL8
XSTDFILL68_832 VDD VSS sg13g2_FILL8
XSTDFILL68_840 VDD VSS sg13g2_FILL8
XSTDFILL68_848 VDD VSS sg13g2_FILL8
XSTDFILL68_856 VDD VSS sg13g2_FILL8
XSTDFILL68_864 VDD VSS sg13g2_FILL8
XSTDFILL68_872 VDD VSS sg13g2_FILL8
XSTDFILL68_880 VDD VSS sg13g2_FILL8
XSTDFILL68_888 VDD VSS sg13g2_FILL8
XSTDFILL68_896 VDD VSS sg13g2_FILL8
XSTDFILL68_904 VDD VSS sg13g2_FILL8
XSTDFILL68_912 VDD VSS sg13g2_FILL8
XSTDFILL68_920 VDD VSS sg13g2_FILL8
XSTDFILL68_928 VDD VSS sg13g2_FILL8
XSTDFILL68_936 VDD VSS sg13g2_FILL8
XSTDFILL68_944 VDD VSS sg13g2_FILL8
XSTDFILL68_952 VDD VSS sg13g2_FILL8
XSTDFILL68_960 VDD VSS sg13g2_FILL8
XSTDFILL68_968 VDD VSS sg13g2_FILL8
XSTDFILL68_976 VDD VSS sg13g2_FILL8
XSTDFILL68_984 VDD VSS sg13g2_FILL8
XSTDFILL68_992 VDD VSS sg13g2_FILL8
XSTDFILL68_1000 VDD VSS sg13g2_FILL8
XSTDFILL68_1008 VDD VSS sg13g2_FILL8
XSTDFILL68_1016 VDD VSS sg13g2_FILL8
XSTDFILL68_1024 VDD VSS sg13g2_FILL8
XSTDFILL68_1032 VDD VSS sg13g2_FILL8
XSTDFILL68_1040 VDD VSS sg13g2_FILL8
XSTDFILL68_1048 VDD VSS sg13g2_FILL8
XSTDFILL68_1056 VDD VSS sg13g2_FILL8
XSTDFILL68_1064 VDD VSS sg13g2_FILL8
XSTDFILL68_1072 VDD VSS sg13g2_FILL8
XSTDFILL68_1080 VDD VSS sg13g2_FILL8
XSTDFILL68_1088 VDD VSS sg13g2_FILL8
XSTDFILL68_1096 VDD VSS sg13g2_FILL8
XSTDFILL68_1104 VDD VSS sg13g2_FILL8
XSTDFILL68_1112 VDD VSS sg13g2_FILL8
XSTDFILL68_1120 VDD VSS sg13g2_FILL8
XSTDFILL68_1128 VDD VSS sg13g2_FILL8
XSTDFILL68_1136 VDD VSS sg13g2_FILL8
XSTDFILL68_1144 VDD VSS sg13g2_FILL8
XSTDFILL68_1152 VDD VSS sg13g2_FILL8
XSTDFILL68_1160 VDD VSS sg13g2_FILL8
XSTDFILL68_1168 VDD VSS sg13g2_FILL8
XSTDFILL68_1176 VDD VSS sg13g2_FILL8
XSTDFILL68_1184 VDD VSS sg13g2_FILL8
XSTDFILL68_1192 VDD VSS sg13g2_FILL8
XSTDFILL68_1200 VDD VSS sg13g2_FILL8
XSTDFILL68_1208 VDD VSS sg13g2_FILL8
XSTDFILL68_1216 VDD VSS sg13g2_FILL8
XSTDFILL68_1224 VDD VSS sg13g2_FILL8
XSTDFILL68_1232 VDD VSS sg13g2_FILL8
XSTDFILL68_1240 VDD VSS sg13g2_FILL8
XSTDFILL68_1248 VDD VSS sg13g2_FILL8
XSTDFILL68_1256 VDD VSS sg13g2_FILL8
XSTDFILL68_1264 VDD VSS sg13g2_FILL8
XSTDFILL68_1272 VDD VSS sg13g2_FILL8
XSTDFILL68_1280 VDD VSS sg13g2_FILL8
XSTDFILL68_1288 VDD VSS sg13g2_FILL8
XSTDFILL68_1296 VDD VSS sg13g2_FILL8
XSTDFILL68_1304 VDD VSS sg13g2_FILL8
XSTDFILL68_1312 VDD VSS sg13g2_FILL8
XSTDFILL68_1320 VDD VSS sg13g2_FILL8
XSTDFILL68_1328 VDD VSS sg13g2_FILL8
XSTDFILL68_1336 VDD VSS sg13g2_FILL8
XSTDFILL68_1344 VDD VSS sg13g2_FILL8
XSTDFILL68_1352 VDD VSS sg13g2_FILL8
XSTDFILL68_1360 VDD VSS sg13g2_FILL8
XSTDFILL68_1368 VDD VSS sg13g2_FILL8
XSTDFILL68_1376 VDD VSS sg13g2_FILL8
XSTDFILL68_1384 VDD VSS sg13g2_FILL8
XSTDFILL68_1392 VDD VSS sg13g2_FILL8
XSTDFILL68_1400 VDD VSS sg13g2_FILL8
XSTDFILL68_1408 VDD VSS sg13g2_FILL8
XSTDFILL68_1416 VDD VSS sg13g2_FILL8
XSTDFILL68_1424 VDD VSS sg13g2_FILL8
XSTDFILL68_1432 VDD VSS sg13g2_FILL8
XSTDFILL68_1440 VDD VSS sg13g2_FILL8
XSTDFILL68_1448 VDD VSS sg13g2_FILL8
XSTDFILL68_1456 VDD VSS sg13g2_FILL8
XSTDFILL68_1464 VDD VSS sg13g2_FILL8
XSTDFILL68_1472 VDD VSS sg13g2_FILL8
XSTDFILL68_1480 VDD VSS sg13g2_FILL8
XSTDFILL68_1488 VDD VSS sg13g2_FILL8
XSTDFILL68_1496 VDD VSS sg13g2_FILL8
XSTDFILL68_1504 VDD VSS sg13g2_FILL8
XSTDFILL68_1512 VDD VSS sg13g2_FILL8
XSTDFILL68_1520 VDD VSS sg13g2_FILL8
XSTDFILL68_1528 VDD VSS sg13g2_FILL8
XSTDFILL68_1536 VDD VSS sg13g2_FILL8
XSTDFILL68_1544 VDD VSS sg13g2_FILL8
XSTDFILL68_1552 VDD VSS sg13g2_FILL8
XSTDFILL68_1560 VDD VSS sg13g2_FILL8
XSTDFILL68_1568 VDD VSS sg13g2_FILL8
XSTDFILL68_1576 VDD VSS sg13g2_FILL8
XSTDFILL68_1584 VDD VSS sg13g2_FILL8
XSTDFILL68_1592 VDD VSS sg13g2_FILL8
XSTDFILL68_1600 VDD VSS sg13g2_FILL8
XSTDFILL68_1608 VDD VSS sg13g2_FILL8
XSTDFILL68_1616 VDD VSS sg13g2_FILL8
XSTDFILL68_1624 VDD VSS sg13g2_FILL8
XSTDFILL68_1632 VDD VSS sg13g2_FILL8
XSTDFILL68_1640 VDD VSS sg13g2_FILL8
XSTDFILL68_1648 VDD VSS sg13g2_FILL8
XSTDFILL68_1656 VDD VSS sg13g2_FILL8
XSTDFILL68_1664 VDD VSS sg13g2_FILL8
XSTDFILL68_1672 VDD VSS sg13g2_FILL8
XSTDFILL68_1680 VDD VSS sg13g2_FILL8
XSTDFILL68_1688 VDD VSS sg13g2_FILL8
XSTDFILL68_1696 VDD VSS sg13g2_FILL8
XSTDFILL68_1704 VDD VSS sg13g2_FILL8
XSTDFILL68_1712 VDD VSS sg13g2_FILL8
XSTDFILL68_1720 VDD VSS sg13g2_FILL8
XSTDFILL68_1728 VDD VSS sg13g2_FILL8
XSTDFILL68_1736 VDD VSS sg13g2_FILL8
XSTDFILL68_1744 VDD VSS sg13g2_FILL8
XSTDFILL68_1752 VDD VSS sg13g2_FILL8
XSTDFILL68_1760 VDD VSS sg13g2_FILL8
XSTDFILL68_1768 VDD VSS sg13g2_FILL8
XSTDFILL68_1776 VDD VSS sg13g2_FILL8
XSTDFILL68_1784 VDD VSS sg13g2_FILL8
XSTDFILL68_1792 VDD VSS sg13g2_FILL8
XSTDFILL68_1800 VDD VSS sg13g2_FILL8
XSTDFILL68_1808 VDD VSS sg13g2_FILL8
XSTDFILL68_1816 VDD VSS sg13g2_FILL8
XSTDFILL68_1824 VDD VSS sg13g2_FILL8
XSTDFILL68_1832 VDD VSS sg13g2_FILL8
XSTDFILL68_1840 VDD VSS sg13g2_FILL8
XSTDFILL68_1848 VDD VSS sg13g2_FILL8
XSTDFILL68_1856 VDD VSS sg13g2_FILL8
XSTDFILL68_1864 VDD VSS sg13g2_FILL8
XSTDFILL68_1872 VDD VSS sg13g2_FILL8
XSTDFILL68_1880 VDD VSS sg13g2_FILL8
XSTDFILL68_1888 VDD VSS sg13g2_FILL8
XSTDFILL68_1896 VDD VSS sg13g2_FILL8
XSTDFILL68_1904 VDD VSS sg13g2_FILL8
XSTDFILL68_1912 VDD VSS sg13g2_FILL8
XSTDFILL68_1920 VDD VSS sg13g2_FILL8
XSTDFILL68_1928 VDD VSS sg13g2_FILL8
XSTDFILL68_1936 VDD VSS sg13g2_FILL8
XSTDFILL68_1944 VDD VSS sg13g2_FILL8
XSTDFILL68_1952 VDD VSS sg13g2_FILL8
XSTDFILL68_1960 VDD VSS sg13g2_FILL8
XSTDFILL68_1968 VDD VSS sg13g2_FILL8
XSTDFILL68_1976 VDD VSS sg13g2_FILL8
XSTDFILL68_1984 VDD VSS sg13g2_FILL8
XSTDFILL68_1992 VDD VSS sg13g2_FILL8
XSTDFILL68_2000 VDD VSS sg13g2_FILL8
XSTDFILL68_2008 VDD VSS sg13g2_FILL8
XSTDFILL68_2016 VDD VSS sg13g2_FILL8
XSTDFILL68_2024 VDD VSS sg13g2_FILL8
XSTDFILL68_2032 VDD VSS sg13g2_FILL8
XSTDFILL68_2040 VDD VSS sg13g2_FILL8
XSTDFILL68_2048 VDD VSS sg13g2_FILL8
XSTDFILL68_2056 VDD VSS sg13g2_FILL8
XSTDFILL68_2064 VDD VSS sg13g2_FILL8
XSTDFILL68_2072 VDD VSS sg13g2_FILL8
XSTDFILL68_2080 VDD VSS sg13g2_FILL8
XSTDFILL68_2088 VDD VSS sg13g2_FILL8
XSTDFILL68_2096 VDD VSS sg13g2_FILL8
XSTDFILL68_2104 VDD VSS sg13g2_FILL8
XSTDFILL68_2112 VDD VSS sg13g2_FILL8
XSTDFILL68_2120 VDD VSS sg13g2_FILL8
XSTDFILL68_2128 VDD VSS sg13g2_FILL8
XSTDFILL68_2136 VDD VSS sg13g2_FILL8
XSTDFILL68_2144 VDD VSS sg13g2_FILL8
XSTDFILL68_2152 VDD VSS sg13g2_FILL2
XSTDFILL69_0 VDD VSS sg13g2_FILL8
XSTDFILL69_8 VDD VSS sg13g2_FILL8
XSTDFILL69_16 VDD VSS sg13g2_FILL8
XSTDFILL69_24 VDD VSS sg13g2_FILL8
XSTDFILL69_32 VDD VSS sg13g2_FILL8
XSTDFILL69_40 VDD VSS sg13g2_FILL8
XSTDFILL69_48 VDD VSS sg13g2_FILL8
XSTDFILL69_56 VDD VSS sg13g2_FILL8
XSTDFILL69_64 VDD VSS sg13g2_FILL8
XSTDFILL69_72 VDD VSS sg13g2_FILL8
XSTDFILL69_80 VDD VSS sg13g2_FILL8
XSTDFILL69_88 VDD VSS sg13g2_FILL8
XSTDFILL69_96 VDD VSS sg13g2_FILL8
XSTDFILL69_104 VDD VSS sg13g2_FILL8
XSTDFILL69_112 VDD VSS sg13g2_FILL8
XSTDFILL69_120 VDD VSS sg13g2_FILL8
XSTDFILL69_128 VDD VSS sg13g2_FILL4
XSTDFILL69_1085 VDD VSS sg13g2_FILL8
XSTDFILL69_1093 VDD VSS sg13g2_FILL8
XSTDFILL69_1101 VDD VSS sg13g2_FILL8
XSTDFILL69_1109 VDD VSS sg13g2_FILL8
XSTDFILL69_1117 VDD VSS sg13g2_FILL8
XSTDFILL69_1125 VDD VSS sg13g2_FILL8
XSTDFILL69_1133 VDD VSS sg13g2_FILL8
XSTDFILL69_1141 VDD VSS sg13g2_FILL8
XSTDFILL69_1149 VDD VSS sg13g2_FILL8
XSTDFILL69_1157 VDD VSS sg13g2_FILL8
XSTDFILL69_1165 VDD VSS sg13g2_FILL8
XSTDFILL69_1173 VDD VSS sg13g2_FILL8
XSTDFILL69_1181 VDD VSS sg13g2_FILL8
XSTDFILL69_1189 VDD VSS sg13g2_FILL8
XSTDFILL69_1197 VDD VSS sg13g2_FILL8
XSTDFILL69_1205 VDD VSS sg13g2_FILL8
XSTDFILL69_1213 VDD VSS sg13g2_FILL8
XSTDFILL69_1221 VDD VSS sg13g2_FILL8
XSTDFILL69_1229 VDD VSS sg13g2_FILL8
XSTDFILL69_1237 VDD VSS sg13g2_FILL8
XSTDFILL69_1245 VDD VSS sg13g2_FILL8
XSTDFILL69_1253 VDD VSS sg13g2_FILL8
XSTDFILL69_1261 VDD VSS sg13g2_FILL8
XSTDFILL69_1269 VDD VSS sg13g2_FILL8
XSTDFILL69_1277 VDD VSS sg13g2_FILL8
XSTDFILL69_1285 VDD VSS sg13g2_FILL8
XSTDFILL69_1293 VDD VSS sg13g2_FILL8
XSTDFILL69_1301 VDD VSS sg13g2_FILL8
XSTDFILL69_1309 VDD VSS sg13g2_FILL8
XSTDFILL69_1317 VDD VSS sg13g2_FILL8
XSTDFILL69_1325 VDD VSS sg13g2_FILL8
XSTDFILL69_1333 VDD VSS sg13g2_FILL8
XSTDFILL69_1341 VDD VSS sg13g2_FILL8
XSTDFILL69_1349 VDD VSS sg13g2_FILL8
XSTDFILL69_1357 VDD VSS sg13g2_FILL8
XSTDFILL69_1365 VDD VSS sg13g2_FILL8
XSTDFILL69_1373 VDD VSS sg13g2_FILL8
XSTDFILL69_1381 VDD VSS sg13g2_FILL8
XSTDFILL69_1389 VDD VSS sg13g2_FILL8
XSTDFILL69_1397 VDD VSS sg13g2_FILL8
XSTDFILL69_1405 VDD VSS sg13g2_FILL8
XSTDFILL69_1413 VDD VSS sg13g2_FILL8
XSTDFILL69_1421 VDD VSS sg13g2_FILL8
XSTDFILL69_1429 VDD VSS sg13g2_FILL8
XSTDFILL69_1437 VDD VSS sg13g2_FILL8
XSTDFILL69_1445 VDD VSS sg13g2_FILL8
XSTDFILL69_1453 VDD VSS sg13g2_FILL8
XSTDFILL69_1461 VDD VSS sg13g2_FILL8
XSTDFILL69_1469 VDD VSS sg13g2_FILL8
XSTDFILL69_1477 VDD VSS sg13g2_FILL8
XSTDFILL69_1485 VDD VSS sg13g2_FILL8
XSTDFILL69_1493 VDD VSS sg13g2_FILL8
XSTDFILL69_1501 VDD VSS sg13g2_FILL8
XSTDFILL69_1509 VDD VSS sg13g2_FILL8
XSTDFILL69_1517 VDD VSS sg13g2_FILL8
XSTDFILL69_1525 VDD VSS sg13g2_FILL8
XSTDFILL69_1533 VDD VSS sg13g2_FILL8
XSTDFILL69_1541 VDD VSS sg13g2_FILL8
XSTDFILL69_1549 VDD VSS sg13g2_FILL8
XSTDFILL69_1557 VDD VSS sg13g2_FILL8
XSTDFILL69_1565 VDD VSS sg13g2_FILL8
XSTDFILL69_1573 VDD VSS sg13g2_FILL8
XSTDFILL69_1581 VDD VSS sg13g2_FILL8
XSTDFILL69_1589 VDD VSS sg13g2_FILL8
XSTDFILL69_1597 VDD VSS sg13g2_FILL8
XSTDFILL69_1605 VDD VSS sg13g2_FILL8
XSTDFILL69_1613 VDD VSS sg13g2_FILL8
XSTDFILL69_1621 VDD VSS sg13g2_FILL8
XSTDFILL69_1629 VDD VSS sg13g2_FILL8
XSTDFILL69_1637 VDD VSS sg13g2_FILL8
XSTDFILL69_1645 VDD VSS sg13g2_FILL8
XSTDFILL69_1653 VDD VSS sg13g2_FILL8
XSTDFILL69_1661 VDD VSS sg13g2_FILL8
XSTDFILL69_1669 VDD VSS sg13g2_FILL8
XSTDFILL69_1677 VDD VSS sg13g2_FILL8
XSTDFILL69_1685 VDD VSS sg13g2_FILL8
XSTDFILL69_1693 VDD VSS sg13g2_FILL8
XSTDFILL69_1701 VDD VSS sg13g2_FILL8
XSTDFILL69_1709 VDD VSS sg13g2_FILL8
XSTDFILL69_1717 VDD VSS sg13g2_FILL8
XSTDFILL69_1725 VDD VSS sg13g2_FILL8
XSTDFILL69_1733 VDD VSS sg13g2_FILL8
XSTDFILL69_1741 VDD VSS sg13g2_FILL8
XSTDFILL69_1749 VDD VSS sg13g2_FILL8
XSTDFILL69_1757 VDD VSS sg13g2_FILL8
XSTDFILL69_1765 VDD VSS sg13g2_FILL8
XSTDFILL69_1773 VDD VSS sg13g2_FILL8
XSTDFILL69_1781 VDD VSS sg13g2_FILL8
XSTDFILL69_1789 VDD VSS sg13g2_FILL8
XSTDFILL69_1797 VDD VSS sg13g2_FILL8
XSTDFILL69_1805 VDD VSS sg13g2_FILL8
XSTDFILL69_1813 VDD VSS sg13g2_FILL8
XSTDFILL69_1821 VDD VSS sg13g2_FILL8
XSTDFILL69_1829 VDD VSS sg13g2_FILL8
XSTDFILL69_1837 VDD VSS sg13g2_FILL8
XSTDFILL69_1845 VDD VSS sg13g2_FILL8
XSTDFILL69_1853 VDD VSS sg13g2_FILL8
XSTDFILL69_1861 VDD VSS sg13g2_FILL8
XSTDFILL69_1869 VDD VSS sg13g2_FILL8
XSTDFILL69_1877 VDD VSS sg13g2_FILL8
XSTDFILL69_1885 VDD VSS sg13g2_FILL8
XSTDFILL69_1893 VDD VSS sg13g2_FILL8
XSTDFILL69_1901 VDD VSS sg13g2_FILL8
XSTDFILL69_1909 VDD VSS sg13g2_FILL8
XSTDFILL69_1917 VDD VSS sg13g2_FILL8
XSTDFILL69_1925 VDD VSS sg13g2_FILL8
XSTDFILL69_1933 VDD VSS sg13g2_FILL8
XSTDFILL69_1941 VDD VSS sg13g2_FILL8
XSTDFILL69_1949 VDD VSS sg13g2_FILL8
XSTDFILL69_1957 VDD VSS sg13g2_FILL8
XSTDFILL69_1965 VDD VSS sg13g2_FILL8
XSTDFILL69_1973 VDD VSS sg13g2_FILL8
XSTDFILL69_1981 VDD VSS sg13g2_FILL8
XSTDFILL69_1989 VDD VSS sg13g2_FILL8
XSTDFILL69_1997 VDD VSS sg13g2_FILL8
XSTDFILL69_2005 VDD VSS sg13g2_FILL8
XSTDFILL69_2013 VDD VSS sg13g2_FILL8
XSTDFILL69_2021 VDD VSS sg13g2_FILL8
XSTDFILL69_2029 VDD VSS sg13g2_FILL8
XSTDFILL69_2037 VDD VSS sg13g2_FILL8
XSTDFILL69_2045 VDD VSS sg13g2_FILL8
XSTDFILL69_2053 VDD VSS sg13g2_FILL8
XSTDFILL69_2061 VDD VSS sg13g2_FILL8
XSTDFILL69_2069 VDD VSS sg13g2_FILL8
XSTDFILL69_2077 VDD VSS sg13g2_FILL8
XSTDFILL69_2085 VDD VSS sg13g2_FILL8
XSTDFILL69_2093 VDD VSS sg13g2_FILL8
XSTDFILL69_2101 VDD VSS sg13g2_FILL8
XSTDFILL69_2109 VDD VSS sg13g2_FILL8
XSTDFILL69_2117 VDD VSS sg13g2_FILL8
XSTDFILL69_2125 VDD VSS sg13g2_FILL8
XSTDFILL69_2133 VDD VSS sg13g2_FILL8
XSTDFILL69_2141 VDD VSS sg13g2_FILL8
XSTDFILL69_2149 VDD VSS sg13g2_FILL4
XSTDFILL69_2153 VDD VSS sg13g2_FILL1
XSTDFILL70_0 VDD VSS sg13g2_FILL8
XSTDFILL70_8 VDD VSS sg13g2_FILL8
XSTDFILL70_16 VDD VSS sg13g2_FILL8
XSTDFILL70_24 VDD VSS sg13g2_FILL8
XSTDFILL70_32 VDD VSS sg13g2_FILL8
XSTDFILL70_40 VDD VSS sg13g2_FILL8
XSTDFILL70_48 VDD VSS sg13g2_FILL8
XSTDFILL70_56 VDD VSS sg13g2_FILL8
XSTDFILL70_64 VDD VSS sg13g2_FILL8
XSTDFILL70_72 VDD VSS sg13g2_FILL8
XSTDFILL70_80 VDD VSS sg13g2_FILL8
XSTDFILL70_88 VDD VSS sg13g2_FILL8
XSTDFILL70_96 VDD VSS sg13g2_FILL8
XSTDFILL70_104 VDD VSS sg13g2_FILL8
XSTDFILL70_112 VDD VSS sg13g2_FILL8
XSTDFILL70_120 VDD VSS sg13g2_FILL8
XSTDFILL70_128 VDD VSS sg13g2_FILL4
XSTDFILL70_1085 VDD VSS sg13g2_FILL8
XSTDFILL70_1093 VDD VSS sg13g2_FILL8
XSTDFILL70_1101 VDD VSS sg13g2_FILL8
XSTDFILL70_1109 VDD VSS sg13g2_FILL8
XSTDFILL70_1117 VDD VSS sg13g2_FILL8
XSTDFILL70_1125 VDD VSS sg13g2_FILL8
XSTDFILL70_1133 VDD VSS sg13g2_FILL8
XSTDFILL70_1141 VDD VSS sg13g2_FILL8
XSTDFILL70_1149 VDD VSS sg13g2_FILL8
XSTDFILL70_1157 VDD VSS sg13g2_FILL8
XSTDFILL70_1165 VDD VSS sg13g2_FILL8
XSTDFILL70_1173 VDD VSS sg13g2_FILL8
XSTDFILL70_1181 VDD VSS sg13g2_FILL8
XSTDFILL70_1189 VDD VSS sg13g2_FILL8
XSTDFILL70_1197 VDD VSS sg13g2_FILL8
XSTDFILL70_1205 VDD VSS sg13g2_FILL8
XSTDFILL70_1213 VDD VSS sg13g2_FILL8
XSTDFILL70_1221 VDD VSS sg13g2_FILL8
XSTDFILL70_1229 VDD VSS sg13g2_FILL8
XSTDFILL70_1237 VDD VSS sg13g2_FILL8
XSTDFILL70_1245 VDD VSS sg13g2_FILL8
XSTDFILL70_1253 VDD VSS sg13g2_FILL8
XSTDFILL70_1261 VDD VSS sg13g2_FILL8
XSTDFILL70_1269 VDD VSS sg13g2_FILL8
XSTDFILL70_1277 VDD VSS sg13g2_FILL8
XSTDFILL70_1285 VDD VSS sg13g2_FILL8
XSTDFILL70_1293 VDD VSS sg13g2_FILL8
XSTDFILL70_1301 VDD VSS sg13g2_FILL8
XSTDFILL70_1309 VDD VSS sg13g2_FILL8
XSTDFILL70_1317 VDD VSS sg13g2_FILL8
XSTDFILL70_1325 VDD VSS sg13g2_FILL8
XSTDFILL70_1333 VDD VSS sg13g2_FILL8
XSTDFILL70_1341 VDD VSS sg13g2_FILL8
XSTDFILL70_1349 VDD VSS sg13g2_FILL8
XSTDFILL70_1357 VDD VSS sg13g2_FILL8
XSTDFILL70_1365 VDD VSS sg13g2_FILL8
XSTDFILL70_1373 VDD VSS sg13g2_FILL8
XSTDFILL70_1381 VDD VSS sg13g2_FILL8
XSTDFILL70_1389 VDD VSS sg13g2_FILL8
XSTDFILL70_1397 VDD VSS sg13g2_FILL8
XSTDFILL70_1405 VDD VSS sg13g2_FILL8
XSTDFILL70_1413 VDD VSS sg13g2_FILL8
XSTDFILL70_1421 VDD VSS sg13g2_FILL8
XSTDFILL70_1429 VDD VSS sg13g2_FILL8
XSTDFILL70_1437 VDD VSS sg13g2_FILL8
XSTDFILL70_1445 VDD VSS sg13g2_FILL8
XSTDFILL70_1453 VDD VSS sg13g2_FILL8
XSTDFILL70_1461 VDD VSS sg13g2_FILL8
XSTDFILL70_1469 VDD VSS sg13g2_FILL8
XSTDFILL70_1477 VDD VSS sg13g2_FILL8
XSTDFILL70_1485 VDD VSS sg13g2_FILL8
XSTDFILL70_1493 VDD VSS sg13g2_FILL8
XSTDFILL70_1501 VDD VSS sg13g2_FILL8
XSTDFILL70_1509 VDD VSS sg13g2_FILL8
XSTDFILL70_1517 VDD VSS sg13g2_FILL8
XSTDFILL70_1525 VDD VSS sg13g2_FILL8
XSTDFILL70_1533 VDD VSS sg13g2_FILL8
XSTDFILL70_1541 VDD VSS sg13g2_FILL8
XSTDFILL70_1549 VDD VSS sg13g2_FILL8
XSTDFILL70_1557 VDD VSS sg13g2_FILL8
XSTDFILL70_1565 VDD VSS sg13g2_FILL8
XSTDFILL70_1573 VDD VSS sg13g2_FILL8
XSTDFILL70_1581 VDD VSS sg13g2_FILL8
XSTDFILL70_1589 VDD VSS sg13g2_FILL8
XSTDFILL70_1597 VDD VSS sg13g2_FILL8
XSTDFILL70_1605 VDD VSS sg13g2_FILL8
XSTDFILL70_1613 VDD VSS sg13g2_FILL8
XSTDFILL70_1621 VDD VSS sg13g2_FILL8
XSTDFILL70_1629 VDD VSS sg13g2_FILL8
XSTDFILL70_1637 VDD VSS sg13g2_FILL8
XSTDFILL70_1645 VDD VSS sg13g2_FILL8
XSTDFILL70_1653 VDD VSS sg13g2_FILL8
XSTDFILL70_1661 VDD VSS sg13g2_FILL8
XSTDFILL70_1669 VDD VSS sg13g2_FILL8
XSTDFILL70_1677 VDD VSS sg13g2_FILL8
XSTDFILL70_1685 VDD VSS sg13g2_FILL8
XSTDFILL70_1693 VDD VSS sg13g2_FILL8
XSTDFILL70_1701 VDD VSS sg13g2_FILL8
XSTDFILL70_1709 VDD VSS sg13g2_FILL8
XSTDFILL70_1717 VDD VSS sg13g2_FILL8
XSTDFILL70_1725 VDD VSS sg13g2_FILL8
XSTDFILL70_1733 VDD VSS sg13g2_FILL8
XSTDFILL70_1741 VDD VSS sg13g2_FILL8
XSTDFILL70_1749 VDD VSS sg13g2_FILL8
XSTDFILL70_1757 VDD VSS sg13g2_FILL8
XSTDFILL70_1765 VDD VSS sg13g2_FILL8
XSTDFILL70_1773 VDD VSS sg13g2_FILL8
XSTDFILL70_1781 VDD VSS sg13g2_FILL8
XSTDFILL70_1789 VDD VSS sg13g2_FILL8
XSTDFILL70_1797 VDD VSS sg13g2_FILL8
XSTDFILL70_1805 VDD VSS sg13g2_FILL8
XSTDFILL70_1813 VDD VSS sg13g2_FILL8
XSTDFILL70_1821 VDD VSS sg13g2_FILL8
XSTDFILL70_1829 VDD VSS sg13g2_FILL8
XSTDFILL70_1837 VDD VSS sg13g2_FILL8
XSTDFILL70_1845 VDD VSS sg13g2_FILL8
XSTDFILL70_1853 VDD VSS sg13g2_FILL8
XSTDFILL70_1861 VDD VSS sg13g2_FILL8
XSTDFILL70_1869 VDD VSS sg13g2_FILL8
XSTDFILL70_1877 VDD VSS sg13g2_FILL8
XSTDFILL70_1885 VDD VSS sg13g2_FILL8
XSTDFILL70_1893 VDD VSS sg13g2_FILL8
XSTDFILL70_1901 VDD VSS sg13g2_FILL8
XSTDFILL70_1909 VDD VSS sg13g2_FILL8
XSTDFILL70_1917 VDD VSS sg13g2_FILL8
XSTDFILL70_1925 VDD VSS sg13g2_FILL8
XSTDFILL70_1933 VDD VSS sg13g2_FILL8
XSTDFILL70_1941 VDD VSS sg13g2_FILL8
XSTDFILL70_1949 VDD VSS sg13g2_FILL8
XSTDFILL70_1957 VDD VSS sg13g2_FILL8
XSTDFILL70_1965 VDD VSS sg13g2_FILL8
XSTDFILL70_1973 VDD VSS sg13g2_FILL8
XSTDFILL70_1981 VDD VSS sg13g2_FILL8
XSTDFILL70_1989 VDD VSS sg13g2_FILL8
XSTDFILL70_1997 VDD VSS sg13g2_FILL8
XSTDFILL70_2005 VDD VSS sg13g2_FILL8
XSTDFILL70_2013 VDD VSS sg13g2_FILL8
XSTDFILL70_2021 VDD VSS sg13g2_FILL8
XSTDFILL70_2029 VDD VSS sg13g2_FILL8
XSTDFILL70_2037 VDD VSS sg13g2_FILL8
XSTDFILL70_2045 VDD VSS sg13g2_FILL8
XSTDFILL70_2053 VDD VSS sg13g2_FILL8
XSTDFILL70_2061 VDD VSS sg13g2_FILL8
XSTDFILL70_2069 VDD VSS sg13g2_FILL8
XSTDFILL70_2077 VDD VSS sg13g2_FILL8
XSTDFILL70_2085 VDD VSS sg13g2_FILL8
XSTDFILL70_2093 VDD VSS sg13g2_FILL8
XSTDFILL70_2101 VDD VSS sg13g2_FILL8
XSTDFILL70_2109 VDD VSS sg13g2_FILL8
XSTDFILL70_2117 VDD VSS sg13g2_FILL8
XSTDFILL70_2125 VDD VSS sg13g2_FILL8
XSTDFILL70_2133 VDD VSS sg13g2_FILL8
XSTDFILL70_2141 VDD VSS sg13g2_FILL8
XSTDFILL70_2149 VDD VSS sg13g2_FILL4
XSTDFILL70_2153 VDD VSS sg13g2_FILL1
XSTDFILL71_0 VDD VSS sg13g2_FILL8
XSTDFILL71_8 VDD VSS sg13g2_FILL8
XSTDFILL71_16 VDD VSS sg13g2_FILL8
XSTDFILL71_24 VDD VSS sg13g2_FILL8
XSTDFILL71_32 VDD VSS sg13g2_FILL8
XSTDFILL71_40 VDD VSS sg13g2_FILL8
XSTDFILL71_48 VDD VSS sg13g2_FILL8
XSTDFILL71_56 VDD VSS sg13g2_FILL8
XSTDFILL71_64 VDD VSS sg13g2_FILL8
XSTDFILL71_72 VDD VSS sg13g2_FILL8
XSTDFILL71_80 VDD VSS sg13g2_FILL8
XSTDFILL71_88 VDD VSS sg13g2_FILL8
XSTDFILL71_96 VDD VSS sg13g2_FILL8
XSTDFILL71_104 VDD VSS sg13g2_FILL8
XSTDFILL71_112 VDD VSS sg13g2_FILL8
XSTDFILL71_120 VDD VSS sg13g2_FILL8
XSTDFILL71_128 VDD VSS sg13g2_FILL4
XSTDFILL71_1085 VDD VSS sg13g2_FILL8
XSTDFILL71_1093 VDD VSS sg13g2_FILL8
XSTDFILL71_1101 VDD VSS sg13g2_FILL8
XSTDFILL71_1109 VDD VSS sg13g2_FILL8
XSTDFILL71_1117 VDD VSS sg13g2_FILL8
XSTDFILL71_1125 VDD VSS sg13g2_FILL8
XSTDFILL71_1133 VDD VSS sg13g2_FILL8
XSTDFILL71_1141 VDD VSS sg13g2_FILL8
XSTDFILL71_1149 VDD VSS sg13g2_FILL8
XSTDFILL71_1157 VDD VSS sg13g2_FILL8
XSTDFILL71_1165 VDD VSS sg13g2_FILL8
XSTDFILL71_1173 VDD VSS sg13g2_FILL8
XSTDFILL71_1181 VDD VSS sg13g2_FILL8
XSTDFILL71_1189 VDD VSS sg13g2_FILL8
XSTDFILL71_1197 VDD VSS sg13g2_FILL8
XSTDFILL71_1205 VDD VSS sg13g2_FILL8
XSTDFILL71_1213 VDD VSS sg13g2_FILL8
XSTDFILL71_1221 VDD VSS sg13g2_FILL8
XSTDFILL71_1229 VDD VSS sg13g2_FILL8
XSTDFILL71_1237 VDD VSS sg13g2_FILL8
XSTDFILL71_1245 VDD VSS sg13g2_FILL8
XSTDFILL71_1253 VDD VSS sg13g2_FILL8
XSTDFILL71_1261 VDD VSS sg13g2_FILL8
XSTDFILL71_1269 VDD VSS sg13g2_FILL8
XSTDFILL71_1277 VDD VSS sg13g2_FILL8
XSTDFILL71_1285 VDD VSS sg13g2_FILL8
XSTDFILL71_1293 VDD VSS sg13g2_FILL8
XSTDFILL71_1301 VDD VSS sg13g2_FILL8
XSTDFILL71_1309 VDD VSS sg13g2_FILL8
XSTDFILL71_1317 VDD VSS sg13g2_FILL8
XSTDFILL71_1325 VDD VSS sg13g2_FILL8
XSTDFILL71_1333 VDD VSS sg13g2_FILL8
XSTDFILL71_1341 VDD VSS sg13g2_FILL8
XSTDFILL71_1349 VDD VSS sg13g2_FILL8
XSTDFILL71_1357 VDD VSS sg13g2_FILL8
XSTDFILL71_1365 VDD VSS sg13g2_FILL8
XSTDFILL71_1373 VDD VSS sg13g2_FILL8
XSTDFILL71_1381 VDD VSS sg13g2_FILL8
XSTDFILL71_1389 VDD VSS sg13g2_FILL8
XSTDFILL71_1397 VDD VSS sg13g2_FILL8
XSTDFILL71_1405 VDD VSS sg13g2_FILL8
XSTDFILL71_1413 VDD VSS sg13g2_FILL8
XSTDFILL71_1421 VDD VSS sg13g2_FILL8
XSTDFILL71_1429 VDD VSS sg13g2_FILL8
XSTDFILL71_1437 VDD VSS sg13g2_FILL8
XSTDFILL71_1445 VDD VSS sg13g2_FILL8
XSTDFILL71_1453 VDD VSS sg13g2_FILL8
XSTDFILL71_1461 VDD VSS sg13g2_FILL8
XSTDFILL71_1469 VDD VSS sg13g2_FILL8
XSTDFILL71_1477 VDD VSS sg13g2_FILL8
XSTDFILL71_1485 VDD VSS sg13g2_FILL8
XSTDFILL71_1493 VDD VSS sg13g2_FILL8
XSTDFILL71_1501 VDD VSS sg13g2_FILL8
XSTDFILL71_1509 VDD VSS sg13g2_FILL8
XSTDFILL71_1517 VDD VSS sg13g2_FILL8
XSTDFILL71_1525 VDD VSS sg13g2_FILL8
XSTDFILL71_1533 VDD VSS sg13g2_FILL8
XSTDFILL71_1541 VDD VSS sg13g2_FILL8
XSTDFILL71_1549 VDD VSS sg13g2_FILL8
XSTDFILL71_1557 VDD VSS sg13g2_FILL8
XSTDFILL71_1565 VDD VSS sg13g2_FILL8
XSTDFILL71_1573 VDD VSS sg13g2_FILL8
XSTDFILL71_1581 VDD VSS sg13g2_FILL8
XSTDFILL71_1589 VDD VSS sg13g2_FILL8
XSTDFILL71_1597 VDD VSS sg13g2_FILL8
XSTDFILL71_1605 VDD VSS sg13g2_FILL8
XSTDFILL71_1613 VDD VSS sg13g2_FILL8
XSTDFILL71_1621 VDD VSS sg13g2_FILL8
XSTDFILL71_1629 VDD VSS sg13g2_FILL8
XSTDFILL71_1637 VDD VSS sg13g2_FILL8
XSTDFILL71_1645 VDD VSS sg13g2_FILL8
XSTDFILL71_1653 VDD VSS sg13g2_FILL8
XSTDFILL71_1661 VDD VSS sg13g2_FILL8
XSTDFILL71_1669 VDD VSS sg13g2_FILL8
XSTDFILL71_1677 VDD VSS sg13g2_FILL8
XSTDFILL71_1685 VDD VSS sg13g2_FILL8
XSTDFILL71_1693 VDD VSS sg13g2_FILL8
XSTDFILL71_1701 VDD VSS sg13g2_FILL8
XSTDFILL71_1709 VDD VSS sg13g2_FILL8
XSTDFILL71_1717 VDD VSS sg13g2_FILL8
XSTDFILL71_1725 VDD VSS sg13g2_FILL8
XSTDFILL71_1733 VDD VSS sg13g2_FILL8
XSTDFILL71_1741 VDD VSS sg13g2_FILL8
XSTDFILL71_1749 VDD VSS sg13g2_FILL8
XSTDFILL71_1757 VDD VSS sg13g2_FILL8
XSTDFILL71_1765 VDD VSS sg13g2_FILL8
XSTDFILL71_1773 VDD VSS sg13g2_FILL8
XSTDFILL71_1781 VDD VSS sg13g2_FILL8
XSTDFILL71_1789 VDD VSS sg13g2_FILL8
XSTDFILL71_1797 VDD VSS sg13g2_FILL8
XSTDFILL71_1805 VDD VSS sg13g2_FILL8
XSTDFILL71_1813 VDD VSS sg13g2_FILL8
XSTDFILL71_1821 VDD VSS sg13g2_FILL8
XSTDFILL71_1829 VDD VSS sg13g2_FILL8
XSTDFILL71_1837 VDD VSS sg13g2_FILL8
XSTDFILL71_1845 VDD VSS sg13g2_FILL8
XSTDFILL71_1853 VDD VSS sg13g2_FILL8
XSTDFILL71_1861 VDD VSS sg13g2_FILL8
XSTDFILL71_1869 VDD VSS sg13g2_FILL8
XSTDFILL71_1877 VDD VSS sg13g2_FILL8
XSTDFILL71_1885 VDD VSS sg13g2_FILL8
XSTDFILL71_1893 VDD VSS sg13g2_FILL8
XSTDFILL71_1901 VDD VSS sg13g2_FILL8
XSTDFILL71_1909 VDD VSS sg13g2_FILL8
XSTDFILL71_1917 VDD VSS sg13g2_FILL8
XSTDFILL71_1925 VDD VSS sg13g2_FILL8
XSTDFILL71_1933 VDD VSS sg13g2_FILL8
XSTDFILL71_1941 VDD VSS sg13g2_FILL8
XSTDFILL71_1949 VDD VSS sg13g2_FILL8
XSTDFILL71_1957 VDD VSS sg13g2_FILL8
XSTDFILL71_1965 VDD VSS sg13g2_FILL8
XSTDFILL71_1973 VDD VSS sg13g2_FILL8
XSTDFILL71_1981 VDD VSS sg13g2_FILL8
XSTDFILL71_1989 VDD VSS sg13g2_FILL8
XSTDFILL71_1997 VDD VSS sg13g2_FILL8
XSTDFILL71_2005 VDD VSS sg13g2_FILL8
XSTDFILL71_2013 VDD VSS sg13g2_FILL8
XSTDFILL71_2021 VDD VSS sg13g2_FILL8
XSTDFILL71_2029 VDD VSS sg13g2_FILL8
XSTDFILL71_2037 VDD VSS sg13g2_FILL8
XSTDFILL71_2045 VDD VSS sg13g2_FILL8
XSTDFILL71_2053 VDD VSS sg13g2_FILL8
XSTDFILL71_2061 VDD VSS sg13g2_FILL8
XSTDFILL71_2069 VDD VSS sg13g2_FILL8
XSTDFILL71_2077 VDD VSS sg13g2_FILL8
XSTDFILL71_2085 VDD VSS sg13g2_FILL8
XSTDFILL71_2093 VDD VSS sg13g2_FILL8
XSTDFILL71_2101 VDD VSS sg13g2_FILL8
XSTDFILL71_2109 VDD VSS sg13g2_FILL8
XSTDFILL71_2117 VDD VSS sg13g2_FILL8
XSTDFILL71_2125 VDD VSS sg13g2_FILL8
XSTDFILL71_2133 VDD VSS sg13g2_FILL8
XSTDFILL71_2141 VDD VSS sg13g2_FILL8
XSTDFILL71_2149 VDD VSS sg13g2_FILL4
XSTDFILL71_2153 VDD VSS sg13g2_FILL1
XSTDFILL72_0 VDD VSS sg13g2_FILL8
XSTDFILL72_8 VDD VSS sg13g2_FILL8
XSTDFILL72_16 VDD VSS sg13g2_FILL8
XSTDFILL72_24 VDD VSS sg13g2_FILL8
XSTDFILL72_32 VDD VSS sg13g2_FILL8
XSTDFILL72_40 VDD VSS sg13g2_FILL8
XSTDFILL72_48 VDD VSS sg13g2_FILL8
XSTDFILL72_56 VDD VSS sg13g2_FILL8
XSTDFILL72_64 VDD VSS sg13g2_FILL8
XSTDFILL72_72 VDD VSS sg13g2_FILL8
XSTDFILL72_80 VDD VSS sg13g2_FILL8
XSTDFILL72_88 VDD VSS sg13g2_FILL8
XSTDFILL72_96 VDD VSS sg13g2_FILL8
XSTDFILL72_104 VDD VSS sg13g2_FILL8
XSTDFILL72_112 VDD VSS sg13g2_FILL8
XSTDFILL72_120 VDD VSS sg13g2_FILL8
XSTDFILL72_128 VDD VSS sg13g2_FILL4
XSTDFILL72_1085 VDD VSS sg13g2_FILL8
XSTDFILL72_1093 VDD VSS sg13g2_FILL8
XSTDFILL72_1101 VDD VSS sg13g2_FILL8
XSTDFILL72_1109 VDD VSS sg13g2_FILL8
XSTDFILL72_1117 VDD VSS sg13g2_FILL8
XSTDFILL72_1125 VDD VSS sg13g2_FILL8
XSTDFILL72_1133 VDD VSS sg13g2_FILL8
XSTDFILL72_1141 VDD VSS sg13g2_FILL8
XSTDFILL72_1149 VDD VSS sg13g2_FILL8
XSTDFILL72_1157 VDD VSS sg13g2_FILL8
XSTDFILL72_1165 VDD VSS sg13g2_FILL8
XSTDFILL72_1173 VDD VSS sg13g2_FILL8
XSTDFILL72_1181 VDD VSS sg13g2_FILL8
XSTDFILL72_1189 VDD VSS sg13g2_FILL8
XSTDFILL72_1197 VDD VSS sg13g2_FILL8
XSTDFILL72_1205 VDD VSS sg13g2_FILL8
XSTDFILL72_1213 VDD VSS sg13g2_FILL8
XSTDFILL72_1221 VDD VSS sg13g2_FILL8
XSTDFILL72_1229 VDD VSS sg13g2_FILL8
XSTDFILL72_1237 VDD VSS sg13g2_FILL8
XSTDFILL72_1245 VDD VSS sg13g2_FILL8
XSTDFILL72_1253 VDD VSS sg13g2_FILL8
XSTDFILL72_1261 VDD VSS sg13g2_FILL8
XSTDFILL72_1269 VDD VSS sg13g2_FILL8
XSTDFILL72_1277 VDD VSS sg13g2_FILL8
XSTDFILL72_1285 VDD VSS sg13g2_FILL8
XSTDFILL72_1293 VDD VSS sg13g2_FILL8
XSTDFILL72_1301 VDD VSS sg13g2_FILL8
XSTDFILL72_1309 VDD VSS sg13g2_FILL8
XSTDFILL72_1317 VDD VSS sg13g2_FILL8
XSTDFILL72_1325 VDD VSS sg13g2_FILL8
XSTDFILL72_1333 VDD VSS sg13g2_FILL8
XSTDFILL72_1341 VDD VSS sg13g2_FILL8
XSTDFILL72_1349 VDD VSS sg13g2_FILL8
XSTDFILL72_1357 VDD VSS sg13g2_FILL8
XSTDFILL72_1365 VDD VSS sg13g2_FILL8
XSTDFILL72_1373 VDD VSS sg13g2_FILL8
XSTDFILL72_1381 VDD VSS sg13g2_FILL8
XSTDFILL72_1389 VDD VSS sg13g2_FILL8
XSTDFILL72_1397 VDD VSS sg13g2_FILL8
XSTDFILL72_1405 VDD VSS sg13g2_FILL8
XSTDFILL72_1413 VDD VSS sg13g2_FILL8
XSTDFILL72_1421 VDD VSS sg13g2_FILL8
XSTDFILL72_1429 VDD VSS sg13g2_FILL8
XSTDFILL72_1437 VDD VSS sg13g2_FILL8
XSTDFILL72_1445 VDD VSS sg13g2_FILL8
XSTDFILL72_1453 VDD VSS sg13g2_FILL8
XSTDFILL72_1461 VDD VSS sg13g2_FILL8
XSTDFILL72_1469 VDD VSS sg13g2_FILL8
XSTDFILL72_1477 VDD VSS sg13g2_FILL8
XSTDFILL72_1485 VDD VSS sg13g2_FILL8
XSTDFILL72_1493 VDD VSS sg13g2_FILL8
XSTDFILL72_1501 VDD VSS sg13g2_FILL8
XSTDFILL72_1509 VDD VSS sg13g2_FILL8
XSTDFILL72_1517 VDD VSS sg13g2_FILL8
XSTDFILL72_1525 VDD VSS sg13g2_FILL8
XSTDFILL72_1533 VDD VSS sg13g2_FILL8
XSTDFILL72_1541 VDD VSS sg13g2_FILL8
XSTDFILL72_1549 VDD VSS sg13g2_FILL8
XSTDFILL72_1557 VDD VSS sg13g2_FILL8
XSTDFILL72_1565 VDD VSS sg13g2_FILL8
XSTDFILL72_1573 VDD VSS sg13g2_FILL8
XSTDFILL72_1581 VDD VSS sg13g2_FILL8
XSTDFILL72_1589 VDD VSS sg13g2_FILL8
XSTDFILL72_1597 VDD VSS sg13g2_FILL8
XSTDFILL72_1605 VDD VSS sg13g2_FILL8
XSTDFILL72_1613 VDD VSS sg13g2_FILL8
XSTDFILL72_1621 VDD VSS sg13g2_FILL8
XSTDFILL72_1629 VDD VSS sg13g2_FILL8
XSTDFILL72_1637 VDD VSS sg13g2_FILL8
XSTDFILL72_1645 VDD VSS sg13g2_FILL8
XSTDFILL72_1653 VDD VSS sg13g2_FILL8
XSTDFILL72_1661 VDD VSS sg13g2_FILL8
XSTDFILL72_1669 VDD VSS sg13g2_FILL8
XSTDFILL72_1677 VDD VSS sg13g2_FILL8
XSTDFILL72_1685 VDD VSS sg13g2_FILL8
XSTDFILL72_1693 VDD VSS sg13g2_FILL8
XSTDFILL72_1701 VDD VSS sg13g2_FILL8
XSTDFILL72_1709 VDD VSS sg13g2_FILL8
XSTDFILL72_1717 VDD VSS sg13g2_FILL8
XSTDFILL72_1725 VDD VSS sg13g2_FILL8
XSTDFILL72_1733 VDD VSS sg13g2_FILL8
XSTDFILL72_1741 VDD VSS sg13g2_FILL8
XSTDFILL72_1749 VDD VSS sg13g2_FILL8
XSTDFILL72_1757 VDD VSS sg13g2_FILL8
XSTDFILL72_1765 VDD VSS sg13g2_FILL8
XSTDFILL72_1773 VDD VSS sg13g2_FILL8
XSTDFILL72_1781 VDD VSS sg13g2_FILL8
XSTDFILL72_1789 VDD VSS sg13g2_FILL8
XSTDFILL72_1797 VDD VSS sg13g2_FILL8
XSTDFILL72_1805 VDD VSS sg13g2_FILL8
XSTDFILL72_1813 VDD VSS sg13g2_FILL8
XSTDFILL72_1821 VDD VSS sg13g2_FILL8
XSTDFILL72_1829 VDD VSS sg13g2_FILL8
XSTDFILL72_1837 VDD VSS sg13g2_FILL8
XSTDFILL72_1845 VDD VSS sg13g2_FILL8
XSTDFILL72_1853 VDD VSS sg13g2_FILL8
XSTDFILL72_1861 VDD VSS sg13g2_FILL8
XSTDFILL72_1869 VDD VSS sg13g2_FILL8
XSTDFILL72_1877 VDD VSS sg13g2_FILL8
XSTDFILL72_1885 VDD VSS sg13g2_FILL8
XSTDFILL72_1893 VDD VSS sg13g2_FILL8
XSTDFILL72_1901 VDD VSS sg13g2_FILL8
XSTDFILL72_1909 VDD VSS sg13g2_FILL8
XSTDFILL72_1917 VDD VSS sg13g2_FILL8
XSTDFILL72_1925 VDD VSS sg13g2_FILL8
XSTDFILL72_1933 VDD VSS sg13g2_FILL8
XSTDFILL72_1941 VDD VSS sg13g2_FILL8
XSTDFILL72_1949 VDD VSS sg13g2_FILL8
XSTDFILL72_1957 VDD VSS sg13g2_FILL8
XSTDFILL72_1965 VDD VSS sg13g2_FILL8
XSTDFILL72_1973 VDD VSS sg13g2_FILL8
XSTDFILL72_1981 VDD VSS sg13g2_FILL8
XSTDFILL72_1989 VDD VSS sg13g2_FILL8
XSTDFILL72_1997 VDD VSS sg13g2_FILL8
XSTDFILL72_2005 VDD VSS sg13g2_FILL8
XSTDFILL72_2013 VDD VSS sg13g2_FILL8
XSTDFILL72_2021 VDD VSS sg13g2_FILL8
XSTDFILL72_2029 VDD VSS sg13g2_FILL8
XSTDFILL72_2037 VDD VSS sg13g2_FILL8
XSTDFILL72_2045 VDD VSS sg13g2_FILL8
XSTDFILL72_2053 VDD VSS sg13g2_FILL8
XSTDFILL72_2061 VDD VSS sg13g2_FILL8
XSTDFILL72_2069 VDD VSS sg13g2_FILL8
XSTDFILL72_2077 VDD VSS sg13g2_FILL8
XSTDFILL72_2085 VDD VSS sg13g2_FILL8
XSTDFILL72_2093 VDD VSS sg13g2_FILL8
XSTDFILL72_2101 VDD VSS sg13g2_FILL8
XSTDFILL72_2109 VDD VSS sg13g2_FILL8
XSTDFILL72_2117 VDD VSS sg13g2_FILL8
XSTDFILL72_2125 VDD VSS sg13g2_FILL8
XSTDFILL72_2133 VDD VSS sg13g2_FILL8
XSTDFILL72_2141 VDD VSS sg13g2_FILL8
XSTDFILL72_2149 VDD VSS sg13g2_FILL4
XSTDFILL72_2153 VDD VSS sg13g2_FILL1
XSTDFILL73_0 VDD VSS sg13g2_FILL8
XSTDFILL73_8 VDD VSS sg13g2_FILL8
XSTDFILL73_16 VDD VSS sg13g2_FILL8
XSTDFILL73_24 VDD VSS sg13g2_FILL8
XSTDFILL73_32 VDD VSS sg13g2_FILL8
XSTDFILL73_40 VDD VSS sg13g2_FILL8
XSTDFILL73_48 VDD VSS sg13g2_FILL8
XSTDFILL73_56 VDD VSS sg13g2_FILL8
XSTDFILL73_64 VDD VSS sg13g2_FILL8
XSTDFILL73_72 VDD VSS sg13g2_FILL8
XSTDFILL73_80 VDD VSS sg13g2_FILL8
XSTDFILL73_88 VDD VSS sg13g2_FILL8
XSTDFILL73_96 VDD VSS sg13g2_FILL8
XSTDFILL73_104 VDD VSS sg13g2_FILL8
XSTDFILL73_112 VDD VSS sg13g2_FILL8
XSTDFILL73_120 VDD VSS sg13g2_FILL8
XSTDFILL73_128 VDD VSS sg13g2_FILL4
XSTDFILL73_1085 VDD VSS sg13g2_FILL8
XSTDFILL73_1093 VDD VSS sg13g2_FILL8
XSTDFILL73_1101 VDD VSS sg13g2_FILL8
XSTDFILL73_1109 VDD VSS sg13g2_FILL8
XSTDFILL73_1117 VDD VSS sg13g2_FILL8
XSTDFILL73_1125 VDD VSS sg13g2_FILL8
XSTDFILL73_1133 VDD VSS sg13g2_FILL8
XSTDFILL73_1141 VDD VSS sg13g2_FILL8
XSTDFILL73_1149 VDD VSS sg13g2_FILL8
XSTDFILL73_1157 VDD VSS sg13g2_FILL8
XSTDFILL73_1165 VDD VSS sg13g2_FILL8
XSTDFILL73_1173 VDD VSS sg13g2_FILL8
XSTDFILL73_1181 VDD VSS sg13g2_FILL8
XSTDFILL73_1189 VDD VSS sg13g2_FILL8
XSTDFILL73_1197 VDD VSS sg13g2_FILL8
XSTDFILL73_1205 VDD VSS sg13g2_FILL8
XSTDFILL73_1213 VDD VSS sg13g2_FILL8
XSTDFILL73_1221 VDD VSS sg13g2_FILL8
XSTDFILL73_1229 VDD VSS sg13g2_FILL8
XSTDFILL73_1237 VDD VSS sg13g2_FILL8
XSTDFILL73_1245 VDD VSS sg13g2_FILL8
XSTDFILL73_1253 VDD VSS sg13g2_FILL8
XSTDFILL73_1261 VDD VSS sg13g2_FILL8
XSTDFILL73_1269 VDD VSS sg13g2_FILL8
XSTDFILL73_1277 VDD VSS sg13g2_FILL8
XSTDFILL73_1285 VDD VSS sg13g2_FILL8
XSTDFILL73_1293 VDD VSS sg13g2_FILL8
XSTDFILL73_1301 VDD VSS sg13g2_FILL8
XSTDFILL73_1309 VDD VSS sg13g2_FILL8
XSTDFILL73_1317 VDD VSS sg13g2_FILL8
XSTDFILL73_1325 VDD VSS sg13g2_FILL8
XSTDFILL73_1333 VDD VSS sg13g2_FILL8
XSTDFILL73_1341 VDD VSS sg13g2_FILL8
XSTDFILL73_1349 VDD VSS sg13g2_FILL8
XSTDFILL73_1357 VDD VSS sg13g2_FILL8
XSTDFILL73_1365 VDD VSS sg13g2_FILL8
XSTDFILL73_1373 VDD VSS sg13g2_FILL8
XSTDFILL73_1381 VDD VSS sg13g2_FILL8
XSTDFILL73_1389 VDD VSS sg13g2_FILL8
XSTDFILL73_1397 VDD VSS sg13g2_FILL8
XSTDFILL73_1405 VDD VSS sg13g2_FILL8
XSTDFILL73_1413 VDD VSS sg13g2_FILL8
XSTDFILL73_1421 VDD VSS sg13g2_FILL8
XSTDFILL73_1429 VDD VSS sg13g2_FILL8
XSTDFILL73_1437 VDD VSS sg13g2_FILL8
XSTDFILL73_1445 VDD VSS sg13g2_FILL8
XSTDFILL73_1453 VDD VSS sg13g2_FILL8
XSTDFILL73_1461 VDD VSS sg13g2_FILL8
XSTDFILL73_1469 VDD VSS sg13g2_FILL8
XSTDFILL73_1477 VDD VSS sg13g2_FILL8
XSTDFILL73_1485 VDD VSS sg13g2_FILL8
XSTDFILL73_1493 VDD VSS sg13g2_FILL8
XSTDFILL73_1501 VDD VSS sg13g2_FILL8
XSTDFILL73_1509 VDD VSS sg13g2_FILL8
XSTDFILL73_1517 VDD VSS sg13g2_FILL8
XSTDFILL73_1525 VDD VSS sg13g2_FILL8
XSTDFILL73_1533 VDD VSS sg13g2_FILL8
XSTDFILL73_1541 VDD VSS sg13g2_FILL8
XSTDFILL73_1549 VDD VSS sg13g2_FILL8
XSTDFILL73_1557 VDD VSS sg13g2_FILL8
XSTDFILL73_1565 VDD VSS sg13g2_FILL8
XSTDFILL73_1573 VDD VSS sg13g2_FILL8
XSTDFILL73_1581 VDD VSS sg13g2_FILL8
XSTDFILL73_1589 VDD VSS sg13g2_FILL8
XSTDFILL73_1597 VDD VSS sg13g2_FILL8
XSTDFILL73_1605 VDD VSS sg13g2_FILL8
XSTDFILL73_1613 VDD VSS sg13g2_FILL8
XSTDFILL73_1621 VDD VSS sg13g2_FILL8
XSTDFILL73_1629 VDD VSS sg13g2_FILL8
XSTDFILL73_1637 VDD VSS sg13g2_FILL8
XSTDFILL73_1645 VDD VSS sg13g2_FILL8
XSTDFILL73_1653 VDD VSS sg13g2_FILL8
XSTDFILL73_1661 VDD VSS sg13g2_FILL8
XSTDFILL73_1669 VDD VSS sg13g2_FILL8
XSTDFILL73_1677 VDD VSS sg13g2_FILL8
XSTDFILL73_1685 VDD VSS sg13g2_FILL8
XSTDFILL73_1693 VDD VSS sg13g2_FILL8
XSTDFILL73_1701 VDD VSS sg13g2_FILL8
XSTDFILL73_1709 VDD VSS sg13g2_FILL8
XSTDFILL73_1717 VDD VSS sg13g2_FILL8
XSTDFILL73_1725 VDD VSS sg13g2_FILL8
XSTDFILL73_1733 VDD VSS sg13g2_FILL8
XSTDFILL73_1741 VDD VSS sg13g2_FILL8
XSTDFILL73_1749 VDD VSS sg13g2_FILL8
XSTDFILL73_1757 VDD VSS sg13g2_FILL8
XSTDFILL73_1765 VDD VSS sg13g2_FILL8
XSTDFILL73_1773 VDD VSS sg13g2_FILL8
XSTDFILL73_1781 VDD VSS sg13g2_FILL8
XSTDFILL73_1789 VDD VSS sg13g2_FILL8
XSTDFILL73_1797 VDD VSS sg13g2_FILL8
XSTDFILL73_1805 VDD VSS sg13g2_FILL8
XSTDFILL73_1813 VDD VSS sg13g2_FILL8
XSTDFILL73_1821 VDD VSS sg13g2_FILL8
XSTDFILL73_1829 VDD VSS sg13g2_FILL8
XSTDFILL73_1837 VDD VSS sg13g2_FILL8
XSTDFILL73_1845 VDD VSS sg13g2_FILL8
XSTDFILL73_1853 VDD VSS sg13g2_FILL8
XSTDFILL73_1861 VDD VSS sg13g2_FILL8
XSTDFILL73_1869 VDD VSS sg13g2_FILL8
XSTDFILL73_1877 VDD VSS sg13g2_FILL8
XSTDFILL73_1885 VDD VSS sg13g2_FILL8
XSTDFILL73_1893 VDD VSS sg13g2_FILL8
XSTDFILL73_1901 VDD VSS sg13g2_FILL8
XSTDFILL73_1909 VDD VSS sg13g2_FILL8
XSTDFILL73_1917 VDD VSS sg13g2_FILL8
XSTDFILL73_1925 VDD VSS sg13g2_FILL8
XSTDFILL73_1933 VDD VSS sg13g2_FILL8
XSTDFILL73_1941 VDD VSS sg13g2_FILL8
XSTDFILL73_1949 VDD VSS sg13g2_FILL8
XSTDFILL73_1957 VDD VSS sg13g2_FILL8
XSTDFILL73_1965 VDD VSS sg13g2_FILL8
XSTDFILL73_1973 VDD VSS sg13g2_FILL8
XSTDFILL73_1981 VDD VSS sg13g2_FILL8
XSTDFILL73_1989 VDD VSS sg13g2_FILL8
XSTDFILL73_1997 VDD VSS sg13g2_FILL8
XSTDFILL73_2005 VDD VSS sg13g2_FILL8
XSTDFILL73_2013 VDD VSS sg13g2_FILL8
XSTDFILL73_2021 VDD VSS sg13g2_FILL8
XSTDFILL73_2029 VDD VSS sg13g2_FILL8
XSTDFILL73_2037 VDD VSS sg13g2_FILL8
XSTDFILL73_2045 VDD VSS sg13g2_FILL8
XSTDFILL73_2053 VDD VSS sg13g2_FILL8
XSTDFILL73_2061 VDD VSS sg13g2_FILL8
XSTDFILL73_2069 VDD VSS sg13g2_FILL8
XSTDFILL73_2077 VDD VSS sg13g2_FILL8
XSTDFILL73_2085 VDD VSS sg13g2_FILL8
XSTDFILL73_2093 VDD VSS sg13g2_FILL8
XSTDFILL73_2101 VDD VSS sg13g2_FILL8
XSTDFILL73_2109 VDD VSS sg13g2_FILL8
XSTDFILL73_2117 VDD VSS sg13g2_FILL8
XSTDFILL73_2125 VDD VSS sg13g2_FILL8
XSTDFILL73_2133 VDD VSS sg13g2_FILL8
XSTDFILL73_2141 VDD VSS sg13g2_FILL8
XSTDFILL73_2149 VDD VSS sg13g2_FILL4
XSTDFILL73_2153 VDD VSS sg13g2_FILL1
XSTDFILL74_0 VDD VSS sg13g2_FILL8
XSTDFILL74_8 VDD VSS sg13g2_FILL8
XSTDFILL74_16 VDD VSS sg13g2_FILL8
XSTDFILL74_24 VDD VSS sg13g2_FILL8
XSTDFILL74_32 VDD VSS sg13g2_FILL8
XSTDFILL74_40 VDD VSS sg13g2_FILL8
XSTDFILL74_48 VDD VSS sg13g2_FILL8
XSTDFILL74_56 VDD VSS sg13g2_FILL8
XSTDFILL74_64 VDD VSS sg13g2_FILL8
XSTDFILL74_72 VDD VSS sg13g2_FILL8
XSTDFILL74_80 VDD VSS sg13g2_FILL8
XSTDFILL74_88 VDD VSS sg13g2_FILL8
XSTDFILL74_96 VDD VSS sg13g2_FILL8
XSTDFILL74_104 VDD VSS sg13g2_FILL8
XSTDFILL74_112 VDD VSS sg13g2_FILL8
XSTDFILL74_120 VDD VSS sg13g2_FILL8
XSTDFILL74_128 VDD VSS sg13g2_FILL4
XSTDFILL74_1085 VDD VSS sg13g2_FILL8
XSTDFILL74_1093 VDD VSS sg13g2_FILL8
XSTDFILL74_1101 VDD VSS sg13g2_FILL8
XSTDFILL74_1109 VDD VSS sg13g2_FILL8
XSTDFILL74_1117 VDD VSS sg13g2_FILL8
XSTDFILL74_1125 VDD VSS sg13g2_FILL8
XSTDFILL74_1133 VDD VSS sg13g2_FILL8
XSTDFILL74_1141 VDD VSS sg13g2_FILL8
XSTDFILL74_1149 VDD VSS sg13g2_FILL8
XSTDFILL74_1157 VDD VSS sg13g2_FILL8
XSTDFILL74_1165 VDD VSS sg13g2_FILL8
XSTDFILL74_1173 VDD VSS sg13g2_FILL8
XSTDFILL74_1181 VDD VSS sg13g2_FILL8
XSTDFILL74_1189 VDD VSS sg13g2_FILL8
XSTDFILL74_1197 VDD VSS sg13g2_FILL8
XSTDFILL74_1205 VDD VSS sg13g2_FILL8
XSTDFILL74_1213 VDD VSS sg13g2_FILL8
XSTDFILL74_1221 VDD VSS sg13g2_FILL8
XSTDFILL74_1229 VDD VSS sg13g2_FILL8
XSTDFILL74_1237 VDD VSS sg13g2_FILL8
XSTDFILL74_1245 VDD VSS sg13g2_FILL8
XSTDFILL74_1253 VDD VSS sg13g2_FILL8
XSTDFILL74_1261 VDD VSS sg13g2_FILL8
XSTDFILL74_1269 VDD VSS sg13g2_FILL8
XSTDFILL74_1277 VDD VSS sg13g2_FILL8
XSTDFILL74_1285 VDD VSS sg13g2_FILL8
XSTDFILL74_1293 VDD VSS sg13g2_FILL8
XSTDFILL74_1301 VDD VSS sg13g2_FILL8
XSTDFILL74_1309 VDD VSS sg13g2_FILL8
XSTDFILL74_1317 VDD VSS sg13g2_FILL8
XSTDFILL74_1325 VDD VSS sg13g2_FILL8
XSTDFILL74_1333 VDD VSS sg13g2_FILL8
XSTDFILL74_1341 VDD VSS sg13g2_FILL8
XSTDFILL74_1349 VDD VSS sg13g2_FILL8
XSTDFILL74_1357 VDD VSS sg13g2_FILL8
XSTDFILL74_1365 VDD VSS sg13g2_FILL8
XSTDFILL74_1373 VDD VSS sg13g2_FILL8
XSTDFILL74_1381 VDD VSS sg13g2_FILL8
XSTDFILL74_1389 VDD VSS sg13g2_FILL8
XSTDFILL74_1397 VDD VSS sg13g2_FILL8
XSTDFILL74_1405 VDD VSS sg13g2_FILL8
XSTDFILL74_1413 VDD VSS sg13g2_FILL8
XSTDFILL74_1421 VDD VSS sg13g2_FILL8
XSTDFILL74_1429 VDD VSS sg13g2_FILL8
XSTDFILL74_1437 VDD VSS sg13g2_FILL8
XSTDFILL74_1445 VDD VSS sg13g2_FILL8
XSTDFILL74_1453 VDD VSS sg13g2_FILL8
XSTDFILL74_1461 VDD VSS sg13g2_FILL8
XSTDFILL74_1469 VDD VSS sg13g2_FILL8
XSTDFILL74_1477 VDD VSS sg13g2_FILL8
XSTDFILL74_1485 VDD VSS sg13g2_FILL8
XSTDFILL74_1493 VDD VSS sg13g2_FILL8
XSTDFILL74_1501 VDD VSS sg13g2_FILL8
XSTDFILL74_1509 VDD VSS sg13g2_FILL8
XSTDFILL74_1517 VDD VSS sg13g2_FILL8
XSTDFILL74_1525 VDD VSS sg13g2_FILL8
XSTDFILL74_1533 VDD VSS sg13g2_FILL8
XSTDFILL74_1541 VDD VSS sg13g2_FILL8
XSTDFILL74_1549 VDD VSS sg13g2_FILL8
XSTDFILL74_1557 VDD VSS sg13g2_FILL8
XSTDFILL74_1565 VDD VSS sg13g2_FILL8
XSTDFILL74_1573 VDD VSS sg13g2_FILL8
XSTDFILL74_1581 VDD VSS sg13g2_FILL8
XSTDFILL74_1589 VDD VSS sg13g2_FILL8
XSTDFILL74_1597 VDD VSS sg13g2_FILL8
XSTDFILL74_1605 VDD VSS sg13g2_FILL8
XSTDFILL74_1613 VDD VSS sg13g2_FILL8
XSTDFILL74_1621 VDD VSS sg13g2_FILL8
XSTDFILL74_1629 VDD VSS sg13g2_FILL8
XSTDFILL74_1637 VDD VSS sg13g2_FILL8
XSTDFILL74_1645 VDD VSS sg13g2_FILL8
XSTDFILL74_1653 VDD VSS sg13g2_FILL8
XSTDFILL74_1661 VDD VSS sg13g2_FILL8
XSTDFILL74_1669 VDD VSS sg13g2_FILL8
XSTDFILL74_1677 VDD VSS sg13g2_FILL8
XSTDFILL74_1685 VDD VSS sg13g2_FILL8
XSTDFILL74_1693 VDD VSS sg13g2_FILL8
XSTDFILL74_1701 VDD VSS sg13g2_FILL8
XSTDFILL74_1709 VDD VSS sg13g2_FILL8
XSTDFILL74_1717 VDD VSS sg13g2_FILL8
XSTDFILL74_1725 VDD VSS sg13g2_FILL8
XSTDFILL74_1733 VDD VSS sg13g2_FILL8
XSTDFILL74_1741 VDD VSS sg13g2_FILL8
XSTDFILL74_1749 VDD VSS sg13g2_FILL8
XSTDFILL74_1757 VDD VSS sg13g2_FILL8
XSTDFILL74_1765 VDD VSS sg13g2_FILL8
XSTDFILL74_1773 VDD VSS sg13g2_FILL8
XSTDFILL74_1781 VDD VSS sg13g2_FILL8
XSTDFILL74_1789 VDD VSS sg13g2_FILL8
XSTDFILL74_1797 VDD VSS sg13g2_FILL8
XSTDFILL74_1805 VDD VSS sg13g2_FILL8
XSTDFILL74_1813 VDD VSS sg13g2_FILL8
XSTDFILL74_1821 VDD VSS sg13g2_FILL8
XSTDFILL74_1829 VDD VSS sg13g2_FILL8
XSTDFILL74_1837 VDD VSS sg13g2_FILL8
XSTDFILL74_1845 VDD VSS sg13g2_FILL8
XSTDFILL74_1853 VDD VSS sg13g2_FILL8
XSTDFILL74_1861 VDD VSS sg13g2_FILL8
XSTDFILL74_1869 VDD VSS sg13g2_FILL8
XSTDFILL74_1877 VDD VSS sg13g2_FILL8
XSTDFILL74_1885 VDD VSS sg13g2_FILL8
XSTDFILL74_1893 VDD VSS sg13g2_FILL8
XSTDFILL74_1901 VDD VSS sg13g2_FILL8
XSTDFILL74_1909 VDD VSS sg13g2_FILL8
XSTDFILL74_1917 VDD VSS sg13g2_FILL8
XSTDFILL74_1925 VDD VSS sg13g2_FILL8
XSTDFILL74_1933 VDD VSS sg13g2_FILL8
XSTDFILL74_1941 VDD VSS sg13g2_FILL8
XSTDFILL74_1949 VDD VSS sg13g2_FILL8
XSTDFILL74_1957 VDD VSS sg13g2_FILL8
XSTDFILL74_1965 VDD VSS sg13g2_FILL8
XSTDFILL74_1973 VDD VSS sg13g2_FILL8
XSTDFILL74_1981 VDD VSS sg13g2_FILL8
XSTDFILL74_1989 VDD VSS sg13g2_FILL8
XSTDFILL74_1997 VDD VSS sg13g2_FILL8
XSTDFILL74_2005 VDD VSS sg13g2_FILL8
XSTDFILL74_2013 VDD VSS sg13g2_FILL8
XSTDFILL74_2021 VDD VSS sg13g2_FILL8
XSTDFILL74_2029 VDD VSS sg13g2_FILL8
XSTDFILL74_2037 VDD VSS sg13g2_FILL8
XSTDFILL74_2045 VDD VSS sg13g2_FILL8
XSTDFILL74_2053 VDD VSS sg13g2_FILL8
XSTDFILL74_2061 VDD VSS sg13g2_FILL8
XSTDFILL74_2069 VDD VSS sg13g2_FILL8
XSTDFILL74_2077 VDD VSS sg13g2_FILL8
XSTDFILL74_2085 VDD VSS sg13g2_FILL8
XSTDFILL74_2093 VDD VSS sg13g2_FILL8
XSTDFILL74_2101 VDD VSS sg13g2_FILL8
XSTDFILL74_2109 VDD VSS sg13g2_FILL8
XSTDFILL74_2117 VDD VSS sg13g2_FILL8
XSTDFILL74_2125 VDD VSS sg13g2_FILL8
XSTDFILL74_2133 VDD VSS sg13g2_FILL8
XSTDFILL74_2141 VDD VSS sg13g2_FILL8
XSTDFILL74_2149 VDD VSS sg13g2_FILL4
XSTDFILL74_2153 VDD VSS sg13g2_FILL1
XSTDFILL75_0 VDD VSS sg13g2_FILL8
XSTDFILL75_8 VDD VSS sg13g2_FILL8
XSTDFILL75_16 VDD VSS sg13g2_FILL8
XSTDFILL75_24 VDD VSS sg13g2_FILL8
XSTDFILL75_32 VDD VSS sg13g2_FILL8
XSTDFILL75_40 VDD VSS sg13g2_FILL8
XSTDFILL75_48 VDD VSS sg13g2_FILL8
XSTDFILL75_56 VDD VSS sg13g2_FILL8
XSTDFILL75_64 VDD VSS sg13g2_FILL8
XSTDFILL75_72 VDD VSS sg13g2_FILL8
XSTDFILL75_80 VDD VSS sg13g2_FILL8
XSTDFILL75_88 VDD VSS sg13g2_FILL8
XSTDFILL75_96 VDD VSS sg13g2_FILL8
XSTDFILL75_104 VDD VSS sg13g2_FILL8
XSTDFILL75_112 VDD VSS sg13g2_FILL8
XSTDFILL75_120 VDD VSS sg13g2_FILL8
XSTDFILL75_128 VDD VSS sg13g2_FILL4
XSTDFILL75_1085 VDD VSS sg13g2_FILL8
XSTDFILL75_1093 VDD VSS sg13g2_FILL8
XSTDFILL75_1101 VDD VSS sg13g2_FILL8
XSTDFILL75_1109 VDD VSS sg13g2_FILL8
XSTDFILL75_1117 VDD VSS sg13g2_FILL8
XSTDFILL75_1125 VDD VSS sg13g2_FILL8
XSTDFILL75_1133 VDD VSS sg13g2_FILL8
XSTDFILL75_1141 VDD VSS sg13g2_FILL8
XSTDFILL75_1149 VDD VSS sg13g2_FILL8
XSTDFILL75_1157 VDD VSS sg13g2_FILL8
XSTDFILL75_1165 VDD VSS sg13g2_FILL8
XSTDFILL75_1173 VDD VSS sg13g2_FILL8
XSTDFILL75_1181 VDD VSS sg13g2_FILL8
XSTDFILL75_1189 VDD VSS sg13g2_FILL8
XSTDFILL75_1197 VDD VSS sg13g2_FILL8
XSTDFILL75_1205 VDD VSS sg13g2_FILL8
XSTDFILL75_1213 VDD VSS sg13g2_FILL8
XSTDFILL75_1221 VDD VSS sg13g2_FILL8
XSTDFILL75_1229 VDD VSS sg13g2_FILL8
XSTDFILL75_1237 VDD VSS sg13g2_FILL8
XSTDFILL75_1245 VDD VSS sg13g2_FILL8
XSTDFILL75_1253 VDD VSS sg13g2_FILL8
XSTDFILL75_1261 VDD VSS sg13g2_FILL8
XSTDFILL75_1269 VDD VSS sg13g2_FILL8
XSTDFILL75_1277 VDD VSS sg13g2_FILL8
XSTDFILL75_1285 VDD VSS sg13g2_FILL8
XSTDFILL75_1293 VDD VSS sg13g2_FILL8
XSTDFILL75_1301 VDD VSS sg13g2_FILL8
XSTDFILL75_1309 VDD VSS sg13g2_FILL8
XSTDFILL75_1317 VDD VSS sg13g2_FILL8
XSTDFILL75_1325 VDD VSS sg13g2_FILL8
XSTDFILL75_1333 VDD VSS sg13g2_FILL8
XSTDFILL75_1341 VDD VSS sg13g2_FILL8
XSTDFILL75_1349 VDD VSS sg13g2_FILL8
XSTDFILL75_1357 VDD VSS sg13g2_FILL8
XSTDFILL75_1365 VDD VSS sg13g2_FILL8
XSTDFILL75_1373 VDD VSS sg13g2_FILL8
XSTDFILL75_1381 VDD VSS sg13g2_FILL8
XSTDFILL75_1389 VDD VSS sg13g2_FILL8
XSTDFILL75_1397 VDD VSS sg13g2_FILL8
XSTDFILL75_1405 VDD VSS sg13g2_FILL8
XSTDFILL75_1413 VDD VSS sg13g2_FILL8
XSTDFILL75_1421 VDD VSS sg13g2_FILL8
XSTDFILL75_1429 VDD VSS sg13g2_FILL8
XSTDFILL75_1437 VDD VSS sg13g2_FILL8
XSTDFILL75_1445 VDD VSS sg13g2_FILL8
XSTDFILL75_1453 VDD VSS sg13g2_FILL8
XSTDFILL75_1461 VDD VSS sg13g2_FILL8
XSTDFILL75_1469 VDD VSS sg13g2_FILL8
XSTDFILL75_1477 VDD VSS sg13g2_FILL8
XSTDFILL75_1485 VDD VSS sg13g2_FILL8
XSTDFILL75_1493 VDD VSS sg13g2_FILL8
XSTDFILL75_1501 VDD VSS sg13g2_FILL8
XSTDFILL75_1509 VDD VSS sg13g2_FILL8
XSTDFILL75_1517 VDD VSS sg13g2_FILL8
XSTDFILL75_1525 VDD VSS sg13g2_FILL8
XSTDFILL75_1533 VDD VSS sg13g2_FILL8
XSTDFILL75_1541 VDD VSS sg13g2_FILL8
XSTDFILL75_1549 VDD VSS sg13g2_FILL8
XSTDFILL75_1557 VDD VSS sg13g2_FILL8
XSTDFILL75_1565 VDD VSS sg13g2_FILL8
XSTDFILL75_1573 VDD VSS sg13g2_FILL8
XSTDFILL75_1581 VDD VSS sg13g2_FILL8
XSTDFILL75_1589 VDD VSS sg13g2_FILL8
XSTDFILL75_1597 VDD VSS sg13g2_FILL8
XSTDFILL75_1605 VDD VSS sg13g2_FILL8
XSTDFILL75_1613 VDD VSS sg13g2_FILL8
XSTDFILL75_1621 VDD VSS sg13g2_FILL8
XSTDFILL75_1629 VDD VSS sg13g2_FILL8
XSTDFILL75_1637 VDD VSS sg13g2_FILL8
XSTDFILL75_1645 VDD VSS sg13g2_FILL8
XSTDFILL75_1653 VDD VSS sg13g2_FILL8
XSTDFILL75_1661 VDD VSS sg13g2_FILL8
XSTDFILL75_1669 VDD VSS sg13g2_FILL8
XSTDFILL75_1677 VDD VSS sg13g2_FILL8
XSTDFILL75_1685 VDD VSS sg13g2_FILL8
XSTDFILL75_1693 VDD VSS sg13g2_FILL8
XSTDFILL75_1701 VDD VSS sg13g2_FILL8
XSTDFILL75_1709 VDD VSS sg13g2_FILL8
XSTDFILL75_1717 VDD VSS sg13g2_FILL8
XSTDFILL75_1725 VDD VSS sg13g2_FILL8
XSTDFILL75_1733 VDD VSS sg13g2_FILL8
XSTDFILL75_1741 VDD VSS sg13g2_FILL8
XSTDFILL75_1749 VDD VSS sg13g2_FILL8
XSTDFILL75_1757 VDD VSS sg13g2_FILL8
XSTDFILL75_1765 VDD VSS sg13g2_FILL8
XSTDFILL75_1773 VDD VSS sg13g2_FILL8
XSTDFILL75_1781 VDD VSS sg13g2_FILL8
XSTDFILL75_1789 VDD VSS sg13g2_FILL8
XSTDFILL75_1797 VDD VSS sg13g2_FILL8
XSTDFILL75_1805 VDD VSS sg13g2_FILL8
XSTDFILL75_1813 VDD VSS sg13g2_FILL8
XSTDFILL75_1821 VDD VSS sg13g2_FILL8
XSTDFILL75_1829 VDD VSS sg13g2_FILL8
XSTDFILL75_1837 VDD VSS sg13g2_FILL8
XSTDFILL75_1845 VDD VSS sg13g2_FILL8
XSTDFILL75_1853 VDD VSS sg13g2_FILL8
XSTDFILL75_1861 VDD VSS sg13g2_FILL8
XSTDFILL75_1869 VDD VSS sg13g2_FILL8
XSTDFILL75_1877 VDD VSS sg13g2_FILL8
XSTDFILL75_1885 VDD VSS sg13g2_FILL8
XSTDFILL75_1893 VDD VSS sg13g2_FILL8
XSTDFILL75_1901 VDD VSS sg13g2_FILL8
XSTDFILL75_1909 VDD VSS sg13g2_FILL8
XSTDFILL75_1917 VDD VSS sg13g2_FILL8
XSTDFILL75_1925 VDD VSS sg13g2_FILL8
XSTDFILL75_1933 VDD VSS sg13g2_FILL8
XSTDFILL75_1941 VDD VSS sg13g2_FILL8
XSTDFILL75_1949 VDD VSS sg13g2_FILL8
XSTDFILL75_1957 VDD VSS sg13g2_FILL8
XSTDFILL75_1965 VDD VSS sg13g2_FILL8
XSTDFILL75_1973 VDD VSS sg13g2_FILL8
XSTDFILL75_1981 VDD VSS sg13g2_FILL8
XSTDFILL75_1989 VDD VSS sg13g2_FILL8
XSTDFILL75_1997 VDD VSS sg13g2_FILL8
XSTDFILL75_2005 VDD VSS sg13g2_FILL8
XSTDFILL75_2013 VDD VSS sg13g2_FILL8
XSTDFILL75_2021 VDD VSS sg13g2_FILL8
XSTDFILL75_2029 VDD VSS sg13g2_FILL8
XSTDFILL75_2037 VDD VSS sg13g2_FILL8
XSTDFILL75_2045 VDD VSS sg13g2_FILL8
XSTDFILL75_2053 VDD VSS sg13g2_FILL8
XSTDFILL75_2061 VDD VSS sg13g2_FILL8
XSTDFILL75_2069 VDD VSS sg13g2_FILL8
XSTDFILL75_2077 VDD VSS sg13g2_FILL8
XSTDFILL75_2085 VDD VSS sg13g2_FILL8
XSTDFILL75_2093 VDD VSS sg13g2_FILL8
XSTDFILL75_2101 VDD VSS sg13g2_FILL8
XSTDFILL75_2109 VDD VSS sg13g2_FILL8
XSTDFILL75_2117 VDD VSS sg13g2_FILL8
XSTDFILL75_2125 VDD VSS sg13g2_FILL8
XSTDFILL75_2133 VDD VSS sg13g2_FILL8
XSTDFILL75_2141 VDD VSS sg13g2_FILL8
XSTDFILL75_2149 VDD VSS sg13g2_FILL4
XSTDFILL75_2153 VDD VSS sg13g2_FILL1
XSTDFILL76_0 VDD VSS sg13g2_FILL8
XSTDFILL76_8 VDD VSS sg13g2_FILL8
XSTDFILL76_16 VDD VSS sg13g2_FILL8
XSTDFILL76_24 VDD VSS sg13g2_FILL8
XSTDFILL76_32 VDD VSS sg13g2_FILL8
XSTDFILL76_40 VDD VSS sg13g2_FILL8
XSTDFILL76_48 VDD VSS sg13g2_FILL8
XSTDFILL76_56 VDD VSS sg13g2_FILL8
XSTDFILL76_64 VDD VSS sg13g2_FILL8
XSTDFILL76_72 VDD VSS sg13g2_FILL8
XSTDFILL76_80 VDD VSS sg13g2_FILL8
XSTDFILL76_88 VDD VSS sg13g2_FILL8
XSTDFILL76_96 VDD VSS sg13g2_FILL8
XSTDFILL76_104 VDD VSS sg13g2_FILL8
XSTDFILL76_112 VDD VSS sg13g2_FILL8
XSTDFILL76_120 VDD VSS sg13g2_FILL8
XSTDFILL76_128 VDD VSS sg13g2_FILL4
XSTDFILL76_1085 VDD VSS sg13g2_FILL8
XSTDFILL76_1093 VDD VSS sg13g2_FILL8
XSTDFILL76_1101 VDD VSS sg13g2_FILL8
XSTDFILL76_1109 VDD VSS sg13g2_FILL8
XSTDFILL76_1117 VDD VSS sg13g2_FILL8
XSTDFILL76_1125 VDD VSS sg13g2_FILL8
XSTDFILL76_1133 VDD VSS sg13g2_FILL8
XSTDFILL76_1141 VDD VSS sg13g2_FILL8
XSTDFILL76_1149 VDD VSS sg13g2_FILL8
XSTDFILL76_1157 VDD VSS sg13g2_FILL8
XSTDFILL76_1165 VDD VSS sg13g2_FILL8
XSTDFILL76_1173 VDD VSS sg13g2_FILL8
XSTDFILL76_1181 VDD VSS sg13g2_FILL8
XSTDFILL76_1189 VDD VSS sg13g2_FILL8
XSTDFILL76_1197 VDD VSS sg13g2_FILL8
XSTDFILL76_1205 VDD VSS sg13g2_FILL8
XSTDFILL76_1213 VDD VSS sg13g2_FILL8
XSTDFILL76_1221 VDD VSS sg13g2_FILL8
XSTDFILL76_1229 VDD VSS sg13g2_FILL8
XSTDFILL76_1237 VDD VSS sg13g2_FILL8
XSTDFILL76_1245 VDD VSS sg13g2_FILL8
XSTDFILL76_1253 VDD VSS sg13g2_FILL8
XSTDFILL76_1261 VDD VSS sg13g2_FILL8
XSTDFILL76_1269 VDD VSS sg13g2_FILL8
XSTDFILL76_1277 VDD VSS sg13g2_FILL8
XSTDFILL76_1285 VDD VSS sg13g2_FILL8
XSTDFILL76_1293 VDD VSS sg13g2_FILL8
XSTDFILL76_1301 VDD VSS sg13g2_FILL8
XSTDFILL76_1309 VDD VSS sg13g2_FILL8
XSTDFILL76_1317 VDD VSS sg13g2_FILL8
XSTDFILL76_1325 VDD VSS sg13g2_FILL8
XSTDFILL76_1333 VDD VSS sg13g2_FILL8
XSTDFILL76_1341 VDD VSS sg13g2_FILL8
XSTDFILL76_1349 VDD VSS sg13g2_FILL8
XSTDFILL76_1357 VDD VSS sg13g2_FILL8
XSTDFILL76_1365 VDD VSS sg13g2_FILL8
XSTDFILL76_1373 VDD VSS sg13g2_FILL8
XSTDFILL76_1381 VDD VSS sg13g2_FILL8
XSTDFILL76_1389 VDD VSS sg13g2_FILL8
XSTDFILL76_1397 VDD VSS sg13g2_FILL8
XSTDFILL76_1405 VDD VSS sg13g2_FILL8
XSTDFILL76_1413 VDD VSS sg13g2_FILL8
XSTDFILL76_1421 VDD VSS sg13g2_FILL8
XSTDFILL76_1429 VDD VSS sg13g2_FILL8
XSTDFILL76_1437 VDD VSS sg13g2_FILL8
XSTDFILL76_1445 VDD VSS sg13g2_FILL8
XSTDFILL76_1453 VDD VSS sg13g2_FILL8
XSTDFILL76_1461 VDD VSS sg13g2_FILL8
XSTDFILL76_1469 VDD VSS sg13g2_FILL8
XSTDFILL76_1477 VDD VSS sg13g2_FILL8
XSTDFILL76_1485 VDD VSS sg13g2_FILL8
XSTDFILL76_1493 VDD VSS sg13g2_FILL8
XSTDFILL76_1501 VDD VSS sg13g2_FILL8
XSTDFILL76_1509 VDD VSS sg13g2_FILL8
XSTDFILL76_1517 VDD VSS sg13g2_FILL8
XSTDFILL76_1525 VDD VSS sg13g2_FILL8
XSTDFILL76_1533 VDD VSS sg13g2_FILL8
XSTDFILL76_1541 VDD VSS sg13g2_FILL8
XSTDFILL76_1549 VDD VSS sg13g2_FILL8
XSTDFILL76_1557 VDD VSS sg13g2_FILL8
XSTDFILL76_1565 VDD VSS sg13g2_FILL8
XSTDFILL76_1573 VDD VSS sg13g2_FILL8
XSTDFILL76_1581 VDD VSS sg13g2_FILL8
XSTDFILL76_1589 VDD VSS sg13g2_FILL8
XSTDFILL76_1597 VDD VSS sg13g2_FILL8
XSTDFILL76_1605 VDD VSS sg13g2_FILL8
XSTDFILL76_1613 VDD VSS sg13g2_FILL8
XSTDFILL76_1621 VDD VSS sg13g2_FILL8
XSTDFILL76_1629 VDD VSS sg13g2_FILL8
XSTDFILL76_1637 VDD VSS sg13g2_FILL8
XSTDFILL76_1645 VDD VSS sg13g2_FILL8
XSTDFILL76_1653 VDD VSS sg13g2_FILL8
XSTDFILL76_1661 VDD VSS sg13g2_FILL8
XSTDFILL76_1669 VDD VSS sg13g2_FILL8
XSTDFILL76_1677 VDD VSS sg13g2_FILL8
XSTDFILL76_1685 VDD VSS sg13g2_FILL8
XSTDFILL76_1693 VDD VSS sg13g2_FILL8
XSTDFILL76_1701 VDD VSS sg13g2_FILL8
XSTDFILL76_1709 VDD VSS sg13g2_FILL8
XSTDFILL76_1717 VDD VSS sg13g2_FILL8
XSTDFILL76_1725 VDD VSS sg13g2_FILL8
XSTDFILL76_1733 VDD VSS sg13g2_FILL8
XSTDFILL76_1741 VDD VSS sg13g2_FILL8
XSTDFILL76_1749 VDD VSS sg13g2_FILL8
XSTDFILL76_1757 VDD VSS sg13g2_FILL8
XSTDFILL76_1765 VDD VSS sg13g2_FILL8
XSTDFILL76_1773 VDD VSS sg13g2_FILL8
XSTDFILL76_1781 VDD VSS sg13g2_FILL8
XSTDFILL76_1789 VDD VSS sg13g2_FILL8
XSTDFILL76_1797 VDD VSS sg13g2_FILL8
XSTDFILL76_1805 VDD VSS sg13g2_FILL8
XSTDFILL76_1813 VDD VSS sg13g2_FILL8
XSTDFILL76_1821 VDD VSS sg13g2_FILL8
XSTDFILL76_1829 VDD VSS sg13g2_FILL8
XSTDFILL76_1837 VDD VSS sg13g2_FILL8
XSTDFILL76_1845 VDD VSS sg13g2_FILL8
XSTDFILL76_1853 VDD VSS sg13g2_FILL8
XSTDFILL76_1861 VDD VSS sg13g2_FILL8
XSTDFILL76_1869 VDD VSS sg13g2_FILL8
XSTDFILL76_1877 VDD VSS sg13g2_FILL8
XSTDFILL76_1885 VDD VSS sg13g2_FILL8
XSTDFILL76_1893 VDD VSS sg13g2_FILL8
XSTDFILL76_1901 VDD VSS sg13g2_FILL8
XSTDFILL76_1909 VDD VSS sg13g2_FILL8
XSTDFILL76_1917 VDD VSS sg13g2_FILL8
XSTDFILL76_1925 VDD VSS sg13g2_FILL8
XSTDFILL76_1933 VDD VSS sg13g2_FILL8
XSTDFILL76_1941 VDD VSS sg13g2_FILL8
XSTDFILL76_1949 VDD VSS sg13g2_FILL8
XSTDFILL76_1957 VDD VSS sg13g2_FILL8
XSTDFILL76_1965 VDD VSS sg13g2_FILL8
XSTDFILL76_1973 VDD VSS sg13g2_FILL8
XSTDFILL76_1981 VDD VSS sg13g2_FILL8
XSTDFILL76_1989 VDD VSS sg13g2_FILL8
XSTDFILL76_1997 VDD VSS sg13g2_FILL8
XSTDFILL76_2005 VDD VSS sg13g2_FILL8
XSTDFILL76_2013 VDD VSS sg13g2_FILL8
XSTDFILL76_2021 VDD VSS sg13g2_FILL8
XSTDFILL76_2029 VDD VSS sg13g2_FILL8
XSTDFILL76_2037 VDD VSS sg13g2_FILL8
XSTDFILL76_2045 VDD VSS sg13g2_FILL8
XSTDFILL76_2053 VDD VSS sg13g2_FILL8
XSTDFILL76_2061 VDD VSS sg13g2_FILL8
XSTDFILL76_2069 VDD VSS sg13g2_FILL8
XSTDFILL76_2077 VDD VSS sg13g2_FILL8
XSTDFILL76_2085 VDD VSS sg13g2_FILL8
XSTDFILL76_2093 VDD VSS sg13g2_FILL8
XSTDFILL76_2101 VDD VSS sg13g2_FILL8
XSTDFILL76_2109 VDD VSS sg13g2_FILL8
XSTDFILL76_2117 VDD VSS sg13g2_FILL8
XSTDFILL76_2125 VDD VSS sg13g2_FILL8
XSTDFILL76_2133 VDD VSS sg13g2_FILL8
XSTDFILL76_2141 VDD VSS sg13g2_FILL8
XSTDFILL76_2149 VDD VSS sg13g2_FILL4
XSTDFILL76_2153 VDD VSS sg13g2_FILL1
XSTDFILL77_0 VDD VSS sg13g2_FILL8
XSTDFILL77_8 VDD VSS sg13g2_FILL8
XSTDFILL77_16 VDD VSS sg13g2_FILL8
XSTDFILL77_24 VDD VSS sg13g2_FILL8
XSTDFILL77_32 VDD VSS sg13g2_FILL8
XSTDFILL77_40 VDD VSS sg13g2_FILL8
XSTDFILL77_48 VDD VSS sg13g2_FILL8
XSTDFILL77_56 VDD VSS sg13g2_FILL8
XSTDFILL77_64 VDD VSS sg13g2_FILL8
XSTDFILL77_72 VDD VSS sg13g2_FILL8
XSTDFILL77_80 VDD VSS sg13g2_FILL8
XSTDFILL77_88 VDD VSS sg13g2_FILL8
XSTDFILL77_96 VDD VSS sg13g2_FILL8
XSTDFILL77_104 VDD VSS sg13g2_FILL8
XSTDFILL77_112 VDD VSS sg13g2_FILL8
XSTDFILL77_120 VDD VSS sg13g2_FILL8
XSTDFILL77_128 VDD VSS sg13g2_FILL4
XSTDFILL77_1085 VDD VSS sg13g2_FILL8
XSTDFILL77_1093 VDD VSS sg13g2_FILL8
XSTDFILL77_1101 VDD VSS sg13g2_FILL8
XSTDFILL77_1109 VDD VSS sg13g2_FILL8
XSTDFILL77_1117 VDD VSS sg13g2_FILL8
XSTDFILL77_1125 VDD VSS sg13g2_FILL8
XSTDFILL77_1133 VDD VSS sg13g2_FILL8
XSTDFILL77_1141 VDD VSS sg13g2_FILL8
XSTDFILL77_1149 VDD VSS sg13g2_FILL8
XSTDFILL77_1157 VDD VSS sg13g2_FILL8
XSTDFILL77_1165 VDD VSS sg13g2_FILL8
XSTDFILL77_1173 VDD VSS sg13g2_FILL8
XSTDFILL77_1181 VDD VSS sg13g2_FILL8
XSTDFILL77_1189 VDD VSS sg13g2_FILL8
XSTDFILL77_1197 VDD VSS sg13g2_FILL8
XSTDFILL77_1205 VDD VSS sg13g2_FILL8
XSTDFILL77_1213 VDD VSS sg13g2_FILL8
XSTDFILL77_1221 VDD VSS sg13g2_FILL8
XSTDFILL77_1229 VDD VSS sg13g2_FILL8
XSTDFILL77_1237 VDD VSS sg13g2_FILL8
XSTDFILL77_1245 VDD VSS sg13g2_FILL8
XSTDFILL77_1253 VDD VSS sg13g2_FILL8
XSTDFILL77_1261 VDD VSS sg13g2_FILL8
XSTDFILL77_1269 VDD VSS sg13g2_FILL8
XSTDFILL77_1277 VDD VSS sg13g2_FILL8
XSTDFILL77_1285 VDD VSS sg13g2_FILL8
XSTDFILL77_1293 VDD VSS sg13g2_FILL8
XSTDFILL77_1301 VDD VSS sg13g2_FILL8
XSTDFILL77_1309 VDD VSS sg13g2_FILL8
XSTDFILL77_1317 VDD VSS sg13g2_FILL8
XSTDFILL77_1325 VDD VSS sg13g2_FILL8
XSTDFILL77_1333 VDD VSS sg13g2_FILL8
XSTDFILL77_1341 VDD VSS sg13g2_FILL8
XSTDFILL77_1349 VDD VSS sg13g2_FILL8
XSTDFILL77_1357 VDD VSS sg13g2_FILL8
XSTDFILL77_1365 VDD VSS sg13g2_FILL8
XSTDFILL77_1373 VDD VSS sg13g2_FILL8
XSTDFILL77_1381 VDD VSS sg13g2_FILL8
XSTDFILL77_1389 VDD VSS sg13g2_FILL8
XSTDFILL77_1397 VDD VSS sg13g2_FILL8
XSTDFILL77_1405 VDD VSS sg13g2_FILL8
XSTDFILL77_1413 VDD VSS sg13g2_FILL8
XSTDFILL77_1421 VDD VSS sg13g2_FILL8
XSTDFILL77_1429 VDD VSS sg13g2_FILL8
XSTDFILL77_1437 VDD VSS sg13g2_FILL8
XSTDFILL77_1445 VDD VSS sg13g2_FILL8
XSTDFILL77_1453 VDD VSS sg13g2_FILL8
XSTDFILL77_1461 VDD VSS sg13g2_FILL8
XSTDFILL77_1469 VDD VSS sg13g2_FILL8
XSTDFILL77_1477 VDD VSS sg13g2_FILL8
XSTDFILL77_1485 VDD VSS sg13g2_FILL8
XSTDFILL77_1493 VDD VSS sg13g2_FILL8
XSTDFILL77_1501 VDD VSS sg13g2_FILL8
XSTDFILL77_1509 VDD VSS sg13g2_FILL8
XSTDFILL77_1517 VDD VSS sg13g2_FILL8
XSTDFILL77_1525 VDD VSS sg13g2_FILL8
XSTDFILL77_1533 VDD VSS sg13g2_FILL8
XSTDFILL77_1541 VDD VSS sg13g2_FILL8
XSTDFILL77_1549 VDD VSS sg13g2_FILL8
XSTDFILL77_1557 VDD VSS sg13g2_FILL8
XSTDFILL77_1565 VDD VSS sg13g2_FILL8
XSTDFILL77_1573 VDD VSS sg13g2_FILL8
XSTDFILL77_1581 VDD VSS sg13g2_FILL8
XSTDFILL77_1589 VDD VSS sg13g2_FILL8
XSTDFILL77_1597 VDD VSS sg13g2_FILL8
XSTDFILL77_1605 VDD VSS sg13g2_FILL8
XSTDFILL77_1613 VDD VSS sg13g2_FILL8
XSTDFILL77_1621 VDD VSS sg13g2_FILL8
XSTDFILL77_1629 VDD VSS sg13g2_FILL8
XSTDFILL77_1637 VDD VSS sg13g2_FILL8
XSTDFILL77_1645 VDD VSS sg13g2_FILL8
XSTDFILL77_1653 VDD VSS sg13g2_FILL8
XSTDFILL77_1661 VDD VSS sg13g2_FILL8
XSTDFILL77_1669 VDD VSS sg13g2_FILL8
XSTDFILL77_1677 VDD VSS sg13g2_FILL8
XSTDFILL77_1685 VDD VSS sg13g2_FILL8
XSTDFILL77_1693 VDD VSS sg13g2_FILL8
XSTDFILL77_1701 VDD VSS sg13g2_FILL8
XSTDFILL77_1709 VDD VSS sg13g2_FILL8
XSTDFILL77_1717 VDD VSS sg13g2_FILL8
XSTDFILL77_1725 VDD VSS sg13g2_FILL8
XSTDFILL77_1733 VDD VSS sg13g2_FILL8
XSTDFILL77_1741 VDD VSS sg13g2_FILL8
XSTDFILL77_1749 VDD VSS sg13g2_FILL8
XSTDFILL77_1757 VDD VSS sg13g2_FILL8
XSTDFILL77_1765 VDD VSS sg13g2_FILL8
XSTDFILL77_1773 VDD VSS sg13g2_FILL8
XSTDFILL77_1781 VDD VSS sg13g2_FILL8
XSTDFILL77_1789 VDD VSS sg13g2_FILL8
XSTDFILL77_1797 VDD VSS sg13g2_FILL8
XSTDFILL77_1805 VDD VSS sg13g2_FILL8
XSTDFILL77_1813 VDD VSS sg13g2_FILL8
XSTDFILL77_1821 VDD VSS sg13g2_FILL8
XSTDFILL77_1829 VDD VSS sg13g2_FILL8
XSTDFILL77_1837 VDD VSS sg13g2_FILL8
XSTDFILL77_1845 VDD VSS sg13g2_FILL8
XSTDFILL77_1853 VDD VSS sg13g2_FILL8
XSTDFILL77_1861 VDD VSS sg13g2_FILL8
XSTDFILL77_1869 VDD VSS sg13g2_FILL8
XSTDFILL77_1877 VDD VSS sg13g2_FILL8
XSTDFILL77_1885 VDD VSS sg13g2_FILL8
XSTDFILL77_1893 VDD VSS sg13g2_FILL8
XSTDFILL77_1901 VDD VSS sg13g2_FILL8
XSTDFILL77_1909 VDD VSS sg13g2_FILL8
XSTDFILL77_1917 VDD VSS sg13g2_FILL8
XSTDFILL77_1925 VDD VSS sg13g2_FILL8
XSTDFILL77_1933 VDD VSS sg13g2_FILL8
XSTDFILL77_1941 VDD VSS sg13g2_FILL8
XSTDFILL77_1949 VDD VSS sg13g2_FILL8
XSTDFILL77_1957 VDD VSS sg13g2_FILL8
XSTDFILL77_1965 VDD VSS sg13g2_FILL8
XSTDFILL77_1973 VDD VSS sg13g2_FILL8
XSTDFILL77_1981 VDD VSS sg13g2_FILL8
XSTDFILL77_1989 VDD VSS sg13g2_FILL8
XSTDFILL77_1997 VDD VSS sg13g2_FILL8
XSTDFILL77_2005 VDD VSS sg13g2_FILL8
XSTDFILL77_2013 VDD VSS sg13g2_FILL8
XSTDFILL77_2021 VDD VSS sg13g2_FILL8
XSTDFILL77_2029 VDD VSS sg13g2_FILL8
XSTDFILL77_2037 VDD VSS sg13g2_FILL8
XSTDFILL77_2045 VDD VSS sg13g2_FILL8
XSTDFILL77_2053 VDD VSS sg13g2_FILL8
XSTDFILL77_2061 VDD VSS sg13g2_FILL8
XSTDFILL77_2069 VDD VSS sg13g2_FILL8
XSTDFILL77_2077 VDD VSS sg13g2_FILL8
XSTDFILL77_2085 VDD VSS sg13g2_FILL8
XSTDFILL77_2093 VDD VSS sg13g2_FILL8
XSTDFILL77_2101 VDD VSS sg13g2_FILL8
XSTDFILL77_2109 VDD VSS sg13g2_FILL8
XSTDFILL77_2117 VDD VSS sg13g2_FILL8
XSTDFILL77_2125 VDD VSS sg13g2_FILL8
XSTDFILL77_2133 VDD VSS sg13g2_FILL8
XSTDFILL77_2141 VDD VSS sg13g2_FILL8
XSTDFILL77_2149 VDD VSS sg13g2_FILL4
XSTDFILL77_2153 VDD VSS sg13g2_FILL1
XSTDFILL78_0 VDD VSS sg13g2_FILL8
XSTDFILL78_8 VDD VSS sg13g2_FILL8
XSTDFILL78_16 VDD VSS sg13g2_FILL8
XSTDFILL78_24 VDD VSS sg13g2_FILL8
XSTDFILL78_32 VDD VSS sg13g2_FILL8
XSTDFILL78_40 VDD VSS sg13g2_FILL8
XSTDFILL78_48 VDD VSS sg13g2_FILL8
XSTDFILL78_56 VDD VSS sg13g2_FILL8
XSTDFILL78_64 VDD VSS sg13g2_FILL8
XSTDFILL78_72 VDD VSS sg13g2_FILL8
XSTDFILL78_80 VDD VSS sg13g2_FILL8
XSTDFILL78_88 VDD VSS sg13g2_FILL8
XSTDFILL78_96 VDD VSS sg13g2_FILL8
XSTDFILL78_104 VDD VSS sg13g2_FILL8
XSTDFILL78_112 VDD VSS sg13g2_FILL8
XSTDFILL78_120 VDD VSS sg13g2_FILL8
XSTDFILL78_128 VDD VSS sg13g2_FILL4
XSTDFILL78_1085 VDD VSS sg13g2_FILL8
XSTDFILL78_1093 VDD VSS sg13g2_FILL8
XSTDFILL78_1101 VDD VSS sg13g2_FILL8
XSTDFILL78_1109 VDD VSS sg13g2_FILL8
XSTDFILL78_1117 VDD VSS sg13g2_FILL8
XSTDFILL78_1125 VDD VSS sg13g2_FILL8
XSTDFILL78_1133 VDD VSS sg13g2_FILL8
XSTDFILL78_1141 VDD VSS sg13g2_FILL8
XSTDFILL78_1149 VDD VSS sg13g2_FILL8
XSTDFILL78_1157 VDD VSS sg13g2_FILL8
XSTDFILL78_1165 VDD VSS sg13g2_FILL8
XSTDFILL78_1173 VDD VSS sg13g2_FILL8
XSTDFILL78_1181 VDD VSS sg13g2_FILL8
XSTDFILL78_1189 VDD VSS sg13g2_FILL8
XSTDFILL78_1197 VDD VSS sg13g2_FILL8
XSTDFILL78_1205 VDD VSS sg13g2_FILL8
XSTDFILL78_1213 VDD VSS sg13g2_FILL8
XSTDFILL78_1221 VDD VSS sg13g2_FILL8
XSTDFILL78_1229 VDD VSS sg13g2_FILL8
XSTDFILL78_1237 VDD VSS sg13g2_FILL8
XSTDFILL78_1245 VDD VSS sg13g2_FILL8
XSTDFILL78_1253 VDD VSS sg13g2_FILL8
XSTDFILL78_1261 VDD VSS sg13g2_FILL8
XSTDFILL78_1269 VDD VSS sg13g2_FILL8
XSTDFILL78_1277 VDD VSS sg13g2_FILL8
XSTDFILL78_1285 VDD VSS sg13g2_FILL8
XSTDFILL78_1293 VDD VSS sg13g2_FILL8
XSTDFILL78_1301 VDD VSS sg13g2_FILL8
XSTDFILL78_1309 VDD VSS sg13g2_FILL8
XSTDFILL78_1317 VDD VSS sg13g2_FILL8
XSTDFILL78_1325 VDD VSS sg13g2_FILL8
XSTDFILL78_1333 VDD VSS sg13g2_FILL8
XSTDFILL78_1341 VDD VSS sg13g2_FILL8
XSTDFILL78_1349 VDD VSS sg13g2_FILL8
XSTDFILL78_1357 VDD VSS sg13g2_FILL8
XSTDFILL78_1365 VDD VSS sg13g2_FILL8
XSTDFILL78_1373 VDD VSS sg13g2_FILL8
XSTDFILL78_1381 VDD VSS sg13g2_FILL8
XSTDFILL78_1389 VDD VSS sg13g2_FILL8
XSTDFILL78_1397 VDD VSS sg13g2_FILL8
XSTDFILL78_1405 VDD VSS sg13g2_FILL8
XSTDFILL78_1413 VDD VSS sg13g2_FILL8
XSTDFILL78_1421 VDD VSS sg13g2_FILL8
XSTDFILL78_1429 VDD VSS sg13g2_FILL8
XSTDFILL78_1437 VDD VSS sg13g2_FILL8
XSTDFILL78_1445 VDD VSS sg13g2_FILL8
XSTDFILL78_1453 VDD VSS sg13g2_FILL8
XSTDFILL78_1461 VDD VSS sg13g2_FILL8
XSTDFILL78_1469 VDD VSS sg13g2_FILL8
XSTDFILL78_1477 VDD VSS sg13g2_FILL8
XSTDFILL78_1485 VDD VSS sg13g2_FILL8
XSTDFILL78_1493 VDD VSS sg13g2_FILL8
XSTDFILL78_1501 VDD VSS sg13g2_FILL8
XSTDFILL78_1509 VDD VSS sg13g2_FILL8
XSTDFILL78_1517 VDD VSS sg13g2_FILL8
XSTDFILL78_1525 VDD VSS sg13g2_FILL8
XSTDFILL78_1533 VDD VSS sg13g2_FILL8
XSTDFILL78_1541 VDD VSS sg13g2_FILL8
XSTDFILL78_1549 VDD VSS sg13g2_FILL8
XSTDFILL78_1557 VDD VSS sg13g2_FILL8
XSTDFILL78_1565 VDD VSS sg13g2_FILL8
XSTDFILL78_1573 VDD VSS sg13g2_FILL8
XSTDFILL78_1581 VDD VSS sg13g2_FILL8
XSTDFILL78_1589 VDD VSS sg13g2_FILL8
XSTDFILL78_1597 VDD VSS sg13g2_FILL8
XSTDFILL78_1605 VDD VSS sg13g2_FILL8
XSTDFILL78_1613 VDD VSS sg13g2_FILL8
XSTDFILL78_1621 VDD VSS sg13g2_FILL8
XSTDFILL78_1629 VDD VSS sg13g2_FILL8
XSTDFILL78_1637 VDD VSS sg13g2_FILL8
XSTDFILL78_1645 VDD VSS sg13g2_FILL8
XSTDFILL78_1653 VDD VSS sg13g2_FILL8
XSTDFILL78_1661 VDD VSS sg13g2_FILL8
XSTDFILL78_1669 VDD VSS sg13g2_FILL8
XSTDFILL78_1677 VDD VSS sg13g2_FILL8
XSTDFILL78_1685 VDD VSS sg13g2_FILL8
XSTDFILL78_1693 VDD VSS sg13g2_FILL8
XSTDFILL78_1701 VDD VSS sg13g2_FILL8
XSTDFILL78_1709 VDD VSS sg13g2_FILL8
XSTDFILL78_1717 VDD VSS sg13g2_FILL8
XSTDFILL78_1725 VDD VSS sg13g2_FILL8
XSTDFILL78_1733 VDD VSS sg13g2_FILL8
XSTDFILL78_1741 VDD VSS sg13g2_FILL8
XSTDFILL78_1749 VDD VSS sg13g2_FILL8
XSTDFILL78_1757 VDD VSS sg13g2_FILL8
XSTDFILL78_1765 VDD VSS sg13g2_FILL8
XSTDFILL78_1773 VDD VSS sg13g2_FILL8
XSTDFILL78_1781 VDD VSS sg13g2_FILL8
XSTDFILL78_1789 VDD VSS sg13g2_FILL8
XSTDFILL78_1797 VDD VSS sg13g2_FILL8
XSTDFILL78_1805 VDD VSS sg13g2_FILL8
XSTDFILL78_1813 VDD VSS sg13g2_FILL8
XSTDFILL78_1821 VDD VSS sg13g2_FILL8
XSTDFILL78_1829 VDD VSS sg13g2_FILL8
XSTDFILL78_1837 VDD VSS sg13g2_FILL8
XSTDFILL78_1845 VDD VSS sg13g2_FILL8
XSTDFILL78_1853 VDD VSS sg13g2_FILL8
XSTDFILL78_1861 VDD VSS sg13g2_FILL8
XSTDFILL78_1869 VDD VSS sg13g2_FILL8
XSTDFILL78_1877 VDD VSS sg13g2_FILL8
XSTDFILL78_1885 VDD VSS sg13g2_FILL8
XSTDFILL78_1893 VDD VSS sg13g2_FILL8
XSTDFILL78_1901 VDD VSS sg13g2_FILL8
XSTDFILL78_1909 VDD VSS sg13g2_FILL8
XSTDFILL78_1917 VDD VSS sg13g2_FILL8
XSTDFILL78_1925 VDD VSS sg13g2_FILL8
XSTDFILL78_1933 VDD VSS sg13g2_FILL8
XSTDFILL78_1941 VDD VSS sg13g2_FILL8
XSTDFILL78_1949 VDD VSS sg13g2_FILL8
XSTDFILL78_1957 VDD VSS sg13g2_FILL8
XSTDFILL78_1965 VDD VSS sg13g2_FILL8
XSTDFILL78_1973 VDD VSS sg13g2_FILL8
XSTDFILL78_1981 VDD VSS sg13g2_FILL8
XSTDFILL78_1989 VDD VSS sg13g2_FILL8
XSTDFILL78_1997 VDD VSS sg13g2_FILL8
XSTDFILL78_2005 VDD VSS sg13g2_FILL8
XSTDFILL78_2013 VDD VSS sg13g2_FILL8
XSTDFILL78_2021 VDD VSS sg13g2_FILL8
XSTDFILL78_2029 VDD VSS sg13g2_FILL8
XSTDFILL78_2037 VDD VSS sg13g2_FILL8
XSTDFILL78_2045 VDD VSS sg13g2_FILL8
XSTDFILL78_2053 VDD VSS sg13g2_FILL8
XSTDFILL78_2061 VDD VSS sg13g2_FILL8
XSTDFILL78_2069 VDD VSS sg13g2_FILL8
XSTDFILL78_2077 VDD VSS sg13g2_FILL8
XSTDFILL78_2085 VDD VSS sg13g2_FILL8
XSTDFILL78_2093 VDD VSS sg13g2_FILL8
XSTDFILL78_2101 VDD VSS sg13g2_FILL8
XSTDFILL78_2109 VDD VSS sg13g2_FILL8
XSTDFILL78_2117 VDD VSS sg13g2_FILL8
XSTDFILL78_2125 VDD VSS sg13g2_FILL8
XSTDFILL78_2133 VDD VSS sg13g2_FILL8
XSTDFILL78_2141 VDD VSS sg13g2_FILL8
XSTDFILL78_2149 VDD VSS sg13g2_FILL4
XSTDFILL78_2153 VDD VSS sg13g2_FILL1
XSTDFILL79_0 VDD VSS sg13g2_FILL8
XSTDFILL79_8 VDD VSS sg13g2_FILL8
XSTDFILL79_16 VDD VSS sg13g2_FILL8
XSTDFILL79_24 VDD VSS sg13g2_FILL8
XSTDFILL79_32 VDD VSS sg13g2_FILL8
XSTDFILL79_40 VDD VSS sg13g2_FILL8
XSTDFILL79_48 VDD VSS sg13g2_FILL8
XSTDFILL79_56 VDD VSS sg13g2_FILL8
XSTDFILL79_64 VDD VSS sg13g2_FILL8
XSTDFILL79_72 VDD VSS sg13g2_FILL8
XSTDFILL79_80 VDD VSS sg13g2_FILL8
XSTDFILL79_88 VDD VSS sg13g2_FILL8
XSTDFILL79_96 VDD VSS sg13g2_FILL8
XSTDFILL79_104 VDD VSS sg13g2_FILL8
XSTDFILL79_112 VDD VSS sg13g2_FILL8
XSTDFILL79_120 VDD VSS sg13g2_FILL8
XSTDFILL79_128 VDD VSS sg13g2_FILL4
XSTDFILL79_1085 VDD VSS sg13g2_FILL8
XSTDFILL79_1093 VDD VSS sg13g2_FILL8
XSTDFILL79_1101 VDD VSS sg13g2_FILL8
XSTDFILL79_1109 VDD VSS sg13g2_FILL8
XSTDFILL79_1117 VDD VSS sg13g2_FILL8
XSTDFILL79_1125 VDD VSS sg13g2_FILL8
XSTDFILL79_1133 VDD VSS sg13g2_FILL8
XSTDFILL79_1141 VDD VSS sg13g2_FILL8
XSTDFILL79_1149 VDD VSS sg13g2_FILL8
XSTDFILL79_1157 VDD VSS sg13g2_FILL8
XSTDFILL79_1165 VDD VSS sg13g2_FILL8
XSTDFILL79_1173 VDD VSS sg13g2_FILL8
XSTDFILL79_1181 VDD VSS sg13g2_FILL8
XSTDFILL79_1189 VDD VSS sg13g2_FILL8
XSTDFILL79_1197 VDD VSS sg13g2_FILL8
XSTDFILL79_1205 VDD VSS sg13g2_FILL8
XSTDFILL79_1213 VDD VSS sg13g2_FILL8
XSTDFILL79_1221 VDD VSS sg13g2_FILL8
XSTDFILL79_1229 VDD VSS sg13g2_FILL8
XSTDFILL79_1237 VDD VSS sg13g2_FILL8
XSTDFILL79_1245 VDD VSS sg13g2_FILL8
XSTDFILL79_1253 VDD VSS sg13g2_FILL8
XSTDFILL79_1261 VDD VSS sg13g2_FILL8
XSTDFILL79_1269 VDD VSS sg13g2_FILL8
XSTDFILL79_1277 VDD VSS sg13g2_FILL8
XSTDFILL79_1285 VDD VSS sg13g2_FILL8
XSTDFILL79_1293 VDD VSS sg13g2_FILL8
XSTDFILL79_1301 VDD VSS sg13g2_FILL8
XSTDFILL79_1309 VDD VSS sg13g2_FILL8
XSTDFILL79_1317 VDD VSS sg13g2_FILL8
XSTDFILL79_1325 VDD VSS sg13g2_FILL8
XSTDFILL79_1333 VDD VSS sg13g2_FILL8
XSTDFILL79_1341 VDD VSS sg13g2_FILL8
XSTDFILL79_1349 VDD VSS sg13g2_FILL8
XSTDFILL79_1357 VDD VSS sg13g2_FILL8
XSTDFILL79_1365 VDD VSS sg13g2_FILL8
XSTDFILL79_1373 VDD VSS sg13g2_FILL8
XSTDFILL79_1381 VDD VSS sg13g2_FILL8
XSTDFILL79_1389 VDD VSS sg13g2_FILL8
XSTDFILL79_1397 VDD VSS sg13g2_FILL8
XSTDFILL79_1405 VDD VSS sg13g2_FILL8
XSTDFILL79_1413 VDD VSS sg13g2_FILL8
XSTDFILL79_1421 VDD VSS sg13g2_FILL8
XSTDFILL79_1429 VDD VSS sg13g2_FILL8
XSTDFILL79_1437 VDD VSS sg13g2_FILL8
XSTDFILL79_1445 VDD VSS sg13g2_FILL8
XSTDFILL79_1453 VDD VSS sg13g2_FILL8
XSTDFILL79_1461 VDD VSS sg13g2_FILL8
XSTDFILL79_1469 VDD VSS sg13g2_FILL8
XSTDFILL79_1477 VDD VSS sg13g2_FILL8
XSTDFILL79_1485 VDD VSS sg13g2_FILL8
XSTDFILL79_1493 VDD VSS sg13g2_FILL8
XSTDFILL79_1501 VDD VSS sg13g2_FILL8
XSTDFILL79_1509 VDD VSS sg13g2_FILL8
XSTDFILL79_1517 VDD VSS sg13g2_FILL8
XSTDFILL79_1525 VDD VSS sg13g2_FILL8
XSTDFILL79_1533 VDD VSS sg13g2_FILL8
XSTDFILL79_1541 VDD VSS sg13g2_FILL8
XSTDFILL79_1549 VDD VSS sg13g2_FILL8
XSTDFILL79_1557 VDD VSS sg13g2_FILL8
XSTDFILL79_1565 VDD VSS sg13g2_FILL8
XSTDFILL79_1573 VDD VSS sg13g2_FILL8
XSTDFILL79_1581 VDD VSS sg13g2_FILL8
XSTDFILL79_1589 VDD VSS sg13g2_FILL8
XSTDFILL79_1597 VDD VSS sg13g2_FILL8
XSTDFILL79_1605 VDD VSS sg13g2_FILL8
XSTDFILL79_1613 VDD VSS sg13g2_FILL8
XSTDFILL79_1621 VDD VSS sg13g2_FILL8
XSTDFILL79_1629 VDD VSS sg13g2_FILL8
XSTDFILL79_1637 VDD VSS sg13g2_FILL8
XSTDFILL79_1645 VDD VSS sg13g2_FILL8
XSTDFILL79_1653 VDD VSS sg13g2_FILL8
XSTDFILL79_1661 VDD VSS sg13g2_FILL8
XSTDFILL79_1669 VDD VSS sg13g2_FILL8
XSTDFILL79_1677 VDD VSS sg13g2_FILL8
XSTDFILL79_1685 VDD VSS sg13g2_FILL8
XSTDFILL79_1693 VDD VSS sg13g2_FILL8
XSTDFILL79_1701 VDD VSS sg13g2_FILL8
XSTDFILL79_1709 VDD VSS sg13g2_FILL8
XSTDFILL79_1717 VDD VSS sg13g2_FILL8
XSTDFILL79_1725 VDD VSS sg13g2_FILL8
XSTDFILL79_1733 VDD VSS sg13g2_FILL8
XSTDFILL79_1741 VDD VSS sg13g2_FILL8
XSTDFILL79_1749 VDD VSS sg13g2_FILL8
XSTDFILL79_1757 VDD VSS sg13g2_FILL8
XSTDFILL79_1765 VDD VSS sg13g2_FILL8
XSTDFILL79_1773 VDD VSS sg13g2_FILL8
XSTDFILL79_1781 VDD VSS sg13g2_FILL8
XSTDFILL79_1789 VDD VSS sg13g2_FILL8
XSTDFILL79_1797 VDD VSS sg13g2_FILL8
XSTDFILL79_1805 VDD VSS sg13g2_FILL8
XSTDFILL79_1813 VDD VSS sg13g2_FILL8
XSTDFILL79_1821 VDD VSS sg13g2_FILL8
XSTDFILL79_1829 VDD VSS sg13g2_FILL8
XSTDFILL79_1837 VDD VSS sg13g2_FILL8
XSTDFILL79_1845 VDD VSS sg13g2_FILL8
XSTDFILL79_1853 VDD VSS sg13g2_FILL8
XSTDFILL79_1861 VDD VSS sg13g2_FILL8
XSTDFILL79_1869 VDD VSS sg13g2_FILL8
XSTDFILL79_1877 VDD VSS sg13g2_FILL8
XSTDFILL79_1885 VDD VSS sg13g2_FILL8
XSTDFILL79_1893 VDD VSS sg13g2_FILL8
XSTDFILL79_1901 VDD VSS sg13g2_FILL8
XSTDFILL79_1909 VDD VSS sg13g2_FILL8
XSTDFILL79_1917 VDD VSS sg13g2_FILL8
XSTDFILL79_1925 VDD VSS sg13g2_FILL8
XSTDFILL79_1933 VDD VSS sg13g2_FILL8
XSTDFILL79_1941 VDD VSS sg13g2_FILL8
XSTDFILL79_1949 VDD VSS sg13g2_FILL8
XSTDFILL79_1957 VDD VSS sg13g2_FILL8
XSTDFILL79_1965 VDD VSS sg13g2_FILL8
XSTDFILL79_1973 VDD VSS sg13g2_FILL8
XSTDFILL79_1981 VDD VSS sg13g2_FILL8
XSTDFILL79_1989 VDD VSS sg13g2_FILL8
XSTDFILL79_1997 VDD VSS sg13g2_FILL8
XSTDFILL79_2005 VDD VSS sg13g2_FILL8
XSTDFILL79_2013 VDD VSS sg13g2_FILL8
XSTDFILL79_2021 VDD VSS sg13g2_FILL8
XSTDFILL79_2029 VDD VSS sg13g2_FILL8
XSTDFILL79_2037 VDD VSS sg13g2_FILL8
XSTDFILL79_2045 VDD VSS sg13g2_FILL8
XSTDFILL79_2053 VDD VSS sg13g2_FILL8
XSTDFILL79_2061 VDD VSS sg13g2_FILL8
XSTDFILL79_2069 VDD VSS sg13g2_FILL8
XSTDFILL79_2077 VDD VSS sg13g2_FILL8
XSTDFILL79_2085 VDD VSS sg13g2_FILL8
XSTDFILL79_2093 VDD VSS sg13g2_FILL8
XSTDFILL79_2101 VDD VSS sg13g2_FILL8
XSTDFILL79_2109 VDD VSS sg13g2_FILL8
XSTDFILL79_2117 VDD VSS sg13g2_FILL8
XSTDFILL79_2125 VDD VSS sg13g2_FILL8
XSTDFILL79_2133 VDD VSS sg13g2_FILL8
XSTDFILL79_2141 VDD VSS sg13g2_FILL8
XSTDFILL79_2149 VDD VSS sg13g2_FILL4
XSTDFILL79_2153 VDD VSS sg13g2_FILL1
XSTDFILL80_0 VDD VSS sg13g2_FILL8
XSTDFILL80_8 VDD VSS sg13g2_FILL8
XSTDFILL80_16 VDD VSS sg13g2_FILL8
XSTDFILL80_24 VDD VSS sg13g2_FILL8
XSTDFILL80_32 VDD VSS sg13g2_FILL8
XSTDFILL80_40 VDD VSS sg13g2_FILL8
XSTDFILL80_48 VDD VSS sg13g2_FILL8
XSTDFILL80_56 VDD VSS sg13g2_FILL8
XSTDFILL80_64 VDD VSS sg13g2_FILL8
XSTDFILL80_72 VDD VSS sg13g2_FILL8
XSTDFILL80_80 VDD VSS sg13g2_FILL8
XSTDFILL80_88 VDD VSS sg13g2_FILL8
XSTDFILL80_96 VDD VSS sg13g2_FILL8
XSTDFILL80_104 VDD VSS sg13g2_FILL8
XSTDFILL80_112 VDD VSS sg13g2_FILL8
XSTDFILL80_120 VDD VSS sg13g2_FILL8
XSTDFILL80_128 VDD VSS sg13g2_FILL4
XSTDFILL80_1085 VDD VSS sg13g2_FILL8
XSTDFILL80_1093 VDD VSS sg13g2_FILL8
XSTDFILL80_1101 VDD VSS sg13g2_FILL8
XSTDFILL80_1109 VDD VSS sg13g2_FILL8
XSTDFILL80_1117 VDD VSS sg13g2_FILL8
XSTDFILL80_1125 VDD VSS sg13g2_FILL8
XSTDFILL80_1133 VDD VSS sg13g2_FILL8
XSTDFILL80_1141 VDD VSS sg13g2_FILL8
XSTDFILL80_1149 VDD VSS sg13g2_FILL8
XSTDFILL80_1157 VDD VSS sg13g2_FILL8
XSTDFILL80_1165 VDD VSS sg13g2_FILL8
XSTDFILL80_1173 VDD VSS sg13g2_FILL8
XSTDFILL80_1181 VDD VSS sg13g2_FILL8
XSTDFILL80_1189 VDD VSS sg13g2_FILL8
XSTDFILL80_1197 VDD VSS sg13g2_FILL8
XSTDFILL80_1205 VDD VSS sg13g2_FILL8
XSTDFILL80_1213 VDD VSS sg13g2_FILL8
XSTDFILL80_1221 VDD VSS sg13g2_FILL8
XSTDFILL80_1229 VDD VSS sg13g2_FILL8
XSTDFILL80_1237 VDD VSS sg13g2_FILL8
XSTDFILL80_1245 VDD VSS sg13g2_FILL8
XSTDFILL80_1253 VDD VSS sg13g2_FILL8
XSTDFILL80_1261 VDD VSS sg13g2_FILL8
XSTDFILL80_1269 VDD VSS sg13g2_FILL8
XSTDFILL80_1277 VDD VSS sg13g2_FILL8
XSTDFILL80_1285 VDD VSS sg13g2_FILL8
XSTDFILL80_1293 VDD VSS sg13g2_FILL8
XSTDFILL80_1301 VDD VSS sg13g2_FILL8
XSTDFILL80_1309 VDD VSS sg13g2_FILL8
XSTDFILL80_1317 VDD VSS sg13g2_FILL8
XSTDFILL80_1325 VDD VSS sg13g2_FILL8
XSTDFILL80_1333 VDD VSS sg13g2_FILL8
XSTDFILL80_1341 VDD VSS sg13g2_FILL8
XSTDFILL80_1349 VDD VSS sg13g2_FILL8
XSTDFILL80_1357 VDD VSS sg13g2_FILL8
XSTDFILL80_1365 VDD VSS sg13g2_FILL8
XSTDFILL80_1373 VDD VSS sg13g2_FILL8
XSTDFILL80_1381 VDD VSS sg13g2_FILL8
XSTDFILL80_1389 VDD VSS sg13g2_FILL8
XSTDFILL80_1397 VDD VSS sg13g2_FILL8
XSTDFILL80_1405 VDD VSS sg13g2_FILL8
XSTDFILL80_1413 VDD VSS sg13g2_FILL8
XSTDFILL80_1421 VDD VSS sg13g2_FILL8
XSTDFILL80_1429 VDD VSS sg13g2_FILL8
XSTDFILL80_1437 VDD VSS sg13g2_FILL8
XSTDFILL80_1445 VDD VSS sg13g2_FILL8
XSTDFILL80_1453 VDD VSS sg13g2_FILL8
XSTDFILL80_1461 VDD VSS sg13g2_FILL8
XSTDFILL80_1469 VDD VSS sg13g2_FILL8
XSTDFILL80_1477 VDD VSS sg13g2_FILL8
XSTDFILL80_1485 VDD VSS sg13g2_FILL8
XSTDFILL80_1493 VDD VSS sg13g2_FILL8
XSTDFILL80_1501 VDD VSS sg13g2_FILL8
XSTDFILL80_1509 VDD VSS sg13g2_FILL8
XSTDFILL80_1517 VDD VSS sg13g2_FILL8
XSTDFILL80_1525 VDD VSS sg13g2_FILL8
XSTDFILL80_1533 VDD VSS sg13g2_FILL8
XSTDFILL80_1541 VDD VSS sg13g2_FILL8
XSTDFILL80_1549 VDD VSS sg13g2_FILL8
XSTDFILL80_1557 VDD VSS sg13g2_FILL8
XSTDFILL80_1565 VDD VSS sg13g2_FILL8
XSTDFILL80_1573 VDD VSS sg13g2_FILL8
XSTDFILL80_1581 VDD VSS sg13g2_FILL8
XSTDFILL80_1589 VDD VSS sg13g2_FILL8
XSTDFILL80_1597 VDD VSS sg13g2_FILL8
XSTDFILL80_1605 VDD VSS sg13g2_FILL8
XSTDFILL80_1613 VDD VSS sg13g2_FILL8
XSTDFILL80_1621 VDD VSS sg13g2_FILL8
XSTDFILL80_1629 VDD VSS sg13g2_FILL8
XSTDFILL80_1637 VDD VSS sg13g2_FILL8
XSTDFILL80_1645 VDD VSS sg13g2_FILL8
XSTDFILL80_1653 VDD VSS sg13g2_FILL8
XSTDFILL80_1661 VDD VSS sg13g2_FILL8
XSTDFILL80_1669 VDD VSS sg13g2_FILL8
XSTDFILL80_1677 VDD VSS sg13g2_FILL8
XSTDFILL80_1685 VDD VSS sg13g2_FILL8
XSTDFILL80_1693 VDD VSS sg13g2_FILL8
XSTDFILL80_1701 VDD VSS sg13g2_FILL8
XSTDFILL80_1709 VDD VSS sg13g2_FILL8
XSTDFILL80_1717 VDD VSS sg13g2_FILL8
XSTDFILL80_1725 VDD VSS sg13g2_FILL8
XSTDFILL80_1733 VDD VSS sg13g2_FILL8
XSTDFILL80_1741 VDD VSS sg13g2_FILL8
XSTDFILL80_1749 VDD VSS sg13g2_FILL8
XSTDFILL80_1757 VDD VSS sg13g2_FILL8
XSTDFILL80_1765 VDD VSS sg13g2_FILL8
XSTDFILL80_1773 VDD VSS sg13g2_FILL8
XSTDFILL80_1781 VDD VSS sg13g2_FILL8
XSTDFILL80_1789 VDD VSS sg13g2_FILL8
XSTDFILL80_1797 VDD VSS sg13g2_FILL8
XSTDFILL80_1805 VDD VSS sg13g2_FILL8
XSTDFILL80_1813 VDD VSS sg13g2_FILL8
XSTDFILL80_1821 VDD VSS sg13g2_FILL8
XSTDFILL80_1829 VDD VSS sg13g2_FILL8
XSTDFILL80_1837 VDD VSS sg13g2_FILL8
XSTDFILL80_1845 VDD VSS sg13g2_FILL8
XSTDFILL80_1853 VDD VSS sg13g2_FILL8
XSTDFILL80_1861 VDD VSS sg13g2_FILL8
XSTDFILL80_1869 VDD VSS sg13g2_FILL8
XSTDFILL80_1877 VDD VSS sg13g2_FILL8
XSTDFILL80_1885 VDD VSS sg13g2_FILL8
XSTDFILL80_1893 VDD VSS sg13g2_FILL8
XSTDFILL80_1901 VDD VSS sg13g2_FILL8
XSTDFILL80_1909 VDD VSS sg13g2_FILL8
XSTDFILL80_1917 VDD VSS sg13g2_FILL8
XSTDFILL80_1925 VDD VSS sg13g2_FILL8
XSTDFILL80_1933 VDD VSS sg13g2_FILL8
XSTDFILL80_1941 VDD VSS sg13g2_FILL8
XSTDFILL80_1949 VDD VSS sg13g2_FILL8
XSTDFILL80_1957 VDD VSS sg13g2_FILL8
XSTDFILL80_1965 VDD VSS sg13g2_FILL8
XSTDFILL80_1973 VDD VSS sg13g2_FILL8
XSTDFILL80_1981 VDD VSS sg13g2_FILL8
XSTDFILL80_1989 VDD VSS sg13g2_FILL8
XSTDFILL80_1997 VDD VSS sg13g2_FILL8
XSTDFILL80_2005 VDD VSS sg13g2_FILL8
XSTDFILL80_2013 VDD VSS sg13g2_FILL8
XSTDFILL80_2021 VDD VSS sg13g2_FILL8
XSTDFILL80_2029 VDD VSS sg13g2_FILL8
XSTDFILL80_2037 VDD VSS sg13g2_FILL8
XSTDFILL80_2045 VDD VSS sg13g2_FILL8
XSTDFILL80_2053 VDD VSS sg13g2_FILL8
XSTDFILL80_2061 VDD VSS sg13g2_FILL8
XSTDFILL80_2069 VDD VSS sg13g2_FILL8
XSTDFILL80_2077 VDD VSS sg13g2_FILL8
XSTDFILL80_2085 VDD VSS sg13g2_FILL8
XSTDFILL80_2093 VDD VSS sg13g2_FILL8
XSTDFILL80_2101 VDD VSS sg13g2_FILL8
XSTDFILL80_2109 VDD VSS sg13g2_FILL8
XSTDFILL80_2117 VDD VSS sg13g2_FILL8
XSTDFILL80_2125 VDD VSS sg13g2_FILL8
XSTDFILL80_2133 VDD VSS sg13g2_FILL8
XSTDFILL80_2141 VDD VSS sg13g2_FILL8
XSTDFILL80_2149 VDD VSS sg13g2_FILL4
XSTDFILL80_2153 VDD VSS sg13g2_FILL1
XSTDFILL81_0 VDD VSS sg13g2_FILL8
XSTDFILL81_8 VDD VSS sg13g2_FILL8
XSTDFILL81_16 VDD VSS sg13g2_FILL8
XSTDFILL81_24 VDD VSS sg13g2_FILL8
XSTDFILL81_32 VDD VSS sg13g2_FILL8
XSTDFILL81_40 VDD VSS sg13g2_FILL8
XSTDFILL81_48 VDD VSS sg13g2_FILL8
XSTDFILL81_56 VDD VSS sg13g2_FILL8
XSTDFILL81_64 VDD VSS sg13g2_FILL8
XSTDFILL81_72 VDD VSS sg13g2_FILL8
XSTDFILL81_80 VDD VSS sg13g2_FILL8
XSTDFILL81_88 VDD VSS sg13g2_FILL8
XSTDFILL81_96 VDD VSS sg13g2_FILL8
XSTDFILL81_104 VDD VSS sg13g2_FILL8
XSTDFILL81_112 VDD VSS sg13g2_FILL8
XSTDFILL81_120 VDD VSS sg13g2_FILL8
XSTDFILL81_128 VDD VSS sg13g2_FILL4
XSTDFILL81_1085 VDD VSS sg13g2_FILL8
XSTDFILL81_1093 VDD VSS sg13g2_FILL8
XSTDFILL81_1101 VDD VSS sg13g2_FILL8
XSTDFILL81_1109 VDD VSS sg13g2_FILL8
XSTDFILL81_1117 VDD VSS sg13g2_FILL8
XSTDFILL81_1125 VDD VSS sg13g2_FILL8
XSTDFILL81_1133 VDD VSS sg13g2_FILL8
XSTDFILL81_1141 VDD VSS sg13g2_FILL8
XSTDFILL81_1149 VDD VSS sg13g2_FILL8
XSTDFILL81_1157 VDD VSS sg13g2_FILL8
XSTDFILL81_1165 VDD VSS sg13g2_FILL8
XSTDFILL81_1173 VDD VSS sg13g2_FILL8
XSTDFILL81_1181 VDD VSS sg13g2_FILL8
XSTDFILL81_1189 VDD VSS sg13g2_FILL8
XSTDFILL81_1197 VDD VSS sg13g2_FILL8
XSTDFILL81_1205 VDD VSS sg13g2_FILL8
XSTDFILL81_1213 VDD VSS sg13g2_FILL8
XSTDFILL81_1221 VDD VSS sg13g2_FILL8
XSTDFILL81_1229 VDD VSS sg13g2_FILL8
XSTDFILL81_1237 VDD VSS sg13g2_FILL8
XSTDFILL81_1245 VDD VSS sg13g2_FILL8
XSTDFILL81_1253 VDD VSS sg13g2_FILL8
XSTDFILL81_1261 VDD VSS sg13g2_FILL8
XSTDFILL81_1269 VDD VSS sg13g2_FILL8
XSTDFILL81_1277 VDD VSS sg13g2_FILL8
XSTDFILL81_1285 VDD VSS sg13g2_FILL8
XSTDFILL81_1293 VDD VSS sg13g2_FILL8
XSTDFILL81_1301 VDD VSS sg13g2_FILL8
XSTDFILL81_1309 VDD VSS sg13g2_FILL8
XSTDFILL81_1317 VDD VSS sg13g2_FILL8
XSTDFILL81_1325 VDD VSS sg13g2_FILL8
XSTDFILL81_1333 VDD VSS sg13g2_FILL8
XSTDFILL81_1341 VDD VSS sg13g2_FILL8
XSTDFILL81_1349 VDD VSS sg13g2_FILL8
XSTDFILL81_1357 VDD VSS sg13g2_FILL8
XSTDFILL81_1365 VDD VSS sg13g2_FILL8
XSTDFILL81_1373 VDD VSS sg13g2_FILL8
XSTDFILL81_1381 VDD VSS sg13g2_FILL8
XSTDFILL81_1389 VDD VSS sg13g2_FILL8
XSTDFILL81_1397 VDD VSS sg13g2_FILL8
XSTDFILL81_1405 VDD VSS sg13g2_FILL8
XSTDFILL81_1413 VDD VSS sg13g2_FILL8
XSTDFILL81_1421 VDD VSS sg13g2_FILL8
XSTDFILL81_1429 VDD VSS sg13g2_FILL8
XSTDFILL81_1437 VDD VSS sg13g2_FILL8
XSTDFILL81_1445 VDD VSS sg13g2_FILL8
XSTDFILL81_1453 VDD VSS sg13g2_FILL8
XSTDFILL81_1461 VDD VSS sg13g2_FILL8
XSTDFILL81_1469 VDD VSS sg13g2_FILL8
XSTDFILL81_1477 VDD VSS sg13g2_FILL8
XSTDFILL81_1485 VDD VSS sg13g2_FILL8
XSTDFILL81_1493 VDD VSS sg13g2_FILL8
XSTDFILL81_1501 VDD VSS sg13g2_FILL8
XSTDFILL81_1509 VDD VSS sg13g2_FILL8
XSTDFILL81_1517 VDD VSS sg13g2_FILL8
XSTDFILL81_1525 VDD VSS sg13g2_FILL8
XSTDFILL81_1533 VDD VSS sg13g2_FILL8
XSTDFILL81_1541 VDD VSS sg13g2_FILL8
XSTDFILL81_1549 VDD VSS sg13g2_FILL8
XSTDFILL81_1557 VDD VSS sg13g2_FILL8
XSTDFILL81_1565 VDD VSS sg13g2_FILL8
XSTDFILL81_1573 VDD VSS sg13g2_FILL8
XSTDFILL81_1581 VDD VSS sg13g2_FILL8
XSTDFILL81_1589 VDD VSS sg13g2_FILL8
XSTDFILL81_1597 VDD VSS sg13g2_FILL8
XSTDFILL81_1605 VDD VSS sg13g2_FILL8
XSTDFILL81_1613 VDD VSS sg13g2_FILL8
XSTDFILL81_1621 VDD VSS sg13g2_FILL8
XSTDFILL81_1629 VDD VSS sg13g2_FILL8
XSTDFILL81_1637 VDD VSS sg13g2_FILL8
XSTDFILL81_1645 VDD VSS sg13g2_FILL8
XSTDFILL81_1653 VDD VSS sg13g2_FILL8
XSTDFILL81_1661 VDD VSS sg13g2_FILL8
XSTDFILL81_1669 VDD VSS sg13g2_FILL8
XSTDFILL81_1677 VDD VSS sg13g2_FILL8
XSTDFILL81_1685 VDD VSS sg13g2_FILL8
XSTDFILL81_1693 VDD VSS sg13g2_FILL8
XSTDFILL81_1701 VDD VSS sg13g2_FILL8
XSTDFILL81_1709 VDD VSS sg13g2_FILL8
XSTDFILL81_1717 VDD VSS sg13g2_FILL8
XSTDFILL81_1725 VDD VSS sg13g2_FILL8
XSTDFILL81_1733 VDD VSS sg13g2_FILL8
XSTDFILL81_1741 VDD VSS sg13g2_FILL8
XSTDFILL81_1749 VDD VSS sg13g2_FILL8
XSTDFILL81_1757 VDD VSS sg13g2_FILL8
XSTDFILL81_1765 VDD VSS sg13g2_FILL8
XSTDFILL81_1773 VDD VSS sg13g2_FILL8
XSTDFILL81_1781 VDD VSS sg13g2_FILL8
XSTDFILL81_1789 VDD VSS sg13g2_FILL8
XSTDFILL81_1797 VDD VSS sg13g2_FILL8
XSTDFILL81_1805 VDD VSS sg13g2_FILL8
XSTDFILL81_1813 VDD VSS sg13g2_FILL8
XSTDFILL81_1821 VDD VSS sg13g2_FILL8
XSTDFILL81_1829 VDD VSS sg13g2_FILL8
XSTDFILL81_1837 VDD VSS sg13g2_FILL8
XSTDFILL81_1845 VDD VSS sg13g2_FILL8
XSTDFILL81_1853 VDD VSS sg13g2_FILL8
XSTDFILL81_1861 VDD VSS sg13g2_FILL8
XSTDFILL81_1869 VDD VSS sg13g2_FILL8
XSTDFILL81_1877 VDD VSS sg13g2_FILL8
XSTDFILL81_1885 VDD VSS sg13g2_FILL8
XSTDFILL81_1893 VDD VSS sg13g2_FILL8
XSTDFILL81_1901 VDD VSS sg13g2_FILL8
XSTDFILL81_1909 VDD VSS sg13g2_FILL8
XSTDFILL81_1917 VDD VSS sg13g2_FILL8
XSTDFILL81_1925 VDD VSS sg13g2_FILL8
XSTDFILL81_1933 VDD VSS sg13g2_FILL8
XSTDFILL81_1941 VDD VSS sg13g2_FILL8
XSTDFILL81_1949 VDD VSS sg13g2_FILL8
XSTDFILL81_1957 VDD VSS sg13g2_FILL8
XSTDFILL81_1965 VDD VSS sg13g2_FILL8
XSTDFILL81_1973 VDD VSS sg13g2_FILL8
XSTDFILL81_1981 VDD VSS sg13g2_FILL8
XSTDFILL81_1989 VDD VSS sg13g2_FILL8
XSTDFILL81_1997 VDD VSS sg13g2_FILL8
XSTDFILL81_2005 VDD VSS sg13g2_FILL8
XSTDFILL81_2013 VDD VSS sg13g2_FILL8
XSTDFILL81_2021 VDD VSS sg13g2_FILL8
XSTDFILL81_2029 VDD VSS sg13g2_FILL8
XSTDFILL81_2037 VDD VSS sg13g2_FILL8
XSTDFILL81_2045 VDD VSS sg13g2_FILL8
XSTDFILL81_2053 VDD VSS sg13g2_FILL8
XSTDFILL81_2061 VDD VSS sg13g2_FILL8
XSTDFILL81_2069 VDD VSS sg13g2_FILL8
XSTDFILL81_2077 VDD VSS sg13g2_FILL8
XSTDFILL81_2085 VDD VSS sg13g2_FILL8
XSTDFILL81_2093 VDD VSS sg13g2_FILL8
XSTDFILL81_2101 VDD VSS sg13g2_FILL8
XSTDFILL81_2109 VDD VSS sg13g2_FILL8
XSTDFILL81_2117 VDD VSS sg13g2_FILL8
XSTDFILL81_2125 VDD VSS sg13g2_FILL8
XSTDFILL81_2133 VDD VSS sg13g2_FILL8
XSTDFILL81_2141 VDD VSS sg13g2_FILL8
XSTDFILL81_2149 VDD VSS sg13g2_FILL4
XSTDFILL81_2153 VDD VSS sg13g2_FILL1
XSTDFILL82_0 VDD VSS sg13g2_FILL8
XSTDFILL82_8 VDD VSS sg13g2_FILL8
XSTDFILL82_16 VDD VSS sg13g2_FILL8
XSTDFILL82_24 VDD VSS sg13g2_FILL8
XSTDFILL82_32 VDD VSS sg13g2_FILL8
XSTDFILL82_40 VDD VSS sg13g2_FILL8
XSTDFILL82_48 VDD VSS sg13g2_FILL8
XSTDFILL82_56 VDD VSS sg13g2_FILL8
XSTDFILL82_64 VDD VSS sg13g2_FILL8
XSTDFILL82_72 VDD VSS sg13g2_FILL8
XSTDFILL82_80 VDD VSS sg13g2_FILL8
XSTDFILL82_88 VDD VSS sg13g2_FILL8
XSTDFILL82_96 VDD VSS sg13g2_FILL8
XSTDFILL82_104 VDD VSS sg13g2_FILL8
XSTDFILL82_112 VDD VSS sg13g2_FILL8
XSTDFILL82_120 VDD VSS sg13g2_FILL8
XSTDFILL82_128 VDD VSS sg13g2_FILL4
XSTDFILL82_1085 VDD VSS sg13g2_FILL8
XSTDFILL82_1093 VDD VSS sg13g2_FILL8
XSTDFILL82_1101 VDD VSS sg13g2_FILL8
XSTDFILL82_1109 VDD VSS sg13g2_FILL8
XSTDFILL82_1117 VDD VSS sg13g2_FILL8
XSTDFILL82_1125 VDD VSS sg13g2_FILL8
XSTDFILL82_1133 VDD VSS sg13g2_FILL8
XSTDFILL82_1141 VDD VSS sg13g2_FILL8
XSTDFILL82_1149 VDD VSS sg13g2_FILL8
XSTDFILL82_1157 VDD VSS sg13g2_FILL8
XSTDFILL82_1165 VDD VSS sg13g2_FILL8
XSTDFILL82_1173 VDD VSS sg13g2_FILL8
XSTDFILL82_1181 VDD VSS sg13g2_FILL8
XSTDFILL82_1189 VDD VSS sg13g2_FILL8
XSTDFILL82_1197 VDD VSS sg13g2_FILL8
XSTDFILL82_1205 VDD VSS sg13g2_FILL8
XSTDFILL82_1213 VDD VSS sg13g2_FILL8
XSTDFILL82_1221 VDD VSS sg13g2_FILL8
XSTDFILL82_1229 VDD VSS sg13g2_FILL8
XSTDFILL82_1237 VDD VSS sg13g2_FILL8
XSTDFILL82_1245 VDD VSS sg13g2_FILL8
XSTDFILL82_1253 VDD VSS sg13g2_FILL8
XSTDFILL82_1261 VDD VSS sg13g2_FILL8
XSTDFILL82_1269 VDD VSS sg13g2_FILL8
XSTDFILL82_1277 VDD VSS sg13g2_FILL8
XSTDFILL82_1285 VDD VSS sg13g2_FILL8
XSTDFILL82_1293 VDD VSS sg13g2_FILL8
XSTDFILL82_1301 VDD VSS sg13g2_FILL8
XSTDFILL82_1309 VDD VSS sg13g2_FILL8
XSTDFILL82_1317 VDD VSS sg13g2_FILL8
XSTDFILL82_1325 VDD VSS sg13g2_FILL8
XSTDFILL82_1333 VDD VSS sg13g2_FILL8
XSTDFILL82_1341 VDD VSS sg13g2_FILL8
XSTDFILL82_1349 VDD VSS sg13g2_FILL8
XSTDFILL82_1357 VDD VSS sg13g2_FILL8
XSTDFILL82_1365 VDD VSS sg13g2_FILL8
XSTDFILL82_1373 VDD VSS sg13g2_FILL8
XSTDFILL82_1381 VDD VSS sg13g2_FILL8
XSTDFILL82_1389 VDD VSS sg13g2_FILL8
XSTDFILL82_1397 VDD VSS sg13g2_FILL8
XSTDFILL82_1405 VDD VSS sg13g2_FILL8
XSTDFILL82_1413 VDD VSS sg13g2_FILL8
XSTDFILL82_1421 VDD VSS sg13g2_FILL8
XSTDFILL82_1429 VDD VSS sg13g2_FILL8
XSTDFILL82_1437 VDD VSS sg13g2_FILL8
XSTDFILL82_1445 VDD VSS sg13g2_FILL8
XSTDFILL82_1453 VDD VSS sg13g2_FILL8
XSTDFILL82_1461 VDD VSS sg13g2_FILL8
XSTDFILL82_1469 VDD VSS sg13g2_FILL8
XSTDFILL82_1477 VDD VSS sg13g2_FILL8
XSTDFILL82_1485 VDD VSS sg13g2_FILL8
XSTDFILL82_1493 VDD VSS sg13g2_FILL8
XSTDFILL82_1501 VDD VSS sg13g2_FILL8
XSTDFILL82_1509 VDD VSS sg13g2_FILL8
XSTDFILL82_1517 VDD VSS sg13g2_FILL8
XSTDFILL82_1525 VDD VSS sg13g2_FILL8
XSTDFILL82_1533 VDD VSS sg13g2_FILL8
XSTDFILL82_1541 VDD VSS sg13g2_FILL8
XSTDFILL82_1549 VDD VSS sg13g2_FILL8
XSTDFILL82_1557 VDD VSS sg13g2_FILL8
XSTDFILL82_1565 VDD VSS sg13g2_FILL8
XSTDFILL82_1573 VDD VSS sg13g2_FILL8
XSTDFILL82_1581 VDD VSS sg13g2_FILL8
XSTDFILL82_1589 VDD VSS sg13g2_FILL8
XSTDFILL82_1597 VDD VSS sg13g2_FILL8
XSTDFILL82_1605 VDD VSS sg13g2_FILL8
XSTDFILL82_1613 VDD VSS sg13g2_FILL8
XSTDFILL82_1621 VDD VSS sg13g2_FILL8
XSTDFILL82_1629 VDD VSS sg13g2_FILL8
XSTDFILL82_1637 VDD VSS sg13g2_FILL8
XSTDFILL82_1645 VDD VSS sg13g2_FILL8
XSTDFILL82_1653 VDD VSS sg13g2_FILL8
XSTDFILL82_1661 VDD VSS sg13g2_FILL8
XSTDFILL82_1669 VDD VSS sg13g2_FILL8
XSTDFILL82_1677 VDD VSS sg13g2_FILL8
XSTDFILL82_1685 VDD VSS sg13g2_FILL8
XSTDFILL82_1693 VDD VSS sg13g2_FILL8
XSTDFILL82_1701 VDD VSS sg13g2_FILL8
XSTDFILL82_1709 VDD VSS sg13g2_FILL8
XSTDFILL82_1717 VDD VSS sg13g2_FILL8
XSTDFILL82_1725 VDD VSS sg13g2_FILL8
XSTDFILL82_1733 VDD VSS sg13g2_FILL8
XSTDFILL82_1741 VDD VSS sg13g2_FILL8
XSTDFILL82_1749 VDD VSS sg13g2_FILL8
XSTDFILL82_1757 VDD VSS sg13g2_FILL8
XSTDFILL82_1765 VDD VSS sg13g2_FILL8
XSTDFILL82_1773 VDD VSS sg13g2_FILL8
XSTDFILL82_1781 VDD VSS sg13g2_FILL8
XSTDFILL82_1789 VDD VSS sg13g2_FILL8
XSTDFILL82_1797 VDD VSS sg13g2_FILL8
XSTDFILL82_1805 VDD VSS sg13g2_FILL8
XSTDFILL82_1813 VDD VSS sg13g2_FILL8
XSTDFILL82_1821 VDD VSS sg13g2_FILL8
XSTDFILL82_1829 VDD VSS sg13g2_FILL8
XSTDFILL82_1837 VDD VSS sg13g2_FILL8
XSTDFILL82_1845 VDD VSS sg13g2_FILL8
XSTDFILL82_1853 VDD VSS sg13g2_FILL8
XSTDFILL82_1861 VDD VSS sg13g2_FILL8
XSTDFILL82_1869 VDD VSS sg13g2_FILL8
XSTDFILL82_1877 VDD VSS sg13g2_FILL8
XSTDFILL82_1885 VDD VSS sg13g2_FILL8
XSTDFILL82_1893 VDD VSS sg13g2_FILL8
XSTDFILL82_1901 VDD VSS sg13g2_FILL8
XSTDFILL82_1909 VDD VSS sg13g2_FILL8
XSTDFILL82_1917 VDD VSS sg13g2_FILL8
XSTDFILL82_1925 VDD VSS sg13g2_FILL8
XSTDFILL82_1933 VDD VSS sg13g2_FILL8
XSTDFILL82_1941 VDD VSS sg13g2_FILL8
XSTDFILL82_1949 VDD VSS sg13g2_FILL8
XSTDFILL82_1957 VDD VSS sg13g2_FILL8
XSTDFILL82_1965 VDD VSS sg13g2_FILL8
XSTDFILL82_1973 VDD VSS sg13g2_FILL8
XSTDFILL82_1981 VDD VSS sg13g2_FILL8
XSTDFILL82_1989 VDD VSS sg13g2_FILL8
XSTDFILL82_1997 VDD VSS sg13g2_FILL8
XSTDFILL82_2005 VDD VSS sg13g2_FILL8
XSTDFILL82_2013 VDD VSS sg13g2_FILL8
XSTDFILL82_2021 VDD VSS sg13g2_FILL8
XSTDFILL82_2029 VDD VSS sg13g2_FILL8
XSTDFILL82_2037 VDD VSS sg13g2_FILL8
XSTDFILL82_2045 VDD VSS sg13g2_FILL8
XSTDFILL82_2053 VDD VSS sg13g2_FILL8
XSTDFILL82_2061 VDD VSS sg13g2_FILL8
XSTDFILL82_2069 VDD VSS sg13g2_FILL8
XSTDFILL82_2077 VDD VSS sg13g2_FILL8
XSTDFILL82_2085 VDD VSS sg13g2_FILL8
XSTDFILL82_2093 VDD VSS sg13g2_FILL8
XSTDFILL82_2101 VDD VSS sg13g2_FILL8
XSTDFILL82_2109 VDD VSS sg13g2_FILL8
XSTDFILL82_2117 VDD VSS sg13g2_FILL8
XSTDFILL82_2125 VDD VSS sg13g2_FILL8
XSTDFILL82_2133 VDD VSS sg13g2_FILL8
XSTDFILL82_2141 VDD VSS sg13g2_FILL8
XSTDFILL82_2149 VDD VSS sg13g2_FILL4
XSTDFILL82_2153 VDD VSS sg13g2_FILL1
XSTDFILL83_0 VDD VSS sg13g2_FILL8
XSTDFILL83_8 VDD VSS sg13g2_FILL8
XSTDFILL83_16 VDD VSS sg13g2_FILL8
XSTDFILL83_24 VDD VSS sg13g2_FILL8
XSTDFILL83_32 VDD VSS sg13g2_FILL8
XSTDFILL83_40 VDD VSS sg13g2_FILL8
XSTDFILL83_48 VDD VSS sg13g2_FILL8
XSTDFILL83_56 VDD VSS sg13g2_FILL8
XSTDFILL83_64 VDD VSS sg13g2_FILL8
XSTDFILL83_72 VDD VSS sg13g2_FILL8
XSTDFILL83_80 VDD VSS sg13g2_FILL8
XSTDFILL83_88 VDD VSS sg13g2_FILL8
XSTDFILL83_96 VDD VSS sg13g2_FILL8
XSTDFILL83_104 VDD VSS sg13g2_FILL8
XSTDFILL83_112 VDD VSS sg13g2_FILL8
XSTDFILL83_120 VDD VSS sg13g2_FILL8
XSTDFILL83_128 VDD VSS sg13g2_FILL4
XSTDFILL83_1085 VDD VSS sg13g2_FILL8
XSTDFILL83_1093 VDD VSS sg13g2_FILL8
XSTDFILL83_1101 VDD VSS sg13g2_FILL8
XSTDFILL83_1109 VDD VSS sg13g2_FILL8
XSTDFILL83_1117 VDD VSS sg13g2_FILL8
XSTDFILL83_1125 VDD VSS sg13g2_FILL8
XSTDFILL83_1133 VDD VSS sg13g2_FILL8
XSTDFILL83_1141 VDD VSS sg13g2_FILL8
XSTDFILL83_1149 VDD VSS sg13g2_FILL8
XSTDFILL83_1157 VDD VSS sg13g2_FILL8
XSTDFILL83_1165 VDD VSS sg13g2_FILL8
XSTDFILL83_1173 VDD VSS sg13g2_FILL8
XSTDFILL83_1181 VDD VSS sg13g2_FILL8
XSTDFILL83_1189 VDD VSS sg13g2_FILL8
XSTDFILL83_1197 VDD VSS sg13g2_FILL8
XSTDFILL83_1205 VDD VSS sg13g2_FILL8
XSTDFILL83_1213 VDD VSS sg13g2_FILL8
XSTDFILL83_1221 VDD VSS sg13g2_FILL8
XSTDFILL83_1229 VDD VSS sg13g2_FILL8
XSTDFILL83_1237 VDD VSS sg13g2_FILL8
XSTDFILL83_1245 VDD VSS sg13g2_FILL8
XSTDFILL83_1253 VDD VSS sg13g2_FILL8
XSTDFILL83_1261 VDD VSS sg13g2_FILL8
XSTDFILL83_1269 VDD VSS sg13g2_FILL8
XSTDFILL83_1277 VDD VSS sg13g2_FILL8
XSTDFILL83_1285 VDD VSS sg13g2_FILL8
XSTDFILL83_1293 VDD VSS sg13g2_FILL8
XSTDFILL83_1301 VDD VSS sg13g2_FILL8
XSTDFILL83_1309 VDD VSS sg13g2_FILL8
XSTDFILL83_1317 VDD VSS sg13g2_FILL8
XSTDFILL83_1325 VDD VSS sg13g2_FILL8
XSTDFILL83_1333 VDD VSS sg13g2_FILL8
XSTDFILL83_1341 VDD VSS sg13g2_FILL8
XSTDFILL83_1349 VDD VSS sg13g2_FILL8
XSTDFILL83_1357 VDD VSS sg13g2_FILL8
XSTDFILL83_1365 VDD VSS sg13g2_FILL8
XSTDFILL83_1373 VDD VSS sg13g2_FILL8
XSTDFILL83_1381 VDD VSS sg13g2_FILL8
XSTDFILL83_1389 VDD VSS sg13g2_FILL8
XSTDFILL83_1397 VDD VSS sg13g2_FILL8
XSTDFILL83_1405 VDD VSS sg13g2_FILL8
XSTDFILL83_1413 VDD VSS sg13g2_FILL8
XSTDFILL83_1421 VDD VSS sg13g2_FILL8
XSTDFILL83_1429 VDD VSS sg13g2_FILL8
XSTDFILL83_1437 VDD VSS sg13g2_FILL8
XSTDFILL83_1445 VDD VSS sg13g2_FILL8
XSTDFILL83_1453 VDD VSS sg13g2_FILL8
XSTDFILL83_1461 VDD VSS sg13g2_FILL8
XSTDFILL83_1469 VDD VSS sg13g2_FILL8
XSTDFILL83_1477 VDD VSS sg13g2_FILL8
XSTDFILL83_1485 VDD VSS sg13g2_FILL8
XSTDFILL83_1493 VDD VSS sg13g2_FILL8
XSTDFILL83_1501 VDD VSS sg13g2_FILL8
XSTDFILL83_1509 VDD VSS sg13g2_FILL8
XSTDFILL83_1517 VDD VSS sg13g2_FILL8
XSTDFILL83_1525 VDD VSS sg13g2_FILL8
XSTDFILL83_1533 VDD VSS sg13g2_FILL8
XSTDFILL83_1541 VDD VSS sg13g2_FILL8
XSTDFILL83_1549 VDD VSS sg13g2_FILL8
XSTDFILL83_1557 VDD VSS sg13g2_FILL8
XSTDFILL83_1565 VDD VSS sg13g2_FILL8
XSTDFILL83_1573 VDD VSS sg13g2_FILL8
XSTDFILL83_1581 VDD VSS sg13g2_FILL8
XSTDFILL83_1589 VDD VSS sg13g2_FILL8
XSTDFILL83_1597 VDD VSS sg13g2_FILL8
XSTDFILL83_1605 VDD VSS sg13g2_FILL8
XSTDFILL83_1613 VDD VSS sg13g2_FILL8
XSTDFILL83_1621 VDD VSS sg13g2_FILL8
XSTDFILL83_1629 VDD VSS sg13g2_FILL8
XSTDFILL83_1637 VDD VSS sg13g2_FILL8
XSTDFILL83_1645 VDD VSS sg13g2_FILL8
XSTDFILL83_1653 VDD VSS sg13g2_FILL8
XSTDFILL83_1661 VDD VSS sg13g2_FILL8
XSTDFILL83_1669 VDD VSS sg13g2_FILL8
XSTDFILL83_1677 VDD VSS sg13g2_FILL8
XSTDFILL83_1685 VDD VSS sg13g2_FILL8
XSTDFILL83_1693 VDD VSS sg13g2_FILL8
XSTDFILL83_1701 VDD VSS sg13g2_FILL8
XSTDFILL83_1709 VDD VSS sg13g2_FILL8
XSTDFILL83_1717 VDD VSS sg13g2_FILL8
XSTDFILL83_1725 VDD VSS sg13g2_FILL8
XSTDFILL83_1733 VDD VSS sg13g2_FILL8
XSTDFILL83_1741 VDD VSS sg13g2_FILL8
XSTDFILL83_1749 VDD VSS sg13g2_FILL8
XSTDFILL83_1757 VDD VSS sg13g2_FILL8
XSTDFILL83_1765 VDD VSS sg13g2_FILL8
XSTDFILL83_1773 VDD VSS sg13g2_FILL8
XSTDFILL83_1781 VDD VSS sg13g2_FILL8
XSTDFILL83_1789 VDD VSS sg13g2_FILL8
XSTDFILL83_1797 VDD VSS sg13g2_FILL8
XSTDFILL83_1805 VDD VSS sg13g2_FILL8
XSTDFILL83_1813 VDD VSS sg13g2_FILL8
XSTDFILL83_1821 VDD VSS sg13g2_FILL8
XSTDFILL83_1829 VDD VSS sg13g2_FILL8
XSTDFILL83_1837 VDD VSS sg13g2_FILL8
XSTDFILL83_1845 VDD VSS sg13g2_FILL8
XSTDFILL83_1853 VDD VSS sg13g2_FILL8
XSTDFILL83_1861 VDD VSS sg13g2_FILL8
XSTDFILL83_1869 VDD VSS sg13g2_FILL8
XSTDFILL83_1877 VDD VSS sg13g2_FILL8
XSTDFILL83_1885 VDD VSS sg13g2_FILL8
XSTDFILL83_1893 VDD VSS sg13g2_FILL8
XSTDFILL83_1901 VDD VSS sg13g2_FILL8
XSTDFILL83_1909 VDD VSS sg13g2_FILL8
XSTDFILL83_1917 VDD VSS sg13g2_FILL8
XSTDFILL83_1925 VDD VSS sg13g2_FILL8
XSTDFILL83_1933 VDD VSS sg13g2_FILL8
XSTDFILL83_1941 VDD VSS sg13g2_FILL8
XSTDFILL83_1949 VDD VSS sg13g2_FILL8
XSTDFILL83_1957 VDD VSS sg13g2_FILL8
XSTDFILL83_1965 VDD VSS sg13g2_FILL8
XSTDFILL83_1973 VDD VSS sg13g2_FILL8
XSTDFILL83_1981 VDD VSS sg13g2_FILL8
XSTDFILL83_1989 VDD VSS sg13g2_FILL8
XSTDFILL83_1997 VDD VSS sg13g2_FILL8
XSTDFILL83_2005 VDD VSS sg13g2_FILL8
XSTDFILL83_2013 VDD VSS sg13g2_FILL8
XSTDFILL83_2021 VDD VSS sg13g2_FILL8
XSTDFILL83_2029 VDD VSS sg13g2_FILL8
XSTDFILL83_2037 VDD VSS sg13g2_FILL8
XSTDFILL83_2045 VDD VSS sg13g2_FILL8
XSTDFILL83_2053 VDD VSS sg13g2_FILL8
XSTDFILL83_2061 VDD VSS sg13g2_FILL8
XSTDFILL83_2069 VDD VSS sg13g2_FILL8
XSTDFILL83_2077 VDD VSS sg13g2_FILL8
XSTDFILL83_2085 VDD VSS sg13g2_FILL8
XSTDFILL83_2093 VDD VSS sg13g2_FILL8
XSTDFILL83_2101 VDD VSS sg13g2_FILL8
XSTDFILL83_2109 VDD VSS sg13g2_FILL8
XSTDFILL83_2117 VDD VSS sg13g2_FILL8
XSTDFILL83_2125 VDD VSS sg13g2_FILL8
XSTDFILL83_2133 VDD VSS sg13g2_FILL8
XSTDFILL83_2141 VDD VSS sg13g2_FILL8
XSTDFILL83_2149 VDD VSS sg13g2_FILL4
XSTDFILL83_2153 VDD VSS sg13g2_FILL1
XSTDFILL84_0 VDD VSS sg13g2_FILL8
XSTDFILL84_8 VDD VSS sg13g2_FILL8
XSTDFILL84_16 VDD VSS sg13g2_FILL8
XSTDFILL84_24 VDD VSS sg13g2_FILL8
XSTDFILL84_32 VDD VSS sg13g2_FILL8
XSTDFILL84_40 VDD VSS sg13g2_FILL8
XSTDFILL84_48 VDD VSS sg13g2_FILL8
XSTDFILL84_56 VDD VSS sg13g2_FILL8
XSTDFILL84_64 VDD VSS sg13g2_FILL8
XSTDFILL84_72 VDD VSS sg13g2_FILL8
XSTDFILL84_80 VDD VSS sg13g2_FILL8
XSTDFILL84_88 VDD VSS sg13g2_FILL8
XSTDFILL84_96 VDD VSS sg13g2_FILL8
XSTDFILL84_104 VDD VSS sg13g2_FILL8
XSTDFILL84_112 VDD VSS sg13g2_FILL8
XSTDFILL84_120 VDD VSS sg13g2_FILL8
XSTDFILL84_128 VDD VSS sg13g2_FILL4
XSTDFILL84_1085 VDD VSS sg13g2_FILL8
XSTDFILL84_1093 VDD VSS sg13g2_FILL8
XSTDFILL84_1101 VDD VSS sg13g2_FILL8
XSTDFILL84_1109 VDD VSS sg13g2_FILL8
XSTDFILL84_1117 VDD VSS sg13g2_FILL8
XSTDFILL84_1125 VDD VSS sg13g2_FILL8
XSTDFILL84_1133 VDD VSS sg13g2_FILL8
XSTDFILL84_1141 VDD VSS sg13g2_FILL8
XSTDFILL84_1149 VDD VSS sg13g2_FILL8
XSTDFILL84_1157 VDD VSS sg13g2_FILL8
XSTDFILL84_1165 VDD VSS sg13g2_FILL8
XSTDFILL84_1173 VDD VSS sg13g2_FILL8
XSTDFILL84_1181 VDD VSS sg13g2_FILL8
XSTDFILL84_1189 VDD VSS sg13g2_FILL8
XSTDFILL84_1197 VDD VSS sg13g2_FILL8
XSTDFILL84_1205 VDD VSS sg13g2_FILL8
XSTDFILL84_1213 VDD VSS sg13g2_FILL8
XSTDFILL84_1221 VDD VSS sg13g2_FILL8
XSTDFILL84_1229 VDD VSS sg13g2_FILL8
XSTDFILL84_1237 VDD VSS sg13g2_FILL8
XSTDFILL84_1245 VDD VSS sg13g2_FILL8
XSTDFILL84_1253 VDD VSS sg13g2_FILL8
XSTDFILL84_1261 VDD VSS sg13g2_FILL8
XSTDFILL84_1269 VDD VSS sg13g2_FILL8
XSTDFILL84_1277 VDD VSS sg13g2_FILL8
XSTDFILL84_1285 VDD VSS sg13g2_FILL8
XSTDFILL84_1293 VDD VSS sg13g2_FILL8
XSTDFILL84_1301 VDD VSS sg13g2_FILL8
XSTDFILL84_1309 VDD VSS sg13g2_FILL8
XSTDFILL84_1317 VDD VSS sg13g2_FILL8
XSTDFILL84_1325 VDD VSS sg13g2_FILL8
XSTDFILL84_1333 VDD VSS sg13g2_FILL8
XSTDFILL84_1341 VDD VSS sg13g2_FILL8
XSTDFILL84_1349 VDD VSS sg13g2_FILL8
XSTDFILL84_1357 VDD VSS sg13g2_FILL8
XSTDFILL84_1365 VDD VSS sg13g2_FILL8
XSTDFILL84_1373 VDD VSS sg13g2_FILL8
XSTDFILL84_1381 VDD VSS sg13g2_FILL8
XSTDFILL84_1389 VDD VSS sg13g2_FILL8
XSTDFILL84_1397 VDD VSS sg13g2_FILL8
XSTDFILL84_1405 VDD VSS sg13g2_FILL8
XSTDFILL84_1413 VDD VSS sg13g2_FILL8
XSTDFILL84_1421 VDD VSS sg13g2_FILL8
XSTDFILL84_1429 VDD VSS sg13g2_FILL8
XSTDFILL84_1437 VDD VSS sg13g2_FILL8
XSTDFILL84_1445 VDD VSS sg13g2_FILL8
XSTDFILL84_1453 VDD VSS sg13g2_FILL8
XSTDFILL84_1461 VDD VSS sg13g2_FILL8
XSTDFILL84_1469 VDD VSS sg13g2_FILL8
XSTDFILL84_1477 VDD VSS sg13g2_FILL8
XSTDFILL84_1485 VDD VSS sg13g2_FILL8
XSTDFILL84_1493 VDD VSS sg13g2_FILL8
XSTDFILL84_1501 VDD VSS sg13g2_FILL8
XSTDFILL84_1509 VDD VSS sg13g2_FILL8
XSTDFILL84_1517 VDD VSS sg13g2_FILL8
XSTDFILL85_0 VDD VSS sg13g2_FILL8
XSTDFILL85_8 VDD VSS sg13g2_FILL8
XSTDFILL85_16 VDD VSS sg13g2_FILL8
XSTDFILL85_24 VDD VSS sg13g2_FILL8
XSTDFILL85_32 VDD VSS sg13g2_FILL8
XSTDFILL85_40 VDD VSS sg13g2_FILL8
XSTDFILL85_48 VDD VSS sg13g2_FILL8
XSTDFILL85_56 VDD VSS sg13g2_FILL8
XSTDFILL85_64 VDD VSS sg13g2_FILL8
XSTDFILL85_72 VDD VSS sg13g2_FILL8
XSTDFILL85_80 VDD VSS sg13g2_FILL8
XSTDFILL85_88 VDD VSS sg13g2_FILL8
XSTDFILL85_96 VDD VSS sg13g2_FILL8
XSTDFILL85_104 VDD VSS sg13g2_FILL8
XSTDFILL85_112 VDD VSS sg13g2_FILL8
XSTDFILL85_120 VDD VSS sg13g2_FILL8
XSTDFILL85_128 VDD VSS sg13g2_FILL4
XSTDFILL85_1085 VDD VSS sg13g2_FILL8
XSTDFILL85_1093 VDD VSS sg13g2_FILL8
XSTDFILL85_1101 VDD VSS sg13g2_FILL8
XSTDFILL85_1109 VDD VSS sg13g2_FILL8
XSTDFILL85_1117 VDD VSS sg13g2_FILL8
XSTDFILL85_1125 VDD VSS sg13g2_FILL8
XSTDFILL85_1133 VDD VSS sg13g2_FILL8
XSTDFILL85_1141 VDD VSS sg13g2_FILL8
XSTDFILL85_1149 VDD VSS sg13g2_FILL8
XSTDFILL85_1157 VDD VSS sg13g2_FILL8
XSTDFILL85_1165 VDD VSS sg13g2_FILL8
XSTDFILL85_1173 VDD VSS sg13g2_FILL8
XSTDFILL85_1181 VDD VSS sg13g2_FILL8
XSTDFILL85_1189 VDD VSS sg13g2_FILL8
XSTDFILL85_1197 VDD VSS sg13g2_FILL8
XSTDFILL85_1205 VDD VSS sg13g2_FILL8
XSTDFILL85_1213 VDD VSS sg13g2_FILL8
XSTDFILL85_1221 VDD VSS sg13g2_FILL8
XSTDFILL85_1229 VDD VSS sg13g2_FILL8
XSTDFILL85_1237 VDD VSS sg13g2_FILL8
XSTDFILL85_1245 VDD VSS sg13g2_FILL8
XSTDFILL85_1253 VDD VSS sg13g2_FILL8
XSTDFILL85_1261 VDD VSS sg13g2_FILL8
XSTDFILL85_1269 VDD VSS sg13g2_FILL8
XSTDFILL85_1277 VDD VSS sg13g2_FILL8
XSTDFILL85_1285 VDD VSS sg13g2_FILL8
XSTDFILL85_1293 VDD VSS sg13g2_FILL8
XSTDFILL85_1301 VDD VSS sg13g2_FILL8
XSTDFILL85_1309 VDD VSS sg13g2_FILL8
XSTDFILL85_1317 VDD VSS sg13g2_FILL8
XSTDFILL85_1325 VDD VSS sg13g2_FILL8
XSTDFILL85_1333 VDD VSS sg13g2_FILL8
XSTDFILL85_1341 VDD VSS sg13g2_FILL8
XSTDFILL85_1349 VDD VSS sg13g2_FILL8
XSTDFILL85_1357 VDD VSS sg13g2_FILL8
XSTDFILL85_1365 VDD VSS sg13g2_FILL8
XSTDFILL85_1373 VDD VSS sg13g2_FILL8
XSTDFILL85_1381 VDD VSS sg13g2_FILL8
XSTDFILL85_1389 VDD VSS sg13g2_FILL8
XSTDFILL85_1397 VDD VSS sg13g2_FILL8
XSTDFILL85_1405 VDD VSS sg13g2_FILL8
XSTDFILL85_1413 VDD VSS sg13g2_FILL8
XSTDFILL85_1421 VDD VSS sg13g2_FILL8
XSTDFILL85_1429 VDD VSS sg13g2_FILL8
XSTDFILL85_1437 VDD VSS sg13g2_FILL8
XSTDFILL85_1445 VDD VSS sg13g2_FILL8
XSTDFILL85_1453 VDD VSS sg13g2_FILL8
XSTDFILL85_1461 VDD VSS sg13g2_FILL8
XSTDFILL85_1469 VDD VSS sg13g2_FILL8
XSTDFILL85_1477 VDD VSS sg13g2_FILL8
XSTDFILL85_1485 VDD VSS sg13g2_FILL8
XSTDFILL85_1493 VDD VSS sg13g2_FILL8
XSTDFILL85_1501 VDD VSS sg13g2_FILL8
XSTDFILL85_1509 VDD VSS sg13g2_FILL8
XSTDFILL85_1517 VDD VSS sg13g2_FILL8
XSTDFILL86_0 VDD VSS sg13g2_FILL8
XSTDFILL86_8 VDD VSS sg13g2_FILL8
XSTDFILL86_16 VDD VSS sg13g2_FILL8
XSTDFILL86_24 VDD VSS sg13g2_FILL8
XSTDFILL86_32 VDD VSS sg13g2_FILL8
XSTDFILL86_40 VDD VSS sg13g2_FILL8
XSTDFILL86_48 VDD VSS sg13g2_FILL8
XSTDFILL86_56 VDD VSS sg13g2_FILL8
XSTDFILL86_64 VDD VSS sg13g2_FILL8
XSTDFILL86_72 VDD VSS sg13g2_FILL8
XSTDFILL86_80 VDD VSS sg13g2_FILL8
XSTDFILL86_88 VDD VSS sg13g2_FILL8
XSTDFILL86_96 VDD VSS sg13g2_FILL8
XSTDFILL86_104 VDD VSS sg13g2_FILL8
XSTDFILL86_112 VDD VSS sg13g2_FILL8
XSTDFILL86_120 VDD VSS sg13g2_FILL8
XSTDFILL86_128 VDD VSS sg13g2_FILL4
XSTDFILL86_1085 VDD VSS sg13g2_FILL8
XSTDFILL86_1093 VDD VSS sg13g2_FILL8
XSTDFILL86_1101 VDD VSS sg13g2_FILL8
XSTDFILL86_1109 VDD VSS sg13g2_FILL8
XSTDFILL86_1117 VDD VSS sg13g2_FILL8
XSTDFILL86_1125 VDD VSS sg13g2_FILL8
XSTDFILL86_1133 VDD VSS sg13g2_FILL8
XSTDFILL86_1141 VDD VSS sg13g2_FILL8
XSTDFILL86_1149 VDD VSS sg13g2_FILL8
XSTDFILL86_1157 VDD VSS sg13g2_FILL8
XSTDFILL86_1165 VDD VSS sg13g2_FILL8
XSTDFILL86_1173 VDD VSS sg13g2_FILL8
XSTDFILL86_1181 VDD VSS sg13g2_FILL8
XSTDFILL86_1189 VDD VSS sg13g2_FILL8
XSTDFILL86_1197 VDD VSS sg13g2_FILL8
XSTDFILL86_1205 VDD VSS sg13g2_FILL8
XSTDFILL86_1213 VDD VSS sg13g2_FILL8
XSTDFILL86_1221 VDD VSS sg13g2_FILL8
XSTDFILL86_1229 VDD VSS sg13g2_FILL8
XSTDFILL86_1237 VDD VSS sg13g2_FILL8
XSTDFILL86_1245 VDD VSS sg13g2_FILL8
XSTDFILL86_1253 VDD VSS sg13g2_FILL8
XSTDFILL86_1261 VDD VSS sg13g2_FILL8
XSTDFILL86_1269 VDD VSS sg13g2_FILL8
XSTDFILL86_1277 VDD VSS sg13g2_FILL8
XSTDFILL86_1285 VDD VSS sg13g2_FILL8
XSTDFILL86_1293 VDD VSS sg13g2_FILL8
XSTDFILL86_1301 VDD VSS sg13g2_FILL8
XSTDFILL86_1309 VDD VSS sg13g2_FILL8
XSTDFILL86_1317 VDD VSS sg13g2_FILL8
XSTDFILL86_1325 VDD VSS sg13g2_FILL8
XSTDFILL86_1333 VDD VSS sg13g2_FILL8
XSTDFILL86_1341 VDD VSS sg13g2_FILL8
XSTDFILL86_1349 VDD VSS sg13g2_FILL8
XSTDFILL86_1357 VDD VSS sg13g2_FILL8
XSTDFILL86_1365 VDD VSS sg13g2_FILL8
XSTDFILL86_1373 VDD VSS sg13g2_FILL8
XSTDFILL86_1381 VDD VSS sg13g2_FILL8
XSTDFILL86_1389 VDD VSS sg13g2_FILL8
XSTDFILL86_1397 VDD VSS sg13g2_FILL8
XSTDFILL86_1405 VDD VSS sg13g2_FILL8
XSTDFILL86_1413 VDD VSS sg13g2_FILL8
XSTDFILL86_1421 VDD VSS sg13g2_FILL8
XSTDFILL86_1429 VDD VSS sg13g2_FILL8
XSTDFILL86_1437 VDD VSS sg13g2_FILL8
XSTDFILL86_1445 VDD VSS sg13g2_FILL8
XSTDFILL86_1453 VDD VSS sg13g2_FILL8
XSTDFILL86_1461 VDD VSS sg13g2_FILL8
XSTDFILL86_1469 VDD VSS sg13g2_FILL8
XSTDFILL86_1477 VDD VSS sg13g2_FILL8
XSTDFILL86_1485 VDD VSS sg13g2_FILL8
XSTDFILL86_1493 VDD VSS sg13g2_FILL8
XSTDFILL86_1501 VDD VSS sg13g2_FILL8
XSTDFILL86_1509 VDD VSS sg13g2_FILL8
XSTDFILL86_1517 VDD VSS sg13g2_FILL8
XSTDFILL87_0 VDD VSS sg13g2_FILL8
XSTDFILL87_8 VDD VSS sg13g2_FILL8
XSTDFILL87_16 VDD VSS sg13g2_FILL8
XSTDFILL87_24 VDD VSS sg13g2_FILL8
XSTDFILL87_32 VDD VSS sg13g2_FILL8
XSTDFILL87_40 VDD VSS sg13g2_FILL8
XSTDFILL87_48 VDD VSS sg13g2_FILL8
XSTDFILL87_56 VDD VSS sg13g2_FILL8
XSTDFILL87_64 VDD VSS sg13g2_FILL8
XSTDFILL87_72 VDD VSS sg13g2_FILL8
XSTDFILL87_80 VDD VSS sg13g2_FILL8
XSTDFILL87_88 VDD VSS sg13g2_FILL8
XSTDFILL87_96 VDD VSS sg13g2_FILL8
XSTDFILL87_104 VDD VSS sg13g2_FILL8
XSTDFILL87_112 VDD VSS sg13g2_FILL8
XSTDFILL87_120 VDD VSS sg13g2_FILL8
XSTDFILL87_128 VDD VSS sg13g2_FILL4
XSTDFILL87_1085 VDD VSS sg13g2_FILL8
XSTDFILL87_1093 VDD VSS sg13g2_FILL8
XSTDFILL87_1101 VDD VSS sg13g2_FILL8
XSTDFILL87_1109 VDD VSS sg13g2_FILL8
XSTDFILL87_1117 VDD VSS sg13g2_FILL8
XSTDFILL87_1125 VDD VSS sg13g2_FILL8
XSTDFILL87_1133 VDD VSS sg13g2_FILL8
XSTDFILL87_1141 VDD VSS sg13g2_FILL8
XSTDFILL87_1149 VDD VSS sg13g2_FILL8
XSTDFILL87_1157 VDD VSS sg13g2_FILL8
XSTDFILL87_1165 VDD VSS sg13g2_FILL8
XSTDFILL87_1173 VDD VSS sg13g2_FILL8
XSTDFILL87_1181 VDD VSS sg13g2_FILL8
XSTDFILL87_1189 VDD VSS sg13g2_FILL8
XSTDFILL87_1197 VDD VSS sg13g2_FILL8
XSTDFILL87_1205 VDD VSS sg13g2_FILL8
XSTDFILL87_1213 VDD VSS sg13g2_FILL8
XSTDFILL87_1221 VDD VSS sg13g2_FILL8
XSTDFILL87_1229 VDD VSS sg13g2_FILL8
XSTDFILL87_1237 VDD VSS sg13g2_FILL8
XSTDFILL87_1245 VDD VSS sg13g2_FILL8
XSTDFILL87_1253 VDD VSS sg13g2_FILL8
XSTDFILL87_1261 VDD VSS sg13g2_FILL8
XSTDFILL87_1269 VDD VSS sg13g2_FILL8
XSTDFILL87_1277 VDD VSS sg13g2_FILL8
XSTDFILL87_1285 VDD VSS sg13g2_FILL8
XSTDFILL87_1293 VDD VSS sg13g2_FILL8
XSTDFILL87_1301 VDD VSS sg13g2_FILL8
XSTDFILL87_1309 VDD VSS sg13g2_FILL8
XSTDFILL87_1317 VDD VSS sg13g2_FILL8
XSTDFILL87_1325 VDD VSS sg13g2_FILL8
XSTDFILL87_1333 VDD VSS sg13g2_FILL8
XSTDFILL87_1341 VDD VSS sg13g2_FILL8
XSTDFILL87_1349 VDD VSS sg13g2_FILL8
XSTDFILL87_1357 VDD VSS sg13g2_FILL8
XSTDFILL87_1365 VDD VSS sg13g2_FILL8
XSTDFILL87_1373 VDD VSS sg13g2_FILL8
XSTDFILL87_1381 VDD VSS sg13g2_FILL8
XSTDFILL87_1389 VDD VSS sg13g2_FILL8
XSTDFILL87_1397 VDD VSS sg13g2_FILL8
XSTDFILL87_1405 VDD VSS sg13g2_FILL8
XSTDFILL87_1413 VDD VSS sg13g2_FILL8
XSTDFILL87_1421 VDD VSS sg13g2_FILL8
XSTDFILL87_1429 VDD VSS sg13g2_FILL8
XSTDFILL87_1437 VDD VSS sg13g2_FILL8
XSTDFILL87_1445 VDD VSS sg13g2_FILL8
XSTDFILL87_1453 VDD VSS sg13g2_FILL8
XSTDFILL87_1461 VDD VSS sg13g2_FILL8
XSTDFILL87_1469 VDD VSS sg13g2_FILL8
XSTDFILL87_1477 VDD VSS sg13g2_FILL8
XSTDFILL87_1485 VDD VSS sg13g2_FILL8
XSTDFILL87_1493 VDD VSS sg13g2_FILL8
XSTDFILL87_1501 VDD VSS sg13g2_FILL8
XSTDFILL87_1509 VDD VSS sg13g2_FILL8
XSTDFILL87_1517 VDD VSS sg13g2_FILL8
XSTDFILL88_0 VDD VSS sg13g2_FILL8
XSTDFILL88_8 VDD VSS sg13g2_FILL8
XSTDFILL88_16 VDD VSS sg13g2_FILL8
XSTDFILL88_24 VDD VSS sg13g2_FILL8
XSTDFILL88_32 VDD VSS sg13g2_FILL8
XSTDFILL88_40 VDD VSS sg13g2_FILL8
XSTDFILL88_48 VDD VSS sg13g2_FILL8
XSTDFILL88_56 VDD VSS sg13g2_FILL8
XSTDFILL88_64 VDD VSS sg13g2_FILL8
XSTDFILL88_72 VDD VSS sg13g2_FILL8
XSTDFILL88_80 VDD VSS sg13g2_FILL8
XSTDFILL88_88 VDD VSS sg13g2_FILL8
XSTDFILL88_96 VDD VSS sg13g2_FILL8
XSTDFILL88_104 VDD VSS sg13g2_FILL8
XSTDFILL88_112 VDD VSS sg13g2_FILL8
XSTDFILL88_120 VDD VSS sg13g2_FILL8
XSTDFILL88_128 VDD VSS sg13g2_FILL4
XSTDFILL88_1085 VDD VSS sg13g2_FILL8
XSTDFILL88_1093 VDD VSS sg13g2_FILL8
XSTDFILL88_1101 VDD VSS sg13g2_FILL8
XSTDFILL88_1109 VDD VSS sg13g2_FILL8
XSTDFILL88_1117 VDD VSS sg13g2_FILL8
XSTDFILL88_1125 VDD VSS sg13g2_FILL8
XSTDFILL88_1133 VDD VSS sg13g2_FILL8
XSTDFILL88_1141 VDD VSS sg13g2_FILL8
XSTDFILL88_1149 VDD VSS sg13g2_FILL8
XSTDFILL88_1157 VDD VSS sg13g2_FILL8
XSTDFILL88_1165 VDD VSS sg13g2_FILL8
XSTDFILL88_1173 VDD VSS sg13g2_FILL8
XSTDFILL88_1181 VDD VSS sg13g2_FILL8
XSTDFILL88_1189 VDD VSS sg13g2_FILL8
XSTDFILL88_1197 VDD VSS sg13g2_FILL8
XSTDFILL88_1205 VDD VSS sg13g2_FILL8
XSTDFILL88_1213 VDD VSS sg13g2_FILL8
XSTDFILL88_1221 VDD VSS sg13g2_FILL8
XSTDFILL88_1229 VDD VSS sg13g2_FILL8
XSTDFILL88_1237 VDD VSS sg13g2_FILL8
XSTDFILL88_1245 VDD VSS sg13g2_FILL8
XSTDFILL88_1253 VDD VSS sg13g2_FILL8
XSTDFILL88_1261 VDD VSS sg13g2_FILL8
XSTDFILL88_1269 VDD VSS sg13g2_FILL8
XSTDFILL88_1277 VDD VSS sg13g2_FILL8
XSTDFILL88_1285 VDD VSS sg13g2_FILL8
XSTDFILL88_1293 VDD VSS sg13g2_FILL8
XSTDFILL88_1301 VDD VSS sg13g2_FILL8
XSTDFILL88_1309 VDD VSS sg13g2_FILL8
XSTDFILL88_1317 VDD VSS sg13g2_FILL8
XSTDFILL88_1325 VDD VSS sg13g2_FILL8
XSTDFILL88_1333 VDD VSS sg13g2_FILL8
XSTDFILL88_1341 VDD VSS sg13g2_FILL8
XSTDFILL88_1349 VDD VSS sg13g2_FILL8
XSTDFILL88_1357 VDD VSS sg13g2_FILL8
XSTDFILL88_1365 VDD VSS sg13g2_FILL8
XSTDFILL88_1373 VDD VSS sg13g2_FILL8
XSTDFILL88_1381 VDD VSS sg13g2_FILL8
XSTDFILL88_1389 VDD VSS sg13g2_FILL8
XSTDFILL88_1397 VDD VSS sg13g2_FILL8
XSTDFILL88_1405 VDD VSS sg13g2_FILL8
XSTDFILL88_1413 VDD VSS sg13g2_FILL8
XSTDFILL88_1421 VDD VSS sg13g2_FILL8
XSTDFILL88_1429 VDD VSS sg13g2_FILL8
XSTDFILL88_1437 VDD VSS sg13g2_FILL8
XSTDFILL88_1445 VDD VSS sg13g2_FILL8
XSTDFILL88_1453 VDD VSS sg13g2_FILL8
XSTDFILL88_1461 VDD VSS sg13g2_FILL8
XSTDFILL88_1469 VDD VSS sg13g2_FILL8
XSTDFILL88_1477 VDD VSS sg13g2_FILL8
XSTDFILL88_1485 VDD VSS sg13g2_FILL8
XSTDFILL88_1493 VDD VSS sg13g2_FILL8
XSTDFILL88_1501 VDD VSS sg13g2_FILL8
XSTDFILL88_1509 VDD VSS sg13g2_FILL8
XSTDFILL88_1517 VDD VSS sg13g2_FILL8
XSTDFILL89_0 VDD VSS sg13g2_FILL8
XSTDFILL89_8 VDD VSS sg13g2_FILL8
XSTDFILL89_16 VDD VSS sg13g2_FILL8
XSTDFILL89_24 VDD VSS sg13g2_FILL8
XSTDFILL89_32 VDD VSS sg13g2_FILL8
XSTDFILL89_40 VDD VSS sg13g2_FILL8
XSTDFILL89_48 VDD VSS sg13g2_FILL8
XSTDFILL89_56 VDD VSS sg13g2_FILL8
XSTDFILL89_64 VDD VSS sg13g2_FILL8
XSTDFILL89_72 VDD VSS sg13g2_FILL8
XSTDFILL89_80 VDD VSS sg13g2_FILL8
XSTDFILL89_88 VDD VSS sg13g2_FILL8
XSTDFILL89_96 VDD VSS sg13g2_FILL8
XSTDFILL89_104 VDD VSS sg13g2_FILL8
XSTDFILL89_112 VDD VSS sg13g2_FILL8
XSTDFILL89_120 VDD VSS sg13g2_FILL8
XSTDFILL89_128 VDD VSS sg13g2_FILL4
XSTDFILL89_1085 VDD VSS sg13g2_FILL8
XSTDFILL89_1093 VDD VSS sg13g2_FILL8
XSTDFILL89_1101 VDD VSS sg13g2_FILL8
XSTDFILL89_1109 VDD VSS sg13g2_FILL8
XSTDFILL89_1117 VDD VSS sg13g2_FILL8
XSTDFILL89_1125 VDD VSS sg13g2_FILL8
XSTDFILL89_1133 VDD VSS sg13g2_FILL8
XSTDFILL89_1141 VDD VSS sg13g2_FILL8
XSTDFILL89_1149 VDD VSS sg13g2_FILL8
XSTDFILL89_1157 VDD VSS sg13g2_FILL8
XSTDFILL89_1165 VDD VSS sg13g2_FILL8
XSTDFILL89_1173 VDD VSS sg13g2_FILL8
XSTDFILL89_1181 VDD VSS sg13g2_FILL8
XSTDFILL89_1189 VDD VSS sg13g2_FILL8
XSTDFILL89_1197 VDD VSS sg13g2_FILL8
XSTDFILL89_1205 VDD VSS sg13g2_FILL8
XSTDFILL89_1213 VDD VSS sg13g2_FILL8
XSTDFILL89_1221 VDD VSS sg13g2_FILL8
XSTDFILL89_1229 VDD VSS sg13g2_FILL8
XSTDFILL89_1237 VDD VSS sg13g2_FILL8
XSTDFILL89_1245 VDD VSS sg13g2_FILL8
XSTDFILL89_1253 VDD VSS sg13g2_FILL8
XSTDFILL89_1261 VDD VSS sg13g2_FILL8
XSTDFILL89_1269 VDD VSS sg13g2_FILL8
XSTDFILL89_1277 VDD VSS sg13g2_FILL8
XSTDFILL89_1285 VDD VSS sg13g2_FILL8
XSTDFILL89_1293 VDD VSS sg13g2_FILL8
XSTDFILL89_1301 VDD VSS sg13g2_FILL8
XSTDFILL89_1309 VDD VSS sg13g2_FILL8
XSTDFILL89_1317 VDD VSS sg13g2_FILL8
XSTDFILL89_1325 VDD VSS sg13g2_FILL8
XSTDFILL89_1333 VDD VSS sg13g2_FILL8
XSTDFILL89_1341 VDD VSS sg13g2_FILL8
XSTDFILL89_1349 VDD VSS sg13g2_FILL8
XSTDFILL89_1357 VDD VSS sg13g2_FILL8
XSTDFILL89_1365 VDD VSS sg13g2_FILL8
XSTDFILL89_1373 VDD VSS sg13g2_FILL8
XSTDFILL89_1381 VDD VSS sg13g2_FILL8
XSTDFILL89_1389 VDD VSS sg13g2_FILL8
XSTDFILL89_1397 VDD VSS sg13g2_FILL8
XSTDFILL89_1405 VDD VSS sg13g2_FILL8
XSTDFILL89_1413 VDD VSS sg13g2_FILL8
XSTDFILL89_1421 VDD VSS sg13g2_FILL8
XSTDFILL89_1429 VDD VSS sg13g2_FILL8
XSTDFILL89_1437 VDD VSS sg13g2_FILL8
XSTDFILL89_1445 VDD VSS sg13g2_FILL8
XSTDFILL89_1453 VDD VSS sg13g2_FILL8
XSTDFILL89_1461 VDD VSS sg13g2_FILL8
XSTDFILL89_1469 VDD VSS sg13g2_FILL8
XSTDFILL89_1477 VDD VSS sg13g2_FILL8
XSTDFILL89_1485 VDD VSS sg13g2_FILL8
XSTDFILL89_1493 VDD VSS sg13g2_FILL8
XSTDFILL89_1501 VDD VSS sg13g2_FILL8
XSTDFILL89_1509 VDD VSS sg13g2_FILL8
XSTDFILL89_1517 VDD VSS sg13g2_FILL8
XSTDFILL90_0 VDD VSS sg13g2_FILL8
XSTDFILL90_8 VDD VSS sg13g2_FILL8
XSTDFILL90_16 VDD VSS sg13g2_FILL8
XSTDFILL90_24 VDD VSS sg13g2_FILL8
XSTDFILL90_32 VDD VSS sg13g2_FILL8
XSTDFILL90_40 VDD VSS sg13g2_FILL8
XSTDFILL90_48 VDD VSS sg13g2_FILL8
XSTDFILL90_56 VDD VSS sg13g2_FILL8
XSTDFILL90_64 VDD VSS sg13g2_FILL8
XSTDFILL90_72 VDD VSS sg13g2_FILL8
XSTDFILL90_80 VDD VSS sg13g2_FILL8
XSTDFILL90_88 VDD VSS sg13g2_FILL8
XSTDFILL90_96 VDD VSS sg13g2_FILL8
XSTDFILL90_104 VDD VSS sg13g2_FILL8
XSTDFILL90_112 VDD VSS sg13g2_FILL8
XSTDFILL90_120 VDD VSS sg13g2_FILL8
XSTDFILL90_128 VDD VSS sg13g2_FILL4
XSTDFILL90_1085 VDD VSS sg13g2_FILL8
XSTDFILL90_1093 VDD VSS sg13g2_FILL8
XSTDFILL90_1101 VDD VSS sg13g2_FILL8
XSTDFILL90_1109 VDD VSS sg13g2_FILL8
XSTDFILL90_1117 VDD VSS sg13g2_FILL8
XSTDFILL90_1125 VDD VSS sg13g2_FILL8
XSTDFILL90_1133 VDD VSS sg13g2_FILL8
XSTDFILL90_1141 VDD VSS sg13g2_FILL8
XSTDFILL90_1149 VDD VSS sg13g2_FILL8
XSTDFILL90_1157 VDD VSS sg13g2_FILL8
XSTDFILL90_1165 VDD VSS sg13g2_FILL8
XSTDFILL90_1173 VDD VSS sg13g2_FILL8
XSTDFILL90_1181 VDD VSS sg13g2_FILL8
XSTDFILL90_1189 VDD VSS sg13g2_FILL8
XSTDFILL90_1197 VDD VSS sg13g2_FILL8
XSTDFILL90_1205 VDD VSS sg13g2_FILL8
XSTDFILL90_1213 VDD VSS sg13g2_FILL8
XSTDFILL90_1221 VDD VSS sg13g2_FILL8
XSTDFILL90_1229 VDD VSS sg13g2_FILL8
XSTDFILL90_1237 VDD VSS sg13g2_FILL8
XSTDFILL90_1245 VDD VSS sg13g2_FILL8
XSTDFILL90_1253 VDD VSS sg13g2_FILL8
XSTDFILL90_1261 VDD VSS sg13g2_FILL8
XSTDFILL90_1269 VDD VSS sg13g2_FILL8
XSTDFILL90_1277 VDD VSS sg13g2_FILL8
XSTDFILL90_1285 VDD VSS sg13g2_FILL8
XSTDFILL90_1293 VDD VSS sg13g2_FILL8
XSTDFILL90_1301 VDD VSS sg13g2_FILL8
XSTDFILL90_1309 VDD VSS sg13g2_FILL8
XSTDFILL90_1317 VDD VSS sg13g2_FILL8
XSTDFILL90_1325 VDD VSS sg13g2_FILL8
XSTDFILL90_1333 VDD VSS sg13g2_FILL8
XSTDFILL90_1341 VDD VSS sg13g2_FILL8
XSTDFILL90_1349 VDD VSS sg13g2_FILL8
XSTDFILL90_1357 VDD VSS sg13g2_FILL8
XSTDFILL90_1365 VDD VSS sg13g2_FILL8
XSTDFILL90_1373 VDD VSS sg13g2_FILL8
XSTDFILL90_1381 VDD VSS sg13g2_FILL8
XSTDFILL90_1389 VDD VSS sg13g2_FILL8
XSTDFILL90_1397 VDD VSS sg13g2_FILL8
XSTDFILL90_1405 VDD VSS sg13g2_FILL8
XSTDFILL90_1413 VDD VSS sg13g2_FILL8
XSTDFILL90_1421 VDD VSS sg13g2_FILL8
XSTDFILL90_1429 VDD VSS sg13g2_FILL8
XSTDFILL90_1437 VDD VSS sg13g2_FILL8
XSTDFILL90_1445 VDD VSS sg13g2_FILL8
XSTDFILL90_1453 VDD VSS sg13g2_FILL8
XSTDFILL90_1461 VDD VSS sg13g2_FILL8
XSTDFILL90_1469 VDD VSS sg13g2_FILL8
XSTDFILL90_1477 VDD VSS sg13g2_FILL8
XSTDFILL90_1485 VDD VSS sg13g2_FILL8
XSTDFILL90_1493 VDD VSS sg13g2_FILL8
XSTDFILL90_1501 VDD VSS sg13g2_FILL8
XSTDFILL90_1509 VDD VSS sg13g2_FILL8
XSTDFILL90_1517 VDD VSS sg13g2_FILL8
XSTDFILL91_0 VDD VSS sg13g2_FILL8
XSTDFILL91_8 VDD VSS sg13g2_FILL8
XSTDFILL91_16 VDD VSS sg13g2_FILL8
XSTDFILL91_24 VDD VSS sg13g2_FILL8
XSTDFILL91_32 VDD VSS sg13g2_FILL8
XSTDFILL91_40 VDD VSS sg13g2_FILL8
XSTDFILL91_48 VDD VSS sg13g2_FILL8
XSTDFILL91_56 VDD VSS sg13g2_FILL8
XSTDFILL91_64 VDD VSS sg13g2_FILL8
XSTDFILL91_72 VDD VSS sg13g2_FILL8
XSTDFILL91_80 VDD VSS sg13g2_FILL8
XSTDFILL91_88 VDD VSS sg13g2_FILL8
XSTDFILL91_96 VDD VSS sg13g2_FILL8
XSTDFILL91_104 VDD VSS sg13g2_FILL8
XSTDFILL91_112 VDD VSS sg13g2_FILL8
XSTDFILL91_120 VDD VSS sg13g2_FILL8
XSTDFILL91_128 VDD VSS sg13g2_FILL4
XSTDFILL91_1085 VDD VSS sg13g2_FILL8
XSTDFILL91_1093 VDD VSS sg13g2_FILL8
XSTDFILL91_1101 VDD VSS sg13g2_FILL8
XSTDFILL91_1109 VDD VSS sg13g2_FILL8
XSTDFILL91_1117 VDD VSS sg13g2_FILL8
XSTDFILL91_1125 VDD VSS sg13g2_FILL8
XSTDFILL91_1133 VDD VSS sg13g2_FILL8
XSTDFILL91_1141 VDD VSS sg13g2_FILL8
XSTDFILL91_1149 VDD VSS sg13g2_FILL8
XSTDFILL91_1157 VDD VSS sg13g2_FILL8
XSTDFILL91_1165 VDD VSS sg13g2_FILL8
XSTDFILL91_1173 VDD VSS sg13g2_FILL8
XSTDFILL91_1181 VDD VSS sg13g2_FILL8
XSTDFILL91_1189 VDD VSS sg13g2_FILL8
XSTDFILL91_1197 VDD VSS sg13g2_FILL8
XSTDFILL91_1205 VDD VSS sg13g2_FILL8
XSTDFILL91_1213 VDD VSS sg13g2_FILL8
XSTDFILL91_1221 VDD VSS sg13g2_FILL8
XSTDFILL91_1229 VDD VSS sg13g2_FILL8
XSTDFILL91_1237 VDD VSS sg13g2_FILL8
XSTDFILL91_1245 VDD VSS sg13g2_FILL8
XSTDFILL91_1253 VDD VSS sg13g2_FILL8
XSTDFILL91_1261 VDD VSS sg13g2_FILL8
XSTDFILL91_1269 VDD VSS sg13g2_FILL8
XSTDFILL91_1277 VDD VSS sg13g2_FILL8
XSTDFILL91_1285 VDD VSS sg13g2_FILL8
XSTDFILL91_1293 VDD VSS sg13g2_FILL8
XSTDFILL91_1301 VDD VSS sg13g2_FILL8
XSTDFILL91_1309 VDD VSS sg13g2_FILL8
XSTDFILL91_1317 VDD VSS sg13g2_FILL8
XSTDFILL91_1325 VDD VSS sg13g2_FILL8
XSTDFILL91_1333 VDD VSS sg13g2_FILL8
XSTDFILL91_1341 VDD VSS sg13g2_FILL8
XSTDFILL91_1349 VDD VSS sg13g2_FILL8
XSTDFILL91_1357 VDD VSS sg13g2_FILL8
XSTDFILL91_1365 VDD VSS sg13g2_FILL8
XSTDFILL91_1373 VDD VSS sg13g2_FILL8
XSTDFILL91_1381 VDD VSS sg13g2_FILL8
XSTDFILL91_1389 VDD VSS sg13g2_FILL8
XSTDFILL91_1397 VDD VSS sg13g2_FILL8
XSTDFILL91_1405 VDD VSS sg13g2_FILL8
XSTDFILL91_1413 VDD VSS sg13g2_FILL8
XSTDFILL91_1421 VDD VSS sg13g2_FILL8
XSTDFILL91_1429 VDD VSS sg13g2_FILL8
XSTDFILL91_1437 VDD VSS sg13g2_FILL8
XSTDFILL91_1445 VDD VSS sg13g2_FILL8
XSTDFILL91_1453 VDD VSS sg13g2_FILL8
XSTDFILL91_1461 VDD VSS sg13g2_FILL8
XSTDFILL91_1469 VDD VSS sg13g2_FILL8
XSTDFILL91_1477 VDD VSS sg13g2_FILL8
XSTDFILL91_1485 VDD VSS sg13g2_FILL8
XSTDFILL91_1493 VDD VSS sg13g2_FILL8
XSTDFILL91_1501 VDD VSS sg13g2_FILL8
XSTDFILL91_1509 VDD VSS sg13g2_FILL8
XSTDFILL91_1517 VDD VSS sg13g2_FILL8
XSTDFILL92_0 VDD VSS sg13g2_FILL8
XSTDFILL92_8 VDD VSS sg13g2_FILL8
XSTDFILL92_16 VDD VSS sg13g2_FILL8
XSTDFILL92_24 VDD VSS sg13g2_FILL8
XSTDFILL92_32 VDD VSS sg13g2_FILL8
XSTDFILL92_40 VDD VSS sg13g2_FILL8
XSTDFILL92_48 VDD VSS sg13g2_FILL8
XSTDFILL92_56 VDD VSS sg13g2_FILL8
XSTDFILL92_64 VDD VSS sg13g2_FILL8
XSTDFILL92_72 VDD VSS sg13g2_FILL8
XSTDFILL92_80 VDD VSS sg13g2_FILL8
XSTDFILL92_88 VDD VSS sg13g2_FILL8
XSTDFILL92_96 VDD VSS sg13g2_FILL8
XSTDFILL92_104 VDD VSS sg13g2_FILL8
XSTDFILL92_112 VDD VSS sg13g2_FILL8
XSTDFILL92_120 VDD VSS sg13g2_FILL8
XSTDFILL92_128 VDD VSS sg13g2_FILL4
XSTDFILL92_1085 VDD VSS sg13g2_FILL8
XSTDFILL92_1093 VDD VSS sg13g2_FILL8
XSTDFILL92_1101 VDD VSS sg13g2_FILL8
XSTDFILL92_1109 VDD VSS sg13g2_FILL8
XSTDFILL92_1117 VDD VSS sg13g2_FILL8
XSTDFILL92_1125 VDD VSS sg13g2_FILL8
XSTDFILL92_1133 VDD VSS sg13g2_FILL8
XSTDFILL92_1141 VDD VSS sg13g2_FILL8
XSTDFILL92_1149 VDD VSS sg13g2_FILL8
XSTDFILL92_1157 VDD VSS sg13g2_FILL8
XSTDFILL92_1165 VDD VSS sg13g2_FILL8
XSTDFILL92_1173 VDD VSS sg13g2_FILL8
XSTDFILL92_1181 VDD VSS sg13g2_FILL8
XSTDFILL92_1189 VDD VSS sg13g2_FILL8
XSTDFILL92_1197 VDD VSS sg13g2_FILL8
XSTDFILL92_1205 VDD VSS sg13g2_FILL8
XSTDFILL92_1213 VDD VSS sg13g2_FILL8
XSTDFILL92_1221 VDD VSS sg13g2_FILL8
XSTDFILL92_1229 VDD VSS sg13g2_FILL8
XSTDFILL92_1237 VDD VSS sg13g2_FILL8
XSTDFILL92_1245 VDD VSS sg13g2_FILL8
XSTDFILL92_1253 VDD VSS sg13g2_FILL8
XSTDFILL92_1261 VDD VSS sg13g2_FILL8
XSTDFILL92_1269 VDD VSS sg13g2_FILL8
XSTDFILL92_1277 VDD VSS sg13g2_FILL8
XSTDFILL92_1285 VDD VSS sg13g2_FILL8
XSTDFILL92_1293 VDD VSS sg13g2_FILL8
XSTDFILL92_1301 VDD VSS sg13g2_FILL8
XSTDFILL92_1309 VDD VSS sg13g2_FILL8
XSTDFILL92_1317 VDD VSS sg13g2_FILL8
XSTDFILL92_1325 VDD VSS sg13g2_FILL8
XSTDFILL92_1333 VDD VSS sg13g2_FILL8
XSTDFILL92_1341 VDD VSS sg13g2_FILL8
XSTDFILL92_1349 VDD VSS sg13g2_FILL8
XSTDFILL92_1357 VDD VSS sg13g2_FILL8
XSTDFILL92_1365 VDD VSS sg13g2_FILL8
XSTDFILL92_1373 VDD VSS sg13g2_FILL8
XSTDFILL92_1381 VDD VSS sg13g2_FILL8
XSTDFILL92_1389 VDD VSS sg13g2_FILL8
XSTDFILL92_1397 VDD VSS sg13g2_FILL8
XSTDFILL92_1405 VDD VSS sg13g2_FILL8
XSTDFILL92_1413 VDD VSS sg13g2_FILL8
XSTDFILL92_1421 VDD VSS sg13g2_FILL8
XSTDFILL92_1429 VDD VSS sg13g2_FILL8
XSTDFILL92_1437 VDD VSS sg13g2_FILL8
XSTDFILL92_1445 VDD VSS sg13g2_FILL8
XSTDFILL92_1453 VDD VSS sg13g2_FILL8
XSTDFILL92_1461 VDD VSS sg13g2_FILL8
XSTDFILL92_1469 VDD VSS sg13g2_FILL8
XSTDFILL92_1477 VDD VSS sg13g2_FILL8
XSTDFILL92_1485 VDD VSS sg13g2_FILL8
XSTDFILL92_1493 VDD VSS sg13g2_FILL8
XSTDFILL92_1501 VDD VSS sg13g2_FILL8
XSTDFILL92_1509 VDD VSS sg13g2_FILL8
XSTDFILL92_1517 VDD VSS sg13g2_FILL8
XSTDFILL93_0 VDD VSS sg13g2_FILL8
XSTDFILL93_8 VDD VSS sg13g2_FILL8
XSTDFILL93_16 VDD VSS sg13g2_FILL8
XSTDFILL93_24 VDD VSS sg13g2_FILL8
XSTDFILL93_32 VDD VSS sg13g2_FILL8
XSTDFILL93_40 VDD VSS sg13g2_FILL8
XSTDFILL93_48 VDD VSS sg13g2_FILL8
XSTDFILL93_56 VDD VSS sg13g2_FILL8
XSTDFILL93_64 VDD VSS sg13g2_FILL8
XSTDFILL93_72 VDD VSS sg13g2_FILL8
XSTDFILL93_80 VDD VSS sg13g2_FILL8
XSTDFILL93_88 VDD VSS sg13g2_FILL8
XSTDFILL93_96 VDD VSS sg13g2_FILL8
XSTDFILL93_104 VDD VSS sg13g2_FILL8
XSTDFILL93_112 VDD VSS sg13g2_FILL8
XSTDFILL93_120 VDD VSS sg13g2_FILL8
XSTDFILL93_128 VDD VSS sg13g2_FILL8
XSTDFILL93_136 VDD VSS sg13g2_FILL8
XSTDFILL93_144 VDD VSS sg13g2_FILL8
XSTDFILL93_152 VDD VSS sg13g2_FILL8
XSTDFILL93_160 VDD VSS sg13g2_FILL8
XSTDFILL93_168 VDD VSS sg13g2_FILL8
XSTDFILL93_176 VDD VSS sg13g2_FILL8
XSTDFILL93_184 VDD VSS sg13g2_FILL8
XSTDFILL93_192 VDD VSS sg13g2_FILL8
XSTDFILL93_200 VDD VSS sg13g2_FILL8
XSTDFILL93_208 VDD VSS sg13g2_FILL8
XSTDFILL93_216 VDD VSS sg13g2_FILL8
XSTDFILL93_224 VDD VSS sg13g2_FILL8
XSTDFILL93_232 VDD VSS sg13g2_FILL8
XSTDFILL93_240 VDD VSS sg13g2_FILL8
XSTDFILL93_248 VDD VSS sg13g2_FILL8
XSTDFILL93_256 VDD VSS sg13g2_FILL8
XSTDFILL93_264 VDD VSS sg13g2_FILL8
XSTDFILL93_272 VDD VSS sg13g2_FILL8
XSTDFILL93_280 VDD VSS sg13g2_FILL8
XSTDFILL93_288 VDD VSS sg13g2_FILL8
XSTDFILL93_296 VDD VSS sg13g2_FILL8
XSTDFILL93_304 VDD VSS sg13g2_FILL8
XSTDFILL93_312 VDD VSS sg13g2_FILL8
XSTDFILL93_320 VDD VSS sg13g2_FILL8
XSTDFILL93_328 VDD VSS sg13g2_FILL8
XSTDFILL93_336 VDD VSS sg13g2_FILL8
XSTDFILL93_344 VDD VSS sg13g2_FILL8
XSTDFILL93_352 VDD VSS sg13g2_FILL8
XSTDFILL93_360 VDD VSS sg13g2_FILL8
XSTDFILL93_368 VDD VSS sg13g2_FILL8
XSTDFILL93_376 VDD VSS sg13g2_FILL8
XSTDFILL93_384 VDD VSS sg13g2_FILL8
XSTDFILL93_392 VDD VSS sg13g2_FILL8
XSTDFILL93_400 VDD VSS sg13g2_FILL8
XSTDFILL93_408 VDD VSS sg13g2_FILL8
XSTDFILL93_416 VDD VSS sg13g2_FILL8
XSTDFILL93_424 VDD VSS sg13g2_FILL8
XSTDFILL93_432 VDD VSS sg13g2_FILL8
XSTDFILL93_440 VDD VSS sg13g2_FILL8
XSTDFILL93_448 VDD VSS sg13g2_FILL8
XSTDFILL93_456 VDD VSS sg13g2_FILL8
XSTDFILL93_464 VDD VSS sg13g2_FILL8
XSTDFILL93_472 VDD VSS sg13g2_FILL8
XSTDFILL93_480 VDD VSS sg13g2_FILL1
XSTDFILL93_489 VDD VSS sg13g2_FILL4
XSTDFILL93_493 VDD VSS sg13g2_FILL1
XSTDFILL93_507 VDD VSS sg13g2_FILL2
XSTDFILL93_509 VDD VSS sg13g2_FILL1
XSTDFILL93_518 VDD VSS sg13g2_FILL4
XSTDFILL93_537 VDD VSS sg13g2_FILL8
XSTDFILL93_545 VDD VSS sg13g2_FILL8
XSTDFILL93_553 VDD VSS sg13g2_FILL2
XSTDFILL93_555 VDD VSS sg13g2_FILL1
XSTDFILL93_566 VDD VSS sg13g2_FILL1
XSTDFILL93_580 VDD VSS sg13g2_FILL4
XSTDFILL93_612 VDD VSS sg13g2_FILL1
XSTDFILL93_636 VDD VSS sg13g2_FILL2
XSTDFILL93_638 VDD VSS sg13g2_FILL1
XSTDFILL93_647 VDD VSS sg13g2_FILL2
XSTDFILL93_649 VDD VSS sg13g2_FILL1
XSTDFILL93_663 VDD VSS sg13g2_FILL2
XSTDFILL93_665 VDD VSS sg13g2_FILL1
XSTDFILL93_686 VDD VSS sg13g2_FILL2
XSTDFILL93_688 VDD VSS sg13g2_FILL1
XSTDFILL93_715 VDD VSS sg13g2_FILL2
XSTDFILL93_730 VDD VSS sg13g2_FILL8
XSTDFILL93_738 VDD VSS sg13g2_FILL1
XSTDFILL93_747 VDD VSS sg13g2_FILL8
XSTDFILL93_755 VDD VSS sg13g2_FILL2
XSTDFILL93_765 VDD VSS sg13g2_FILL8
XSTDFILL93_773 VDD VSS sg13g2_FILL8
XSTDFILL93_781 VDD VSS sg13g2_FILL8
XSTDFILL93_789 VDD VSS sg13g2_FILL8
XSTDFILL93_805 VDD VSS sg13g2_FILL8
XSTDFILL93_813 VDD VSS sg13g2_FILL8
XSTDFILL93_821 VDD VSS sg13g2_FILL8
XSTDFILL93_829 VDD VSS sg13g2_FILL1
XSTDFILL93_838 VDD VSS sg13g2_FILL8
XSTDFILL93_846 VDD VSS sg13g2_FILL2
XSTDFILL93_856 VDD VSS sg13g2_FILL4
XSTDFILL93_860 VDD VSS sg13g2_FILL1
XSTDFILL93_869 VDD VSS sg13g2_FILL2
XSTDFILL93_879 VDD VSS sg13g2_FILL8
XSTDFILL93_887 VDD VSS sg13g2_FILL4
XSTDFILL93_891 VDD VSS sg13g2_FILL2
XSTDFILL93_901 VDD VSS sg13g2_FILL8
XSTDFILL93_909 VDD VSS sg13g2_FILL8
XSTDFILL93_917 VDD VSS sg13g2_FILL8
XSTDFILL93_925 VDD VSS sg13g2_FILL2
XSTDFILL93_935 VDD VSS sg13g2_FILL8
XSTDFILL93_943 VDD VSS sg13g2_FILL8
XSTDFILL93_951 VDD VSS sg13g2_FILL4
XSTDFILL93_955 VDD VSS sg13g2_FILL1
XSTDFILL93_964 VDD VSS sg13g2_FILL8
XSTDFILL93_972 VDD VSS sg13g2_FILL8
XSTDFILL93_980 VDD VSS sg13g2_FILL8
XSTDFILL93_988 VDD VSS sg13g2_FILL8
XSTDFILL93_996 VDD VSS sg13g2_FILL8
XSTDFILL93_1004 VDD VSS sg13g2_FILL8
XSTDFILL93_1012 VDD VSS sg13g2_FILL8
XSTDFILL93_1020 VDD VSS sg13g2_FILL8
XSTDFILL93_1028 VDD VSS sg13g2_FILL8
XSTDFILL93_1036 VDD VSS sg13g2_FILL8
XSTDFILL93_1044 VDD VSS sg13g2_FILL8
XSTDFILL93_1052 VDD VSS sg13g2_FILL8
XSTDFILL93_1060 VDD VSS sg13g2_FILL8
XSTDFILL93_1068 VDD VSS sg13g2_FILL8
XSTDFILL93_1076 VDD VSS sg13g2_FILL8
XSTDFILL93_1084 VDD VSS sg13g2_FILL8
XSTDFILL93_1092 VDD VSS sg13g2_FILL8
XSTDFILL93_1100 VDD VSS sg13g2_FILL8
XSTDFILL93_1108 VDD VSS sg13g2_FILL8
XSTDFILL93_1116 VDD VSS sg13g2_FILL8
XSTDFILL93_1124 VDD VSS sg13g2_FILL8
XSTDFILL93_1132 VDD VSS sg13g2_FILL8
XSTDFILL93_1140 VDD VSS sg13g2_FILL8
XSTDFILL93_1148 VDD VSS sg13g2_FILL8
XSTDFILL93_1156 VDD VSS sg13g2_FILL8
XSTDFILL93_1164 VDD VSS sg13g2_FILL8
XSTDFILL93_1172 VDD VSS sg13g2_FILL8
XSTDFILL93_1180 VDD VSS sg13g2_FILL8
XSTDFILL93_1188 VDD VSS sg13g2_FILL8
XSTDFILL93_1196 VDD VSS sg13g2_FILL8
XSTDFILL93_1204 VDD VSS sg13g2_FILL8
XSTDFILL93_1212 VDD VSS sg13g2_FILL8
XSTDFILL93_1220 VDD VSS sg13g2_FILL8
XSTDFILL93_1228 VDD VSS sg13g2_FILL8
XSTDFILL93_1236 VDD VSS sg13g2_FILL8
XSTDFILL93_1244 VDD VSS sg13g2_FILL8
XSTDFILL93_1252 VDD VSS sg13g2_FILL8
XSTDFILL93_1260 VDD VSS sg13g2_FILL8
XSTDFILL93_1268 VDD VSS sg13g2_FILL8
XSTDFILL93_1276 VDD VSS sg13g2_FILL8
XSTDFILL93_1284 VDD VSS sg13g2_FILL8
XSTDFILL93_1292 VDD VSS sg13g2_FILL8
XSTDFILL93_1300 VDD VSS sg13g2_FILL8
XSTDFILL93_1308 VDD VSS sg13g2_FILL8
XSTDFILL93_1316 VDD VSS sg13g2_FILL8
XSTDFILL93_1324 VDD VSS sg13g2_FILL8
XSTDFILL93_1332 VDD VSS sg13g2_FILL8
XSTDFILL93_1340 VDD VSS sg13g2_FILL8
XSTDFILL93_1348 VDD VSS sg13g2_FILL8
XSTDFILL93_1356 VDD VSS sg13g2_FILL8
XSTDFILL93_1364 VDD VSS sg13g2_FILL8
XSTDFILL93_1372 VDD VSS sg13g2_FILL8
XSTDFILL93_1380 VDD VSS sg13g2_FILL8
XSTDFILL93_1388 VDD VSS sg13g2_FILL8
XSTDFILL93_1396 VDD VSS sg13g2_FILL8
XSTDFILL93_1404 VDD VSS sg13g2_FILL8
XSTDFILL93_1412 VDD VSS sg13g2_FILL8
XSTDFILL93_1420 VDD VSS sg13g2_FILL8
XSTDFILL93_1428 VDD VSS sg13g2_FILL8
XSTDFILL93_1436 VDD VSS sg13g2_FILL8
XSTDFILL93_1444 VDD VSS sg13g2_FILL8
XSTDFILL93_1452 VDD VSS sg13g2_FILL8
XSTDFILL93_1460 VDD VSS sg13g2_FILL8
XSTDFILL93_1468 VDD VSS sg13g2_FILL8
XSTDFILL93_1476 VDD VSS sg13g2_FILL8
XSTDFILL93_1484 VDD VSS sg13g2_FILL8
XSTDFILL93_1492 VDD VSS sg13g2_FILL8
XSTDFILL93_1500 VDD VSS sg13g2_FILL8
XSTDFILL93_1508 VDD VSS sg13g2_FILL8
XSTDFILL93_1516 VDD VSS sg13g2_FILL8
XSTDFILL93_1524 VDD VSS sg13g2_FILL8
XSTDFILL93_1532 VDD VSS sg13g2_FILL8
XSTDFILL93_1540 VDD VSS sg13g2_FILL8
XSTDFILL93_1548 VDD VSS sg13g2_FILL8
XSTDFILL93_1556 VDD VSS sg13g2_FILL8
XSTDFILL93_1564 VDD VSS sg13g2_FILL8
XSTDFILL93_1572 VDD VSS sg13g2_FILL8
XSTDFILL93_1580 VDD VSS sg13g2_FILL8
XSTDFILL93_1588 VDD VSS sg13g2_FILL8
XSTDFILL93_1596 VDD VSS sg13g2_FILL8
XSTDFILL93_1604 VDD VSS sg13g2_FILL8
XSTDFILL93_1612 VDD VSS sg13g2_FILL8
XSTDFILL93_1620 VDD VSS sg13g2_FILL8
XSTDFILL93_1628 VDD VSS sg13g2_FILL8
XSTDFILL93_1636 VDD VSS sg13g2_FILL8
XSTDFILL93_1644 VDD VSS sg13g2_FILL8
XSTDFILL93_1652 VDD VSS sg13g2_FILL8
XSTDFILL93_1660 VDD VSS sg13g2_FILL8
XSTDFILL93_1668 VDD VSS sg13g2_FILL8
XSTDFILL93_1676 VDD VSS sg13g2_FILL8
XSTDFILL93_1684 VDD VSS sg13g2_FILL8
XSTDFILL93_1692 VDD VSS sg13g2_FILL8
XSTDFILL93_1700 VDD VSS sg13g2_FILL8
XSTDFILL93_1708 VDD VSS sg13g2_FILL8
XSTDFILL93_1716 VDD VSS sg13g2_FILL8
XSTDFILL93_1724 VDD VSS sg13g2_FILL8
XSTDFILL93_1732 VDD VSS sg13g2_FILL8
XSTDFILL93_1740 VDD VSS sg13g2_FILL8
XSTDFILL93_1748 VDD VSS sg13g2_FILL8
XSTDFILL93_1756 VDD VSS sg13g2_FILL8
XSTDFILL93_1764 VDD VSS sg13g2_FILL8
XSTDFILL93_1772 VDD VSS sg13g2_FILL8
XSTDFILL93_1780 VDD VSS sg13g2_FILL8
XSTDFILL93_1788 VDD VSS sg13g2_FILL8
XSTDFILL93_1796 VDD VSS sg13g2_FILL8
XSTDFILL93_1804 VDD VSS sg13g2_FILL8
XSTDFILL93_1812 VDD VSS sg13g2_FILL8
XSTDFILL93_1820 VDD VSS sg13g2_FILL8
XSTDFILL93_1828 VDD VSS sg13g2_FILL8
XSTDFILL93_1836 VDD VSS sg13g2_FILL8
XSTDFILL93_1844 VDD VSS sg13g2_FILL8
XSTDFILL93_1852 VDD VSS sg13g2_FILL8
XSTDFILL93_1860 VDD VSS sg13g2_FILL8
XSTDFILL93_1868 VDD VSS sg13g2_FILL8
XSTDFILL93_1876 VDD VSS sg13g2_FILL8
XSTDFILL93_1884 VDD VSS sg13g2_FILL8
XSTDFILL93_1892 VDD VSS sg13g2_FILL8
XSTDFILL93_1900 VDD VSS sg13g2_FILL8
XSTDFILL93_1908 VDD VSS sg13g2_FILL8
XSTDFILL93_1916 VDD VSS sg13g2_FILL8
XSTDFILL93_1924 VDD VSS sg13g2_FILL8
XSTDFILL93_1932 VDD VSS sg13g2_FILL8
XSTDFILL93_1940 VDD VSS sg13g2_FILL8
XSTDFILL93_1948 VDD VSS sg13g2_FILL8
XSTDFILL93_1956 VDD VSS sg13g2_FILL8
XSTDFILL93_1964 VDD VSS sg13g2_FILL8
XSTDFILL93_1972 VDD VSS sg13g2_FILL8
XSTDFILL93_1980 VDD VSS sg13g2_FILL8
XSTDFILL93_1988 VDD VSS sg13g2_FILL8
XSTDFILL93_1996 VDD VSS sg13g2_FILL8
XSTDFILL93_2004 VDD VSS sg13g2_FILL8
XSTDFILL93_2012 VDD VSS sg13g2_FILL8
XSTDFILL93_2020 VDD VSS sg13g2_FILL8
XSTDFILL93_2028 VDD VSS sg13g2_FILL8
XSTDFILL93_2036 VDD VSS sg13g2_FILL8
XSTDFILL93_2044 VDD VSS sg13g2_FILL8
XSTDFILL93_2052 VDD VSS sg13g2_FILL8
XSTDFILL93_2060 VDD VSS sg13g2_FILL8
XSTDFILL93_2068 VDD VSS sg13g2_FILL8
XSTDFILL93_2076 VDD VSS sg13g2_FILL8
XSTDFILL93_2084 VDD VSS sg13g2_FILL8
XSTDFILL93_2092 VDD VSS sg13g2_FILL8
XSTDFILL93_2100 VDD VSS sg13g2_FILL8
XSTDFILL93_2108 VDD VSS sg13g2_FILL8
XSTDFILL93_2116 VDD VSS sg13g2_FILL8
XSTDFILL93_2124 VDD VSS sg13g2_FILL8
XSTDFILL93_2132 VDD VSS sg13g2_FILL8
XSTDFILL93_2140 VDD VSS sg13g2_FILL8
XSTDFILL93_2148 VDD VSS sg13g2_FILL4
XSTDFILL93_2152 VDD VSS sg13g2_FILL2
XSTDFILL94_0 VDD VSS sg13g2_FILL8
XSTDFILL94_8 VDD VSS sg13g2_FILL8
XSTDFILL94_16 VDD VSS sg13g2_FILL8
XSTDFILL94_24 VDD VSS sg13g2_FILL8
XSTDFILL94_32 VDD VSS sg13g2_FILL8
XSTDFILL94_40 VDD VSS sg13g2_FILL8
XSTDFILL94_48 VDD VSS sg13g2_FILL8
XSTDFILL94_56 VDD VSS sg13g2_FILL8
XSTDFILL94_64 VDD VSS sg13g2_FILL8
XSTDFILL94_72 VDD VSS sg13g2_FILL8
XSTDFILL94_80 VDD VSS sg13g2_FILL8
XSTDFILL94_88 VDD VSS sg13g2_FILL8
XSTDFILL94_96 VDD VSS sg13g2_FILL8
XSTDFILL94_104 VDD VSS sg13g2_FILL8
XSTDFILL94_112 VDD VSS sg13g2_FILL8
XSTDFILL94_120 VDD VSS sg13g2_FILL8
XSTDFILL94_128 VDD VSS sg13g2_FILL8
XSTDFILL94_136 VDD VSS sg13g2_FILL8
XSTDFILL94_144 VDD VSS sg13g2_FILL8
XSTDFILL94_152 VDD VSS sg13g2_FILL8
XSTDFILL94_160 VDD VSS sg13g2_FILL8
XSTDFILL94_168 VDD VSS sg13g2_FILL8
XSTDFILL94_176 VDD VSS sg13g2_FILL8
XSTDFILL94_184 VDD VSS sg13g2_FILL8
XSTDFILL94_192 VDD VSS sg13g2_FILL8
XSTDFILL94_200 VDD VSS sg13g2_FILL8
XSTDFILL94_208 VDD VSS sg13g2_FILL8
XSTDFILL94_216 VDD VSS sg13g2_FILL8
XSTDFILL94_224 VDD VSS sg13g2_FILL8
XSTDFILL94_232 VDD VSS sg13g2_FILL8
XSTDFILL94_240 VDD VSS sg13g2_FILL8
XSTDFILL94_248 VDD VSS sg13g2_FILL8
XSTDFILL94_256 VDD VSS sg13g2_FILL8
XSTDFILL94_264 VDD VSS sg13g2_FILL8
XSTDFILL94_272 VDD VSS sg13g2_FILL8
XSTDFILL94_280 VDD VSS sg13g2_FILL8
XSTDFILL94_288 VDD VSS sg13g2_FILL8
XSTDFILL94_296 VDD VSS sg13g2_FILL8
XSTDFILL94_304 VDD VSS sg13g2_FILL8
XSTDFILL94_312 VDD VSS sg13g2_FILL8
XSTDFILL94_320 VDD VSS sg13g2_FILL8
XSTDFILL94_328 VDD VSS sg13g2_FILL8
XSTDFILL94_336 VDD VSS sg13g2_FILL8
XSTDFILL94_344 VDD VSS sg13g2_FILL8
XSTDFILL94_352 VDD VSS sg13g2_FILL8
XSTDFILL94_360 VDD VSS sg13g2_FILL8
XSTDFILL94_368 VDD VSS sg13g2_FILL8
XSTDFILL94_376 VDD VSS sg13g2_FILL8
XSTDFILL94_384 VDD VSS sg13g2_FILL8
XSTDFILL94_392 VDD VSS sg13g2_FILL8
XSTDFILL94_400 VDD VSS sg13g2_FILL8
XSTDFILL94_408 VDD VSS sg13g2_FILL8
XSTDFILL94_416 VDD VSS sg13g2_FILL8
XSTDFILL94_424 VDD VSS sg13g2_FILL8
XSTDFILL94_432 VDD VSS sg13g2_FILL8
XSTDFILL94_440 VDD VSS sg13g2_FILL8
XSTDFILL94_448 VDD VSS sg13g2_FILL8
XSTDFILL94_456 VDD VSS sg13g2_FILL8
XSTDFILL94_464 VDD VSS sg13g2_FILL8
XSTDFILL94_472 VDD VSS sg13g2_FILL8
XSTDFILL94_480 VDD VSS sg13g2_FILL8
XSTDFILL94_488 VDD VSS sg13g2_FILL8
XSTDFILL94_496 VDD VSS sg13g2_FILL8
XSTDFILL94_504 VDD VSS sg13g2_FILL8
XSTDFILL94_512 VDD VSS sg13g2_FILL8
XSTDFILL94_520 VDD VSS sg13g2_FILL8
XSTDFILL94_528 VDD VSS sg13g2_FILL8
XSTDFILL94_536 VDD VSS sg13g2_FILL8
XSTDFILL94_544 VDD VSS sg13g2_FILL8
XSTDFILL94_552 VDD VSS sg13g2_FILL8
XSTDFILL94_560 VDD VSS sg13g2_FILL8
XSTDFILL94_568 VDD VSS sg13g2_FILL8
XSTDFILL94_576 VDD VSS sg13g2_FILL8
XSTDFILL94_584 VDD VSS sg13g2_FILL2
XSTDFILL94_586 VDD VSS sg13g2_FILL1
XSTDFILL94_592 VDD VSS sg13g2_FILL8
XSTDFILL94_600 VDD VSS sg13g2_FILL8
XSTDFILL94_608 VDD VSS sg13g2_FILL8
XSTDFILL94_616 VDD VSS sg13g2_FILL1
XSTDFILL94_622 VDD VSS sg13g2_FILL8
XSTDFILL94_630 VDD VSS sg13g2_FILL8
XSTDFILL94_638 VDD VSS sg13g2_FILL8
XSTDFILL94_646 VDD VSS sg13g2_FILL4
XSTDFILL94_650 VDD VSS sg13g2_FILL1
XSTDFILL94_656 VDD VSS sg13g2_FILL8
XSTDFILL94_664 VDD VSS sg13g2_FILL8
XSTDFILL94_672 VDD VSS sg13g2_FILL8
XSTDFILL94_680 VDD VSS sg13g2_FILL8
XSTDFILL94_688 VDD VSS sg13g2_FILL8
XSTDFILL94_696 VDD VSS sg13g2_FILL8
XSTDFILL94_704 VDD VSS sg13g2_FILL8
XSTDFILL94_712 VDD VSS sg13g2_FILL8
XSTDFILL94_720 VDD VSS sg13g2_FILL8
XSTDFILL94_728 VDD VSS sg13g2_FILL8
XSTDFILL94_736 VDD VSS sg13g2_FILL8
XSTDFILL94_744 VDD VSS sg13g2_FILL8
XSTDFILL94_752 VDD VSS sg13g2_FILL8
XSTDFILL94_760 VDD VSS sg13g2_FILL8
XSTDFILL94_768 VDD VSS sg13g2_FILL8
XSTDFILL94_776 VDD VSS sg13g2_FILL8
XSTDFILL94_784 VDD VSS sg13g2_FILL8
XSTDFILL94_792 VDD VSS sg13g2_FILL8
XSTDFILL94_800 VDD VSS sg13g2_FILL8
XSTDFILL94_808 VDD VSS sg13g2_FILL8
XSTDFILL94_816 VDD VSS sg13g2_FILL8
XSTDFILL94_824 VDD VSS sg13g2_FILL8
XSTDFILL94_832 VDD VSS sg13g2_FILL8
XSTDFILL94_840 VDD VSS sg13g2_FILL8
XSTDFILL94_848 VDD VSS sg13g2_FILL8
XSTDFILL94_856 VDD VSS sg13g2_FILL8
XSTDFILL94_864 VDD VSS sg13g2_FILL8
XSTDFILL94_872 VDD VSS sg13g2_FILL8
XSTDFILL94_880 VDD VSS sg13g2_FILL8
XSTDFILL94_888 VDD VSS sg13g2_FILL8
XSTDFILL94_896 VDD VSS sg13g2_FILL8
XSTDFILL94_904 VDD VSS sg13g2_FILL8
XSTDFILL94_912 VDD VSS sg13g2_FILL8
XSTDFILL94_920 VDD VSS sg13g2_FILL8
XSTDFILL94_928 VDD VSS sg13g2_FILL8
XSTDFILL94_936 VDD VSS sg13g2_FILL8
XSTDFILL94_944 VDD VSS sg13g2_FILL8
XSTDFILL94_952 VDD VSS sg13g2_FILL8
XSTDFILL94_960 VDD VSS sg13g2_FILL8
XSTDFILL94_968 VDD VSS sg13g2_FILL8
XSTDFILL94_976 VDD VSS sg13g2_FILL8
XSTDFILL94_984 VDD VSS sg13g2_FILL8
XSTDFILL94_992 VDD VSS sg13g2_FILL8
XSTDFILL94_1000 VDD VSS sg13g2_FILL8
XSTDFILL94_1008 VDD VSS sg13g2_FILL8
XSTDFILL94_1016 VDD VSS sg13g2_FILL8
XSTDFILL94_1024 VDD VSS sg13g2_FILL8
XSTDFILL94_1032 VDD VSS sg13g2_FILL8
XSTDFILL94_1040 VDD VSS sg13g2_FILL8
XSTDFILL94_1048 VDD VSS sg13g2_FILL8
XSTDFILL94_1056 VDD VSS sg13g2_FILL8
XSTDFILL94_1064 VDD VSS sg13g2_FILL8
XSTDFILL94_1072 VDD VSS sg13g2_FILL8
XSTDFILL94_1080 VDD VSS sg13g2_FILL8
XSTDFILL94_1088 VDD VSS sg13g2_FILL8
XSTDFILL94_1096 VDD VSS sg13g2_FILL8
XSTDFILL94_1104 VDD VSS sg13g2_FILL8
XSTDFILL94_1112 VDD VSS sg13g2_FILL8
XSTDFILL94_1120 VDD VSS sg13g2_FILL8
XSTDFILL94_1128 VDD VSS sg13g2_FILL8
XSTDFILL94_1136 VDD VSS sg13g2_FILL8
XSTDFILL94_1144 VDD VSS sg13g2_FILL8
XSTDFILL94_1152 VDD VSS sg13g2_FILL8
XSTDFILL94_1160 VDD VSS sg13g2_FILL8
XSTDFILL94_1168 VDD VSS sg13g2_FILL8
XSTDFILL94_1176 VDD VSS sg13g2_FILL8
XSTDFILL94_1184 VDD VSS sg13g2_FILL8
XSTDFILL94_1192 VDD VSS sg13g2_FILL8
XSTDFILL94_1200 VDD VSS sg13g2_FILL8
XSTDFILL94_1208 VDD VSS sg13g2_FILL8
XSTDFILL94_1216 VDD VSS sg13g2_FILL8
XSTDFILL94_1224 VDD VSS sg13g2_FILL8
XSTDFILL94_1232 VDD VSS sg13g2_FILL8
XSTDFILL94_1240 VDD VSS sg13g2_FILL8
XSTDFILL94_1248 VDD VSS sg13g2_FILL8
XSTDFILL94_1256 VDD VSS sg13g2_FILL8
XSTDFILL94_1264 VDD VSS sg13g2_FILL8
XSTDFILL94_1272 VDD VSS sg13g2_FILL8
XSTDFILL94_1280 VDD VSS sg13g2_FILL8
XSTDFILL94_1288 VDD VSS sg13g2_FILL8
XSTDFILL94_1296 VDD VSS sg13g2_FILL8
XSTDFILL94_1304 VDD VSS sg13g2_FILL8
XSTDFILL94_1312 VDD VSS sg13g2_FILL8
XSTDFILL94_1320 VDD VSS sg13g2_FILL8
XSTDFILL94_1328 VDD VSS sg13g2_FILL8
XSTDFILL94_1336 VDD VSS sg13g2_FILL8
XSTDFILL94_1344 VDD VSS sg13g2_FILL8
XSTDFILL94_1352 VDD VSS sg13g2_FILL8
XSTDFILL94_1360 VDD VSS sg13g2_FILL8
XSTDFILL94_1368 VDD VSS sg13g2_FILL8
XSTDFILL94_1376 VDD VSS sg13g2_FILL8
XSTDFILL94_1384 VDD VSS sg13g2_FILL8
XSTDFILL94_1392 VDD VSS sg13g2_FILL8
XSTDFILL94_1400 VDD VSS sg13g2_FILL8
XSTDFILL94_1408 VDD VSS sg13g2_FILL8
XSTDFILL94_1416 VDD VSS sg13g2_FILL8
XSTDFILL94_1424 VDD VSS sg13g2_FILL8
XSTDFILL94_1432 VDD VSS sg13g2_FILL8
XSTDFILL94_1440 VDD VSS sg13g2_FILL8
XSTDFILL94_1448 VDD VSS sg13g2_FILL8
XSTDFILL94_1456 VDD VSS sg13g2_FILL8
XSTDFILL94_1464 VDD VSS sg13g2_FILL8
XSTDFILL94_1472 VDD VSS sg13g2_FILL8
XSTDFILL94_1480 VDD VSS sg13g2_FILL8
XSTDFILL94_1488 VDD VSS sg13g2_FILL8
XSTDFILL94_1496 VDD VSS sg13g2_FILL8
XSTDFILL94_1504 VDD VSS sg13g2_FILL8
XSTDFILL94_1512 VDD VSS sg13g2_FILL8
XSTDFILL94_1520 VDD VSS sg13g2_FILL8
XSTDFILL94_1528 VDD VSS sg13g2_FILL8
XSTDFILL94_1536 VDD VSS sg13g2_FILL8
XSTDFILL94_1544 VDD VSS sg13g2_FILL8
XSTDFILL94_1552 VDD VSS sg13g2_FILL8
XSTDFILL94_1560 VDD VSS sg13g2_FILL8
XSTDFILL94_1568 VDD VSS sg13g2_FILL8
XSTDFILL94_1576 VDD VSS sg13g2_FILL8
XSTDFILL94_1584 VDD VSS sg13g2_FILL8
XSTDFILL94_1592 VDD VSS sg13g2_FILL8
XSTDFILL94_1600 VDD VSS sg13g2_FILL8
XSTDFILL94_1608 VDD VSS sg13g2_FILL8
XSTDFILL94_1616 VDD VSS sg13g2_FILL8
XSTDFILL94_1624 VDD VSS sg13g2_FILL8
XSTDFILL94_1632 VDD VSS sg13g2_FILL8
XSTDFILL94_1640 VDD VSS sg13g2_FILL8
XSTDFILL94_1648 VDD VSS sg13g2_FILL8
XSTDFILL94_1656 VDD VSS sg13g2_FILL8
XSTDFILL94_1664 VDD VSS sg13g2_FILL8
XSTDFILL94_1672 VDD VSS sg13g2_FILL8
XSTDFILL94_1680 VDD VSS sg13g2_FILL8
XSTDFILL94_1688 VDD VSS sg13g2_FILL8
XSTDFILL94_1696 VDD VSS sg13g2_FILL8
XSTDFILL94_1704 VDD VSS sg13g2_FILL8
XSTDFILL94_1712 VDD VSS sg13g2_FILL8
XSTDFILL94_1720 VDD VSS sg13g2_FILL8
XSTDFILL94_1728 VDD VSS sg13g2_FILL8
XSTDFILL94_1736 VDD VSS sg13g2_FILL8
XSTDFILL94_1744 VDD VSS sg13g2_FILL8
XSTDFILL94_1752 VDD VSS sg13g2_FILL8
XSTDFILL94_1760 VDD VSS sg13g2_FILL8
XSTDFILL94_1768 VDD VSS sg13g2_FILL8
XSTDFILL94_1776 VDD VSS sg13g2_FILL8
XSTDFILL94_1784 VDD VSS sg13g2_FILL8
XSTDFILL94_1792 VDD VSS sg13g2_FILL8
XSTDFILL94_1800 VDD VSS sg13g2_FILL8
XSTDFILL94_1808 VDD VSS sg13g2_FILL8
XSTDFILL94_1816 VDD VSS sg13g2_FILL8
XSTDFILL94_1824 VDD VSS sg13g2_FILL8
XSTDFILL94_1832 VDD VSS sg13g2_FILL8
XSTDFILL94_1840 VDD VSS sg13g2_FILL8
XSTDFILL94_1848 VDD VSS sg13g2_FILL8
XSTDFILL94_1856 VDD VSS sg13g2_FILL8
XSTDFILL94_1864 VDD VSS sg13g2_FILL8
XSTDFILL94_1872 VDD VSS sg13g2_FILL8
XSTDFILL94_1880 VDD VSS sg13g2_FILL8
XSTDFILL94_1888 VDD VSS sg13g2_FILL8
XSTDFILL94_1896 VDD VSS sg13g2_FILL8
XSTDFILL94_1904 VDD VSS sg13g2_FILL8
XSTDFILL94_1912 VDD VSS sg13g2_FILL8
XSTDFILL94_1920 VDD VSS sg13g2_FILL8
XSTDFILL94_1928 VDD VSS sg13g2_FILL8
XSTDFILL94_1936 VDD VSS sg13g2_FILL8
XSTDFILL94_1944 VDD VSS sg13g2_FILL8
XSTDFILL94_1952 VDD VSS sg13g2_FILL8
XSTDFILL94_1960 VDD VSS sg13g2_FILL8
XSTDFILL94_1968 VDD VSS sg13g2_FILL8
XSTDFILL94_1976 VDD VSS sg13g2_FILL8
XSTDFILL94_1984 VDD VSS sg13g2_FILL8
XSTDFILL94_1992 VDD VSS sg13g2_FILL8
XSTDFILL94_2000 VDD VSS sg13g2_FILL8
XSTDFILL94_2008 VDD VSS sg13g2_FILL8
XSTDFILL94_2016 VDD VSS sg13g2_FILL8
XSTDFILL94_2024 VDD VSS sg13g2_FILL8
XSTDFILL94_2032 VDD VSS sg13g2_FILL8
XSTDFILL94_2040 VDD VSS sg13g2_FILL8
XSTDFILL94_2048 VDD VSS sg13g2_FILL8
XSTDFILL94_2056 VDD VSS sg13g2_FILL8
XSTDFILL94_2064 VDD VSS sg13g2_FILL8
XSTDFILL94_2072 VDD VSS sg13g2_FILL8
XSTDFILL94_2080 VDD VSS sg13g2_FILL8
XSTDFILL94_2088 VDD VSS sg13g2_FILL8
XSTDFILL94_2096 VDD VSS sg13g2_FILL8
XSTDFILL94_2104 VDD VSS sg13g2_FILL8
XSTDFILL94_2112 VDD VSS sg13g2_FILL8
XSTDFILL94_2120 VDD VSS sg13g2_FILL8
XSTDFILL94_2128 VDD VSS sg13g2_FILL8
XSTDFILL94_2136 VDD VSS sg13g2_FILL8
XSTDFILL94_2144 VDD VSS sg13g2_FILL8
XSTDFILL94_2152 VDD VSS sg13g2_FILL2
XSTDFILL95_0 VDD VSS sg13g2_FILL8
XSTDFILL95_8 VDD VSS sg13g2_FILL8
XSTDFILL95_16 VDD VSS sg13g2_FILL8
XSTDFILL95_24 VDD VSS sg13g2_FILL8
XSTDFILL95_32 VDD VSS sg13g2_FILL8
XSTDFILL95_40 VDD VSS sg13g2_FILL8
XSTDFILL95_48 VDD VSS sg13g2_FILL8
XSTDFILL95_56 VDD VSS sg13g2_FILL8
XSTDFILL95_64 VDD VSS sg13g2_FILL8
XSTDFILL95_72 VDD VSS sg13g2_FILL8
XSTDFILL95_80 VDD VSS sg13g2_FILL8
XSTDFILL95_88 VDD VSS sg13g2_FILL8
XSTDFILL95_96 VDD VSS sg13g2_FILL8
XSTDFILL95_104 VDD VSS sg13g2_FILL8
XSTDFILL95_112 VDD VSS sg13g2_FILL8
XSTDFILL95_120 VDD VSS sg13g2_FILL8
XSTDFILL95_128 VDD VSS sg13g2_FILL8
XSTDFILL95_136 VDD VSS sg13g2_FILL8
XSTDFILL95_144 VDD VSS sg13g2_FILL8
XSTDFILL95_152 VDD VSS sg13g2_FILL8
XSTDFILL95_160 VDD VSS sg13g2_FILL8
XSTDFILL95_168 VDD VSS sg13g2_FILL8
XSTDFILL95_176 VDD VSS sg13g2_FILL8
XSTDFILL95_184 VDD VSS sg13g2_FILL8
XSTDFILL95_192 VDD VSS sg13g2_FILL8
XSTDFILL95_200 VDD VSS sg13g2_FILL8
XSTDFILL95_208 VDD VSS sg13g2_FILL8
XSTDFILL95_216 VDD VSS sg13g2_FILL8
XSTDFILL95_224 VDD VSS sg13g2_FILL8
XSTDFILL95_232 VDD VSS sg13g2_FILL8
XSTDFILL95_240 VDD VSS sg13g2_FILL8
XSTDFILL95_248 VDD VSS sg13g2_FILL8
XSTDFILL95_256 VDD VSS sg13g2_FILL8
XSTDFILL95_264 VDD VSS sg13g2_FILL8
XSTDFILL95_272 VDD VSS sg13g2_FILL8
XSTDFILL95_280 VDD VSS sg13g2_FILL8
XSTDFILL95_288 VDD VSS sg13g2_FILL8
XSTDFILL95_296 VDD VSS sg13g2_FILL8
XSTDFILL95_304 VDD VSS sg13g2_FILL8
XSTDFILL95_312 VDD VSS sg13g2_FILL8
XSTDFILL95_320 VDD VSS sg13g2_FILL8
XSTDFILL95_328 VDD VSS sg13g2_FILL8
XSTDFILL95_336 VDD VSS sg13g2_FILL8
XSTDFILL95_344 VDD VSS sg13g2_FILL8
XSTDFILL95_352 VDD VSS sg13g2_FILL8
XSTDFILL95_360 VDD VSS sg13g2_FILL8
XSTDFILL95_368 VDD VSS sg13g2_FILL8
XSTDFILL95_376 VDD VSS sg13g2_FILL8
XSTDFILL95_384 VDD VSS sg13g2_FILL8
XSTDFILL95_392 VDD VSS sg13g2_FILL8
XSTDFILL95_400 VDD VSS sg13g2_FILL8
XSTDFILL95_408 VDD VSS sg13g2_FILL8
XSTDFILL95_416 VDD VSS sg13g2_FILL8
XSTDFILL95_424 VDD VSS sg13g2_FILL8
XSTDFILL95_432 VDD VSS sg13g2_FILL8
XSTDFILL95_440 VDD VSS sg13g2_FILL8
XSTDFILL95_448 VDD VSS sg13g2_FILL8
XSTDFILL95_456 VDD VSS sg13g2_FILL8
XSTDFILL95_464 VDD VSS sg13g2_FILL8
XSTDFILL95_472 VDD VSS sg13g2_FILL8
XSTDFILL95_480 VDD VSS sg13g2_FILL8
XSTDFILL95_488 VDD VSS sg13g2_FILL8
XSTDFILL95_496 VDD VSS sg13g2_FILL8
XSTDFILL95_504 VDD VSS sg13g2_FILL8
XSTDFILL95_512 VDD VSS sg13g2_FILL8
XSTDFILL95_520 VDD VSS sg13g2_FILL8
XSTDFILL95_528 VDD VSS sg13g2_FILL8
XSTDFILL95_536 VDD VSS sg13g2_FILL8
XSTDFILL95_544 VDD VSS sg13g2_FILL8
XSTDFILL95_552 VDD VSS sg13g2_FILL8
XSTDFILL95_560 VDD VSS sg13g2_FILL8
XSTDFILL95_568 VDD VSS sg13g2_FILL8
XSTDFILL95_576 VDD VSS sg13g2_FILL8
XSTDFILL95_584 VDD VSS sg13g2_FILL8
XSTDFILL95_592 VDD VSS sg13g2_FILL8
XSTDFILL95_600 VDD VSS sg13g2_FILL8
XSTDFILL95_608 VDD VSS sg13g2_FILL8
XSTDFILL95_616 VDD VSS sg13g2_FILL8
XSTDFILL95_624 VDD VSS sg13g2_FILL8
XSTDFILL95_632 VDD VSS sg13g2_FILL8
XSTDFILL95_640 VDD VSS sg13g2_FILL8
XSTDFILL95_648 VDD VSS sg13g2_FILL8
XSTDFILL95_656 VDD VSS sg13g2_FILL8
XSTDFILL95_664 VDD VSS sg13g2_FILL8
XSTDFILL95_672 VDD VSS sg13g2_FILL8
XSTDFILL95_680 VDD VSS sg13g2_FILL8
XSTDFILL95_688 VDD VSS sg13g2_FILL8
XSTDFILL95_696 VDD VSS sg13g2_FILL8
XSTDFILL95_704 VDD VSS sg13g2_FILL8
XSTDFILL95_712 VDD VSS sg13g2_FILL8
XSTDFILL95_720 VDD VSS sg13g2_FILL8
XSTDFILL95_728 VDD VSS sg13g2_FILL8
XSTDFILL95_736 VDD VSS sg13g2_FILL8
XSTDFILL95_744 VDD VSS sg13g2_FILL8
XSTDFILL95_752 VDD VSS sg13g2_FILL8
XSTDFILL95_760 VDD VSS sg13g2_FILL8
XSTDFILL95_768 VDD VSS sg13g2_FILL8
XSTDFILL95_776 VDD VSS sg13g2_FILL8
XSTDFILL95_784 VDD VSS sg13g2_FILL8
XSTDFILL95_792 VDD VSS sg13g2_FILL8
XSTDFILL95_800 VDD VSS sg13g2_FILL8
XSTDFILL95_808 VDD VSS sg13g2_FILL8
XSTDFILL95_816 VDD VSS sg13g2_FILL8
XSTDFILL95_824 VDD VSS sg13g2_FILL8
XSTDFILL95_832 VDD VSS sg13g2_FILL8
XSTDFILL95_840 VDD VSS sg13g2_FILL8
XSTDFILL95_848 VDD VSS sg13g2_FILL8
XSTDFILL95_856 VDD VSS sg13g2_FILL8
XSTDFILL95_864 VDD VSS sg13g2_FILL8
XSTDFILL95_872 VDD VSS sg13g2_FILL8
XSTDFILL95_880 VDD VSS sg13g2_FILL8
XSTDFILL95_888 VDD VSS sg13g2_FILL8
XSTDFILL95_896 VDD VSS sg13g2_FILL8
XSTDFILL95_904 VDD VSS sg13g2_FILL8
XSTDFILL95_912 VDD VSS sg13g2_FILL8
XSTDFILL95_920 VDD VSS sg13g2_FILL8
XSTDFILL95_928 VDD VSS sg13g2_FILL8
XSTDFILL95_936 VDD VSS sg13g2_FILL8
XSTDFILL95_944 VDD VSS sg13g2_FILL8
XSTDFILL95_952 VDD VSS sg13g2_FILL8
XSTDFILL95_960 VDD VSS sg13g2_FILL8
XSTDFILL95_968 VDD VSS sg13g2_FILL8
XSTDFILL95_976 VDD VSS sg13g2_FILL8
XSTDFILL95_984 VDD VSS sg13g2_FILL8
XSTDFILL95_992 VDD VSS sg13g2_FILL8
XSTDFILL95_1000 VDD VSS sg13g2_FILL8
XSTDFILL95_1008 VDD VSS sg13g2_FILL8
XSTDFILL95_1016 VDD VSS sg13g2_FILL8
XSTDFILL95_1024 VDD VSS sg13g2_FILL8
XSTDFILL95_1032 VDD VSS sg13g2_FILL8
XSTDFILL95_1040 VDD VSS sg13g2_FILL8
XSTDFILL95_1048 VDD VSS sg13g2_FILL8
XSTDFILL95_1056 VDD VSS sg13g2_FILL8
XSTDFILL95_1064 VDD VSS sg13g2_FILL8
XSTDFILL95_1072 VDD VSS sg13g2_FILL8
XSTDFILL95_1080 VDD VSS sg13g2_FILL8
XSTDFILL95_1088 VDD VSS sg13g2_FILL8
XSTDFILL95_1096 VDD VSS sg13g2_FILL8
XSTDFILL95_1104 VDD VSS sg13g2_FILL8
XSTDFILL95_1112 VDD VSS sg13g2_FILL8
XSTDFILL95_1120 VDD VSS sg13g2_FILL8
XSTDFILL95_1128 VDD VSS sg13g2_FILL8
XSTDFILL95_1136 VDD VSS sg13g2_FILL8
XSTDFILL95_1144 VDD VSS sg13g2_FILL8
XSTDFILL95_1152 VDD VSS sg13g2_FILL8
XSTDFILL95_1160 VDD VSS sg13g2_FILL8
XSTDFILL95_1168 VDD VSS sg13g2_FILL8
XSTDFILL95_1176 VDD VSS sg13g2_FILL8
XSTDFILL95_1184 VDD VSS sg13g2_FILL8
XSTDFILL95_1192 VDD VSS sg13g2_FILL8
XSTDFILL95_1200 VDD VSS sg13g2_FILL8
XSTDFILL95_1208 VDD VSS sg13g2_FILL8
XSTDFILL95_1216 VDD VSS sg13g2_FILL8
XSTDFILL95_1224 VDD VSS sg13g2_FILL8
XSTDFILL95_1232 VDD VSS sg13g2_FILL8
XSTDFILL95_1240 VDD VSS sg13g2_FILL8
XSTDFILL95_1248 VDD VSS sg13g2_FILL8
XSTDFILL95_1256 VDD VSS sg13g2_FILL8
XSTDFILL95_1264 VDD VSS sg13g2_FILL8
XSTDFILL95_1272 VDD VSS sg13g2_FILL8
XSTDFILL95_1280 VDD VSS sg13g2_FILL8
XSTDFILL95_1288 VDD VSS sg13g2_FILL8
XSTDFILL95_1296 VDD VSS sg13g2_FILL8
XSTDFILL95_1304 VDD VSS sg13g2_FILL8
XSTDFILL95_1312 VDD VSS sg13g2_FILL8
XSTDFILL95_1320 VDD VSS sg13g2_FILL8
XSTDFILL95_1328 VDD VSS sg13g2_FILL8
XSTDFILL95_1336 VDD VSS sg13g2_FILL8
XSTDFILL95_1344 VDD VSS sg13g2_FILL8
XSTDFILL95_1352 VDD VSS sg13g2_FILL8
XSTDFILL95_1360 VDD VSS sg13g2_FILL8
XSTDFILL95_1368 VDD VSS sg13g2_FILL8
XSTDFILL95_1376 VDD VSS sg13g2_FILL8
XSTDFILL95_1384 VDD VSS sg13g2_FILL8
XSTDFILL95_1392 VDD VSS sg13g2_FILL8
XSTDFILL95_1400 VDD VSS sg13g2_FILL8
XSTDFILL95_1408 VDD VSS sg13g2_FILL8
XSTDFILL95_1416 VDD VSS sg13g2_FILL8
XSTDFILL95_1424 VDD VSS sg13g2_FILL8
XSTDFILL95_1432 VDD VSS sg13g2_FILL8
XSTDFILL95_1440 VDD VSS sg13g2_FILL8
XSTDFILL95_1448 VDD VSS sg13g2_FILL8
XSTDFILL95_1456 VDD VSS sg13g2_FILL8
XSTDFILL95_1464 VDD VSS sg13g2_FILL8
XSTDFILL95_1472 VDD VSS sg13g2_FILL8
XSTDFILL95_1480 VDD VSS sg13g2_FILL8
XSTDFILL95_1488 VDD VSS sg13g2_FILL8
XSTDFILL95_1496 VDD VSS sg13g2_FILL8
XSTDFILL95_1504 VDD VSS sg13g2_FILL8
XSTDFILL95_1512 VDD VSS sg13g2_FILL8
XSTDFILL95_1520 VDD VSS sg13g2_FILL8
XSTDFILL95_1528 VDD VSS sg13g2_FILL8
XSTDFILL95_1536 VDD VSS sg13g2_FILL8
XSTDFILL95_1544 VDD VSS sg13g2_FILL8
XSTDFILL95_1552 VDD VSS sg13g2_FILL8
XSTDFILL95_1560 VDD VSS sg13g2_FILL8
XSTDFILL95_1568 VDD VSS sg13g2_FILL8
XSTDFILL95_1576 VDD VSS sg13g2_FILL8
XSTDFILL95_1584 VDD VSS sg13g2_FILL8
XSTDFILL95_1592 VDD VSS sg13g2_FILL8
XSTDFILL95_1600 VDD VSS sg13g2_FILL8
XSTDFILL95_1608 VDD VSS sg13g2_FILL8
XSTDFILL95_1616 VDD VSS sg13g2_FILL8
XSTDFILL95_1624 VDD VSS sg13g2_FILL8
XSTDFILL95_1632 VDD VSS sg13g2_FILL8
XSTDFILL95_1640 VDD VSS sg13g2_FILL8
XSTDFILL95_1648 VDD VSS sg13g2_FILL8
XSTDFILL95_1656 VDD VSS sg13g2_FILL8
XSTDFILL95_1664 VDD VSS sg13g2_FILL8
XSTDFILL95_1672 VDD VSS sg13g2_FILL8
XSTDFILL95_1680 VDD VSS sg13g2_FILL8
XSTDFILL95_1688 VDD VSS sg13g2_FILL8
XSTDFILL95_1696 VDD VSS sg13g2_FILL8
XSTDFILL95_1704 VDD VSS sg13g2_FILL8
XSTDFILL95_1712 VDD VSS sg13g2_FILL8
XSTDFILL95_1720 VDD VSS sg13g2_FILL8
XSTDFILL95_1728 VDD VSS sg13g2_FILL8
XSTDFILL95_1736 VDD VSS sg13g2_FILL8
XSTDFILL95_1744 VDD VSS sg13g2_FILL8
XSTDFILL95_1752 VDD VSS sg13g2_FILL8
XSTDFILL95_1760 VDD VSS sg13g2_FILL8
XSTDFILL95_1768 VDD VSS sg13g2_FILL8
XSTDFILL95_1776 VDD VSS sg13g2_FILL8
XSTDFILL95_1784 VDD VSS sg13g2_FILL8
XSTDFILL95_1792 VDD VSS sg13g2_FILL8
XSTDFILL95_1800 VDD VSS sg13g2_FILL8
XSTDFILL95_1808 VDD VSS sg13g2_FILL8
XSTDFILL95_1816 VDD VSS sg13g2_FILL8
XSTDFILL95_1824 VDD VSS sg13g2_FILL8
XSTDFILL95_1832 VDD VSS sg13g2_FILL8
XSTDFILL95_1840 VDD VSS sg13g2_FILL8
XSTDFILL95_1848 VDD VSS sg13g2_FILL8
XSTDFILL95_1856 VDD VSS sg13g2_FILL8
XSTDFILL95_1864 VDD VSS sg13g2_FILL8
XSTDFILL95_1872 VDD VSS sg13g2_FILL8
XSTDFILL95_1880 VDD VSS sg13g2_FILL8
XSTDFILL95_1888 VDD VSS sg13g2_FILL8
XSTDFILL95_1896 VDD VSS sg13g2_FILL8
XSTDFILL95_1904 VDD VSS sg13g2_FILL8
XSTDFILL95_1912 VDD VSS sg13g2_FILL8
XSTDFILL95_1920 VDD VSS sg13g2_FILL8
XSTDFILL95_1928 VDD VSS sg13g2_FILL8
XSTDFILL95_1936 VDD VSS sg13g2_FILL8
XSTDFILL95_1944 VDD VSS sg13g2_FILL8
XSTDFILL95_1952 VDD VSS sg13g2_FILL8
XSTDFILL95_1960 VDD VSS sg13g2_FILL8
XSTDFILL95_1968 VDD VSS sg13g2_FILL8
XSTDFILL95_1976 VDD VSS sg13g2_FILL8
XSTDFILL95_1984 VDD VSS sg13g2_FILL8
XSTDFILL95_1992 VDD VSS sg13g2_FILL8
XSTDFILL95_2000 VDD VSS sg13g2_FILL8
XSTDFILL95_2008 VDD VSS sg13g2_FILL8
XSTDFILL95_2016 VDD VSS sg13g2_FILL8
XSTDFILL95_2024 VDD VSS sg13g2_FILL8
XSTDFILL95_2032 VDD VSS sg13g2_FILL8
XSTDFILL95_2040 VDD VSS sg13g2_FILL8
XSTDFILL95_2048 VDD VSS sg13g2_FILL8
XSTDFILL95_2056 VDD VSS sg13g2_FILL8
XSTDFILL95_2064 VDD VSS sg13g2_FILL8
XSTDFILL95_2072 VDD VSS sg13g2_FILL8
XSTDFILL95_2080 VDD VSS sg13g2_FILL8
XSTDFILL95_2088 VDD VSS sg13g2_FILL8
XSTDFILL95_2096 VDD VSS sg13g2_FILL8
XSTDFILL95_2104 VDD VSS sg13g2_FILL8
XSTDFILL95_2112 VDD VSS sg13g2_FILL8
XSTDFILL95_2120 VDD VSS sg13g2_FILL8
XSTDFILL95_2128 VDD VSS sg13g2_FILL8
XSTDFILL95_2136 VDD VSS sg13g2_FILL8
XSTDFILL95_2144 VDD VSS sg13g2_FILL8
XSTDFILL95_2152 VDD VSS sg13g2_FILL2
XSTDFILL96_0 VDD VSS sg13g2_FILL8
XSTDFILL96_8 VDD VSS sg13g2_FILL8
XSTDFILL96_16 VDD VSS sg13g2_FILL8
XSTDFILL96_24 VDD VSS sg13g2_FILL8
XSTDFILL96_32 VDD VSS sg13g2_FILL8
XSTDFILL96_40 VDD VSS sg13g2_FILL8
XSTDFILL96_48 VDD VSS sg13g2_FILL8
XSTDFILL96_56 VDD VSS sg13g2_FILL8
XSTDFILL96_64 VDD VSS sg13g2_FILL8
XSTDFILL96_72 VDD VSS sg13g2_FILL8
XSTDFILL96_80 VDD VSS sg13g2_FILL8
XSTDFILL96_88 VDD VSS sg13g2_FILL8
XSTDFILL96_96 VDD VSS sg13g2_FILL8
XSTDFILL96_104 VDD VSS sg13g2_FILL8
XSTDFILL96_112 VDD VSS sg13g2_FILL8
XSTDFILL96_120 VDD VSS sg13g2_FILL8
XSTDFILL96_128 VDD VSS sg13g2_FILL8
XSTDFILL96_136 VDD VSS sg13g2_FILL8
XSTDFILL96_144 VDD VSS sg13g2_FILL8
XSTDFILL96_152 VDD VSS sg13g2_FILL8
XSTDFILL96_160 VDD VSS sg13g2_FILL8
XSTDFILL96_168 VDD VSS sg13g2_FILL8
XSTDFILL96_176 VDD VSS sg13g2_FILL8
XSTDFILL96_184 VDD VSS sg13g2_FILL8
XSTDFILL96_192 VDD VSS sg13g2_FILL8
XSTDFILL96_200 VDD VSS sg13g2_FILL8
XSTDFILL96_208 VDD VSS sg13g2_FILL8
XSTDFILL96_216 VDD VSS sg13g2_FILL8
XSTDFILL96_224 VDD VSS sg13g2_FILL8
XSTDFILL96_232 VDD VSS sg13g2_FILL8
XSTDFILL96_240 VDD VSS sg13g2_FILL8
XSTDFILL96_248 VDD VSS sg13g2_FILL8
XSTDFILL96_256 VDD VSS sg13g2_FILL8
XSTDFILL96_264 VDD VSS sg13g2_FILL8
XSTDFILL96_272 VDD VSS sg13g2_FILL8
XSTDFILL96_280 VDD VSS sg13g2_FILL8
XSTDFILL96_288 VDD VSS sg13g2_FILL8
XSTDFILL96_296 VDD VSS sg13g2_FILL8
XSTDFILL96_304 VDD VSS sg13g2_FILL8
XSTDFILL96_312 VDD VSS sg13g2_FILL8
XSTDFILL96_320 VDD VSS sg13g2_FILL8
XSTDFILL96_328 VDD VSS sg13g2_FILL8
XSTDFILL96_336 VDD VSS sg13g2_FILL8
XSTDFILL96_344 VDD VSS sg13g2_FILL8
XSTDFILL96_352 VDD VSS sg13g2_FILL8
XSTDFILL96_360 VDD VSS sg13g2_FILL8
XSTDFILL96_368 VDD VSS sg13g2_FILL8
XSTDFILL96_376 VDD VSS sg13g2_FILL8
XSTDFILL96_384 VDD VSS sg13g2_FILL8
XSTDFILL96_392 VDD VSS sg13g2_FILL8
XSTDFILL96_400 VDD VSS sg13g2_FILL8
XSTDFILL96_408 VDD VSS sg13g2_FILL8
XSTDFILL96_416 VDD VSS sg13g2_FILL8
XSTDFILL96_424 VDD VSS sg13g2_FILL8
XSTDFILL96_432 VDD VSS sg13g2_FILL8
XSTDFILL96_440 VDD VSS sg13g2_FILL8
XSTDFILL96_448 VDD VSS sg13g2_FILL8
XSTDFILL96_456 VDD VSS sg13g2_FILL8
XSTDFILL96_464 VDD VSS sg13g2_FILL8
XSTDFILL96_472 VDD VSS sg13g2_FILL8
XSTDFILL96_480 VDD VSS sg13g2_FILL8
XSTDFILL96_488 VDD VSS sg13g2_FILL8
XSTDFILL96_496 VDD VSS sg13g2_FILL8
XSTDFILL96_504 VDD VSS sg13g2_FILL8
XSTDFILL96_512 VDD VSS sg13g2_FILL8
XSTDFILL96_520 VDD VSS sg13g2_FILL8
XSTDFILL96_528 VDD VSS sg13g2_FILL8
XSTDFILL96_536 VDD VSS sg13g2_FILL8
XSTDFILL96_544 VDD VSS sg13g2_FILL8
XSTDFILL96_552 VDD VSS sg13g2_FILL8
XSTDFILL96_560 VDD VSS sg13g2_FILL8
XSTDFILL96_568 VDD VSS sg13g2_FILL8
XSTDFILL96_576 VDD VSS sg13g2_FILL8
XSTDFILL96_584 VDD VSS sg13g2_FILL8
XSTDFILL96_592 VDD VSS sg13g2_FILL8
XSTDFILL96_600 VDD VSS sg13g2_FILL8
XSTDFILL96_608 VDD VSS sg13g2_FILL8
XSTDFILL96_616 VDD VSS sg13g2_FILL8
XSTDFILL96_624 VDD VSS sg13g2_FILL8
XSTDFILL96_632 VDD VSS sg13g2_FILL8
XSTDFILL96_640 VDD VSS sg13g2_FILL8
XSTDFILL96_648 VDD VSS sg13g2_FILL8
XSTDFILL96_656 VDD VSS sg13g2_FILL8
XSTDFILL96_664 VDD VSS sg13g2_FILL8
XSTDFILL96_672 VDD VSS sg13g2_FILL8
XSTDFILL96_680 VDD VSS sg13g2_FILL8
XSTDFILL96_688 VDD VSS sg13g2_FILL8
XSTDFILL96_696 VDD VSS sg13g2_FILL8
XSTDFILL96_704 VDD VSS sg13g2_FILL8
XSTDFILL96_712 VDD VSS sg13g2_FILL8
XSTDFILL96_720 VDD VSS sg13g2_FILL8
XSTDFILL96_728 VDD VSS sg13g2_FILL8
XSTDFILL96_736 VDD VSS sg13g2_FILL8
XSTDFILL96_744 VDD VSS sg13g2_FILL8
XSTDFILL96_752 VDD VSS sg13g2_FILL8
XSTDFILL96_760 VDD VSS sg13g2_FILL8
XSTDFILL96_768 VDD VSS sg13g2_FILL8
XSTDFILL96_776 VDD VSS sg13g2_FILL8
XSTDFILL96_784 VDD VSS sg13g2_FILL8
XSTDFILL96_792 VDD VSS sg13g2_FILL8
XSTDFILL96_800 VDD VSS sg13g2_FILL8
XSTDFILL96_808 VDD VSS sg13g2_FILL8
XSTDFILL96_816 VDD VSS sg13g2_FILL8
XSTDFILL96_824 VDD VSS sg13g2_FILL8
XSTDFILL96_832 VDD VSS sg13g2_FILL8
XSTDFILL96_840 VDD VSS sg13g2_FILL8
XSTDFILL96_848 VDD VSS sg13g2_FILL8
XSTDFILL96_856 VDD VSS sg13g2_FILL8
XSTDFILL96_864 VDD VSS sg13g2_FILL8
XSTDFILL96_872 VDD VSS sg13g2_FILL8
XSTDFILL96_880 VDD VSS sg13g2_FILL8
XSTDFILL96_888 VDD VSS sg13g2_FILL8
XSTDFILL96_896 VDD VSS sg13g2_FILL8
XSTDFILL96_904 VDD VSS sg13g2_FILL8
XSTDFILL96_912 VDD VSS sg13g2_FILL8
XSTDFILL96_920 VDD VSS sg13g2_FILL8
XSTDFILL96_928 VDD VSS sg13g2_FILL8
XSTDFILL96_936 VDD VSS sg13g2_FILL8
XSTDFILL96_944 VDD VSS sg13g2_FILL8
XSTDFILL96_952 VDD VSS sg13g2_FILL8
XSTDFILL96_960 VDD VSS sg13g2_FILL8
XSTDFILL96_968 VDD VSS sg13g2_FILL8
XSTDFILL96_976 VDD VSS sg13g2_FILL8
XSTDFILL96_984 VDD VSS sg13g2_FILL8
XSTDFILL96_992 VDD VSS sg13g2_FILL8
XSTDFILL96_1000 VDD VSS sg13g2_FILL8
XSTDFILL96_1008 VDD VSS sg13g2_FILL8
XSTDFILL96_1016 VDD VSS sg13g2_FILL8
XSTDFILL96_1024 VDD VSS sg13g2_FILL8
XSTDFILL96_1032 VDD VSS sg13g2_FILL8
XSTDFILL96_1040 VDD VSS sg13g2_FILL8
XSTDFILL96_1048 VDD VSS sg13g2_FILL8
XSTDFILL96_1056 VDD VSS sg13g2_FILL8
XSTDFILL96_1064 VDD VSS sg13g2_FILL8
XSTDFILL96_1072 VDD VSS sg13g2_FILL8
XSTDFILL96_1080 VDD VSS sg13g2_FILL8
XSTDFILL96_1088 VDD VSS sg13g2_FILL8
XSTDFILL96_1096 VDD VSS sg13g2_FILL8
XSTDFILL96_1104 VDD VSS sg13g2_FILL8
XSTDFILL96_1112 VDD VSS sg13g2_FILL8
XSTDFILL96_1120 VDD VSS sg13g2_FILL8
XSTDFILL96_1128 VDD VSS sg13g2_FILL8
XSTDFILL96_1136 VDD VSS sg13g2_FILL8
XSTDFILL96_1144 VDD VSS sg13g2_FILL8
XSTDFILL96_1152 VDD VSS sg13g2_FILL8
XSTDFILL96_1160 VDD VSS sg13g2_FILL8
XSTDFILL96_1168 VDD VSS sg13g2_FILL8
XSTDFILL96_1176 VDD VSS sg13g2_FILL8
XSTDFILL96_1184 VDD VSS sg13g2_FILL8
XSTDFILL96_1192 VDD VSS sg13g2_FILL8
XSTDFILL96_1200 VDD VSS sg13g2_FILL8
XSTDFILL96_1208 VDD VSS sg13g2_FILL8
XSTDFILL96_1216 VDD VSS sg13g2_FILL8
XSTDFILL96_1224 VDD VSS sg13g2_FILL8
XSTDFILL96_1232 VDD VSS sg13g2_FILL8
XSTDFILL96_1240 VDD VSS sg13g2_FILL8
XSTDFILL96_1248 VDD VSS sg13g2_FILL8
XSTDFILL96_1256 VDD VSS sg13g2_FILL8
XSTDFILL96_1264 VDD VSS sg13g2_FILL8
XSTDFILL96_1272 VDD VSS sg13g2_FILL8
XSTDFILL96_1280 VDD VSS sg13g2_FILL8
XSTDFILL96_1288 VDD VSS sg13g2_FILL8
XSTDFILL96_1296 VDD VSS sg13g2_FILL8
XSTDFILL96_1304 VDD VSS sg13g2_FILL8
XSTDFILL96_1312 VDD VSS sg13g2_FILL8
XSTDFILL96_1320 VDD VSS sg13g2_FILL8
XSTDFILL96_1328 VDD VSS sg13g2_FILL8
XSTDFILL96_1336 VDD VSS sg13g2_FILL8
XSTDFILL96_1344 VDD VSS sg13g2_FILL8
XSTDFILL96_1352 VDD VSS sg13g2_FILL8
XSTDFILL96_1360 VDD VSS sg13g2_FILL8
XSTDFILL96_1368 VDD VSS sg13g2_FILL8
XSTDFILL96_1376 VDD VSS sg13g2_FILL8
XSTDFILL96_1384 VDD VSS sg13g2_FILL8
XSTDFILL96_1392 VDD VSS sg13g2_FILL8
XSTDFILL96_1400 VDD VSS sg13g2_FILL8
XSTDFILL96_1408 VDD VSS sg13g2_FILL8
XSTDFILL96_1416 VDD VSS sg13g2_FILL8
XSTDFILL96_1424 VDD VSS sg13g2_FILL8
XSTDFILL96_1432 VDD VSS sg13g2_FILL8
XSTDFILL96_1440 VDD VSS sg13g2_FILL8
XSTDFILL96_1448 VDD VSS sg13g2_FILL8
XSTDFILL96_1456 VDD VSS sg13g2_FILL8
XSTDFILL96_1464 VDD VSS sg13g2_FILL8
XSTDFILL96_1472 VDD VSS sg13g2_FILL8
XSTDFILL96_1480 VDD VSS sg13g2_FILL8
XSTDFILL96_1488 VDD VSS sg13g2_FILL8
XSTDFILL96_1496 VDD VSS sg13g2_FILL8
XSTDFILL96_1504 VDD VSS sg13g2_FILL8
XSTDFILL96_1512 VDD VSS sg13g2_FILL8
XSTDFILL96_1520 VDD VSS sg13g2_FILL8
XSTDFILL96_1528 VDD VSS sg13g2_FILL8
XSTDFILL96_1536 VDD VSS sg13g2_FILL8
XSTDFILL96_1544 VDD VSS sg13g2_FILL8
XSTDFILL96_1552 VDD VSS sg13g2_FILL8
XSTDFILL96_1560 VDD VSS sg13g2_FILL8
XSTDFILL96_1568 VDD VSS sg13g2_FILL8
XSTDFILL96_1576 VDD VSS sg13g2_FILL8
XSTDFILL96_1584 VDD VSS sg13g2_FILL8
XSTDFILL96_1592 VDD VSS sg13g2_FILL8
XSTDFILL96_1600 VDD VSS sg13g2_FILL8
XSTDFILL96_1608 VDD VSS sg13g2_FILL8
XSTDFILL96_1616 VDD VSS sg13g2_FILL8
XSTDFILL96_1624 VDD VSS sg13g2_FILL8
XSTDFILL96_1632 VDD VSS sg13g2_FILL8
XSTDFILL96_1640 VDD VSS sg13g2_FILL8
XSTDFILL96_1648 VDD VSS sg13g2_FILL8
XSTDFILL96_1656 VDD VSS sg13g2_FILL8
XSTDFILL96_1664 VDD VSS sg13g2_FILL8
XSTDFILL96_1672 VDD VSS sg13g2_FILL8
XSTDFILL96_1680 VDD VSS sg13g2_FILL8
XSTDFILL96_1688 VDD VSS sg13g2_FILL8
XSTDFILL96_1696 VDD VSS sg13g2_FILL8
XSTDFILL96_1704 VDD VSS sg13g2_FILL8
XSTDFILL96_1712 VDD VSS sg13g2_FILL8
XSTDFILL96_1720 VDD VSS sg13g2_FILL8
XSTDFILL96_1728 VDD VSS sg13g2_FILL8
XSTDFILL96_1736 VDD VSS sg13g2_FILL8
XSTDFILL96_1744 VDD VSS sg13g2_FILL8
XSTDFILL96_1752 VDD VSS sg13g2_FILL8
XSTDFILL96_1760 VDD VSS sg13g2_FILL8
XSTDFILL96_1768 VDD VSS sg13g2_FILL8
XSTDFILL96_1776 VDD VSS sg13g2_FILL8
XSTDFILL96_1784 VDD VSS sg13g2_FILL8
XSTDFILL96_1792 VDD VSS sg13g2_FILL8
XSTDFILL96_1800 VDD VSS sg13g2_FILL8
XSTDFILL96_1808 VDD VSS sg13g2_FILL8
XSTDFILL96_1816 VDD VSS sg13g2_FILL8
XSTDFILL96_1824 VDD VSS sg13g2_FILL8
XSTDFILL96_1832 VDD VSS sg13g2_FILL8
XSTDFILL96_1840 VDD VSS sg13g2_FILL8
XSTDFILL96_1848 VDD VSS sg13g2_FILL8
XSTDFILL96_1856 VDD VSS sg13g2_FILL8
XSTDFILL96_1864 VDD VSS sg13g2_FILL8
XSTDFILL96_1872 VDD VSS sg13g2_FILL8
XSTDFILL96_1880 VDD VSS sg13g2_FILL8
XSTDFILL96_1888 VDD VSS sg13g2_FILL8
XSTDFILL96_1896 VDD VSS sg13g2_FILL8
XSTDFILL96_1904 VDD VSS sg13g2_FILL8
XSTDFILL96_1912 VDD VSS sg13g2_FILL8
XSTDFILL96_1920 VDD VSS sg13g2_FILL8
XSTDFILL96_1928 VDD VSS sg13g2_FILL8
XSTDFILL96_1936 VDD VSS sg13g2_FILL8
XSTDFILL96_1944 VDD VSS sg13g2_FILL8
XSTDFILL96_1952 VDD VSS sg13g2_FILL8
XSTDFILL96_1960 VDD VSS sg13g2_FILL8
XSTDFILL96_1968 VDD VSS sg13g2_FILL8
XSTDFILL96_1976 VDD VSS sg13g2_FILL8
XSTDFILL96_1984 VDD VSS sg13g2_FILL8
XSTDFILL96_1992 VDD VSS sg13g2_FILL8
XSTDFILL96_2000 VDD VSS sg13g2_FILL8
XSTDFILL96_2008 VDD VSS sg13g2_FILL8
XSTDFILL96_2016 VDD VSS sg13g2_FILL8
XSTDFILL96_2024 VDD VSS sg13g2_FILL8
XSTDFILL96_2032 VDD VSS sg13g2_FILL8
XSTDFILL96_2040 VDD VSS sg13g2_FILL8
XSTDFILL96_2048 VDD VSS sg13g2_FILL8
XSTDFILL96_2056 VDD VSS sg13g2_FILL8
XSTDFILL96_2064 VDD VSS sg13g2_FILL8
XSTDFILL96_2072 VDD VSS sg13g2_FILL8
XSTDFILL96_2080 VDD VSS sg13g2_FILL8
XSTDFILL96_2088 VDD VSS sg13g2_FILL8
XSTDFILL96_2096 VDD VSS sg13g2_FILL8
XSTDFILL96_2104 VDD VSS sg13g2_FILL8
XSTDFILL96_2112 VDD VSS sg13g2_FILL8
XSTDFILL96_2120 VDD VSS sg13g2_FILL8
XSTDFILL96_2128 VDD VSS sg13g2_FILL8
XSTDFILL96_2136 VDD VSS sg13g2_FILL8
XSTDFILL96_2144 VDD VSS sg13g2_FILL8
XSTDFILL96_2152 VDD VSS sg13g2_FILL2
XSTDFILL97_0 VDD VSS sg13g2_FILL8
XSTDFILL97_8 VDD VSS sg13g2_FILL8
XSTDFILL97_16 VDD VSS sg13g2_FILL8
XSTDFILL97_24 VDD VSS sg13g2_FILL8
XSTDFILL97_32 VDD VSS sg13g2_FILL8
XSTDFILL97_40 VDD VSS sg13g2_FILL8
XSTDFILL97_48 VDD VSS sg13g2_FILL8
XSTDFILL97_56 VDD VSS sg13g2_FILL8
XSTDFILL97_64 VDD VSS sg13g2_FILL8
XSTDFILL97_72 VDD VSS sg13g2_FILL8
XSTDFILL97_80 VDD VSS sg13g2_FILL8
XSTDFILL97_88 VDD VSS sg13g2_FILL8
XSTDFILL97_96 VDD VSS sg13g2_FILL8
XSTDFILL97_104 VDD VSS sg13g2_FILL8
XSTDFILL97_112 VDD VSS sg13g2_FILL8
XSTDFILL97_120 VDD VSS sg13g2_FILL8
XSTDFILL97_128 VDD VSS sg13g2_FILL8
XSTDFILL97_136 VDD VSS sg13g2_FILL8
XSTDFILL97_144 VDD VSS sg13g2_FILL8
XSTDFILL97_152 VDD VSS sg13g2_FILL8
XSTDFILL97_160 VDD VSS sg13g2_FILL8
XSTDFILL97_168 VDD VSS sg13g2_FILL8
XSTDFILL97_176 VDD VSS sg13g2_FILL8
XSTDFILL97_184 VDD VSS sg13g2_FILL8
XSTDFILL97_192 VDD VSS sg13g2_FILL8
XSTDFILL97_200 VDD VSS sg13g2_FILL8
XSTDFILL97_208 VDD VSS sg13g2_FILL8
XSTDFILL97_216 VDD VSS sg13g2_FILL8
XSTDFILL97_224 VDD VSS sg13g2_FILL8
XSTDFILL97_232 VDD VSS sg13g2_FILL8
XSTDFILL97_240 VDD VSS sg13g2_FILL8
XSTDFILL97_248 VDD VSS sg13g2_FILL8
XSTDFILL97_256 VDD VSS sg13g2_FILL8
XSTDFILL97_264 VDD VSS sg13g2_FILL8
XSTDFILL97_272 VDD VSS sg13g2_FILL8
XSTDFILL97_280 VDD VSS sg13g2_FILL8
XSTDFILL97_288 VDD VSS sg13g2_FILL8
XSTDFILL97_296 VDD VSS sg13g2_FILL8
XSTDFILL97_304 VDD VSS sg13g2_FILL8
XSTDFILL97_312 VDD VSS sg13g2_FILL8
XSTDFILL97_320 VDD VSS sg13g2_FILL8
XSTDFILL97_328 VDD VSS sg13g2_FILL8
XSTDFILL97_336 VDD VSS sg13g2_FILL8
XSTDFILL97_344 VDD VSS sg13g2_FILL8
XSTDFILL97_352 VDD VSS sg13g2_FILL8
XSTDFILL97_360 VDD VSS sg13g2_FILL8
XSTDFILL97_368 VDD VSS sg13g2_FILL8
XSTDFILL97_376 VDD VSS sg13g2_FILL8
XSTDFILL97_384 VDD VSS sg13g2_FILL8
XSTDFILL97_392 VDD VSS sg13g2_FILL8
XSTDFILL97_400 VDD VSS sg13g2_FILL8
XSTDFILL97_408 VDD VSS sg13g2_FILL8
XSTDFILL97_416 VDD VSS sg13g2_FILL8
XSTDFILL97_424 VDD VSS sg13g2_FILL8
XSTDFILL97_432 VDD VSS sg13g2_FILL8
XSTDFILL97_440 VDD VSS sg13g2_FILL8
XSTDFILL97_448 VDD VSS sg13g2_FILL8
XSTDFILL97_456 VDD VSS sg13g2_FILL8
XSTDFILL97_464 VDD VSS sg13g2_FILL8
XSTDFILL97_472 VDD VSS sg13g2_FILL8
XSTDFILL97_480 VDD VSS sg13g2_FILL8
XSTDFILL97_488 VDD VSS sg13g2_FILL8
XSTDFILL97_496 VDD VSS sg13g2_FILL8
XSTDFILL97_504 VDD VSS sg13g2_FILL8
XSTDFILL97_512 VDD VSS sg13g2_FILL8
XSTDFILL97_520 VDD VSS sg13g2_FILL8
XSTDFILL97_528 VDD VSS sg13g2_FILL8
XSTDFILL97_536 VDD VSS sg13g2_FILL8
XSTDFILL97_544 VDD VSS sg13g2_FILL8
XSTDFILL97_552 VDD VSS sg13g2_FILL8
XSTDFILL97_560 VDD VSS sg13g2_FILL8
XSTDFILL97_568 VDD VSS sg13g2_FILL8
XSTDFILL97_576 VDD VSS sg13g2_FILL8
XSTDFILL97_584 VDD VSS sg13g2_FILL8
XSTDFILL97_592 VDD VSS sg13g2_FILL8
XSTDFILL97_600 VDD VSS sg13g2_FILL8
XSTDFILL97_608 VDD VSS sg13g2_FILL8
XSTDFILL97_616 VDD VSS sg13g2_FILL8
XSTDFILL97_624 VDD VSS sg13g2_FILL8
XSTDFILL97_632 VDD VSS sg13g2_FILL8
XSTDFILL97_640 VDD VSS sg13g2_FILL8
XSTDFILL97_648 VDD VSS sg13g2_FILL8
XSTDFILL97_656 VDD VSS sg13g2_FILL8
XSTDFILL97_664 VDD VSS sg13g2_FILL8
XSTDFILL97_672 VDD VSS sg13g2_FILL8
XSTDFILL97_680 VDD VSS sg13g2_FILL8
XSTDFILL97_688 VDD VSS sg13g2_FILL8
XSTDFILL97_696 VDD VSS sg13g2_FILL8
XSTDFILL97_704 VDD VSS sg13g2_FILL8
XSTDFILL97_712 VDD VSS sg13g2_FILL8
XSTDFILL97_720 VDD VSS sg13g2_FILL8
XSTDFILL97_728 VDD VSS sg13g2_FILL8
XSTDFILL97_736 VDD VSS sg13g2_FILL8
XSTDFILL97_744 VDD VSS sg13g2_FILL8
XSTDFILL97_752 VDD VSS sg13g2_FILL8
XSTDFILL97_760 VDD VSS sg13g2_FILL8
XSTDFILL97_768 VDD VSS sg13g2_FILL8
XSTDFILL97_776 VDD VSS sg13g2_FILL8
XSTDFILL97_784 VDD VSS sg13g2_FILL8
XSTDFILL97_792 VDD VSS sg13g2_FILL8
XSTDFILL97_800 VDD VSS sg13g2_FILL8
XSTDFILL97_808 VDD VSS sg13g2_FILL8
XSTDFILL97_816 VDD VSS sg13g2_FILL8
XSTDFILL97_824 VDD VSS sg13g2_FILL8
XSTDFILL97_832 VDD VSS sg13g2_FILL8
XSTDFILL97_840 VDD VSS sg13g2_FILL8
XSTDFILL97_848 VDD VSS sg13g2_FILL8
XSTDFILL97_856 VDD VSS sg13g2_FILL8
XSTDFILL97_864 VDD VSS sg13g2_FILL8
XSTDFILL97_872 VDD VSS sg13g2_FILL8
XSTDFILL97_880 VDD VSS sg13g2_FILL8
XSTDFILL97_888 VDD VSS sg13g2_FILL8
XSTDFILL97_896 VDD VSS sg13g2_FILL8
XSTDFILL97_904 VDD VSS sg13g2_FILL8
XSTDFILL97_912 VDD VSS sg13g2_FILL8
XSTDFILL97_920 VDD VSS sg13g2_FILL8
XSTDFILL97_928 VDD VSS sg13g2_FILL8
XSTDFILL97_936 VDD VSS sg13g2_FILL8
XSTDFILL97_944 VDD VSS sg13g2_FILL8
XSTDFILL97_952 VDD VSS sg13g2_FILL8
XSTDFILL97_960 VDD VSS sg13g2_FILL8
XSTDFILL97_968 VDD VSS sg13g2_FILL8
XSTDFILL97_976 VDD VSS sg13g2_FILL8
XSTDFILL97_984 VDD VSS sg13g2_FILL8
XSTDFILL97_992 VDD VSS sg13g2_FILL8
XSTDFILL97_1000 VDD VSS sg13g2_FILL8
XSTDFILL97_1008 VDD VSS sg13g2_FILL8
XSTDFILL97_1016 VDD VSS sg13g2_FILL8
XSTDFILL97_1024 VDD VSS sg13g2_FILL8
XSTDFILL97_1032 VDD VSS sg13g2_FILL8
XSTDFILL97_1040 VDD VSS sg13g2_FILL8
XSTDFILL97_1048 VDD VSS sg13g2_FILL8
XSTDFILL97_1056 VDD VSS sg13g2_FILL8
XSTDFILL97_1064 VDD VSS sg13g2_FILL8
XSTDFILL97_1072 VDD VSS sg13g2_FILL8
XSTDFILL97_1080 VDD VSS sg13g2_FILL8
XSTDFILL97_1088 VDD VSS sg13g2_FILL8
XSTDFILL97_1096 VDD VSS sg13g2_FILL8
XSTDFILL97_1104 VDD VSS sg13g2_FILL8
XSTDFILL97_1112 VDD VSS sg13g2_FILL8
XSTDFILL97_1120 VDD VSS sg13g2_FILL8
XSTDFILL97_1128 VDD VSS sg13g2_FILL8
XSTDFILL97_1136 VDD VSS sg13g2_FILL8
XSTDFILL97_1144 VDD VSS sg13g2_FILL8
XSTDFILL97_1152 VDD VSS sg13g2_FILL8
XSTDFILL97_1160 VDD VSS sg13g2_FILL8
XSTDFILL97_1168 VDD VSS sg13g2_FILL8
XSTDFILL97_1176 VDD VSS sg13g2_FILL8
XSTDFILL97_1184 VDD VSS sg13g2_FILL8
XSTDFILL97_1192 VDD VSS sg13g2_FILL8
XSTDFILL97_1200 VDD VSS sg13g2_FILL8
XSTDFILL97_1208 VDD VSS sg13g2_FILL8
XSTDFILL97_1216 VDD VSS sg13g2_FILL8
XSTDFILL97_1224 VDD VSS sg13g2_FILL8
XSTDFILL97_1232 VDD VSS sg13g2_FILL8
XSTDFILL97_1240 VDD VSS sg13g2_FILL8
XSTDFILL97_1248 VDD VSS sg13g2_FILL8
XSTDFILL97_1256 VDD VSS sg13g2_FILL8
XSTDFILL97_1264 VDD VSS sg13g2_FILL8
XSTDFILL97_1272 VDD VSS sg13g2_FILL8
XSTDFILL97_1280 VDD VSS sg13g2_FILL8
XSTDFILL97_1288 VDD VSS sg13g2_FILL8
XSTDFILL97_1296 VDD VSS sg13g2_FILL8
XSTDFILL97_1304 VDD VSS sg13g2_FILL8
XSTDFILL97_1312 VDD VSS sg13g2_FILL8
XSTDFILL97_1320 VDD VSS sg13g2_FILL8
XSTDFILL97_1328 VDD VSS sg13g2_FILL8
XSTDFILL97_1336 VDD VSS sg13g2_FILL8
XSTDFILL97_1344 VDD VSS sg13g2_FILL8
XSTDFILL97_1352 VDD VSS sg13g2_FILL8
XSTDFILL97_1360 VDD VSS sg13g2_FILL8
XSTDFILL97_1368 VDD VSS sg13g2_FILL8
XSTDFILL97_1376 VDD VSS sg13g2_FILL8
XSTDFILL97_1384 VDD VSS sg13g2_FILL8
XSTDFILL97_1392 VDD VSS sg13g2_FILL8
XSTDFILL97_1400 VDD VSS sg13g2_FILL8
XSTDFILL97_1408 VDD VSS sg13g2_FILL8
XSTDFILL97_1416 VDD VSS sg13g2_FILL8
XSTDFILL97_1424 VDD VSS sg13g2_FILL8
XSTDFILL97_1432 VDD VSS sg13g2_FILL8
XSTDFILL97_1440 VDD VSS sg13g2_FILL8
XSTDFILL97_1448 VDD VSS sg13g2_FILL8
XSTDFILL97_1456 VDD VSS sg13g2_FILL8
XSTDFILL97_1464 VDD VSS sg13g2_FILL8
XSTDFILL97_1472 VDD VSS sg13g2_FILL8
XSTDFILL97_1480 VDD VSS sg13g2_FILL8
XSTDFILL97_1488 VDD VSS sg13g2_FILL8
XSTDFILL97_1496 VDD VSS sg13g2_FILL8
XSTDFILL97_1504 VDD VSS sg13g2_FILL8
XSTDFILL97_1512 VDD VSS sg13g2_FILL8
XSTDFILL97_1520 VDD VSS sg13g2_FILL8
XSTDFILL97_1528 VDD VSS sg13g2_FILL8
XSTDFILL97_1536 VDD VSS sg13g2_FILL8
XSTDFILL97_1544 VDD VSS sg13g2_FILL8
XSTDFILL97_1552 VDD VSS sg13g2_FILL8
XSTDFILL97_1560 VDD VSS sg13g2_FILL8
XSTDFILL97_1568 VDD VSS sg13g2_FILL8
XSTDFILL97_1576 VDD VSS sg13g2_FILL8
XSTDFILL97_1584 VDD VSS sg13g2_FILL8
XSTDFILL97_1592 VDD VSS sg13g2_FILL8
XSTDFILL97_1600 VDD VSS sg13g2_FILL8
XSTDFILL97_1608 VDD VSS sg13g2_FILL8
XSTDFILL97_1616 VDD VSS sg13g2_FILL8
XSTDFILL97_1624 VDD VSS sg13g2_FILL8
XSTDFILL97_1632 VDD VSS sg13g2_FILL8
XSTDFILL97_1640 VDD VSS sg13g2_FILL8
XSTDFILL97_1648 VDD VSS sg13g2_FILL8
XSTDFILL97_1656 VDD VSS sg13g2_FILL8
XSTDFILL97_1664 VDD VSS sg13g2_FILL8
XSTDFILL97_1672 VDD VSS sg13g2_FILL8
XSTDFILL97_1680 VDD VSS sg13g2_FILL8
XSTDFILL97_1688 VDD VSS sg13g2_FILL8
XSTDFILL97_1696 VDD VSS sg13g2_FILL8
XSTDFILL97_1704 VDD VSS sg13g2_FILL8
XSTDFILL97_1712 VDD VSS sg13g2_FILL8
XSTDFILL97_1720 VDD VSS sg13g2_FILL8
XSTDFILL97_1728 VDD VSS sg13g2_FILL8
XSTDFILL97_1736 VDD VSS sg13g2_FILL8
XSTDFILL97_1744 VDD VSS sg13g2_FILL8
XSTDFILL97_1752 VDD VSS sg13g2_FILL8
XSTDFILL97_1760 VDD VSS sg13g2_FILL8
XSTDFILL97_1768 VDD VSS sg13g2_FILL8
XSTDFILL97_1776 VDD VSS sg13g2_FILL8
XSTDFILL97_1784 VDD VSS sg13g2_FILL8
XSTDFILL97_1792 VDD VSS sg13g2_FILL8
XSTDFILL97_1800 VDD VSS sg13g2_FILL8
XSTDFILL97_1808 VDD VSS sg13g2_FILL8
XSTDFILL97_1816 VDD VSS sg13g2_FILL8
XSTDFILL97_1824 VDD VSS sg13g2_FILL8
XSTDFILL97_1832 VDD VSS sg13g2_FILL8
XSTDFILL97_1840 VDD VSS sg13g2_FILL8
XSTDFILL97_1848 VDD VSS sg13g2_FILL8
XSTDFILL97_1856 VDD VSS sg13g2_FILL8
XSTDFILL97_1864 VDD VSS sg13g2_FILL8
XSTDFILL97_1872 VDD VSS sg13g2_FILL8
XSTDFILL97_1880 VDD VSS sg13g2_FILL8
XSTDFILL97_1888 VDD VSS sg13g2_FILL8
XSTDFILL97_1896 VDD VSS sg13g2_FILL8
XSTDFILL97_1904 VDD VSS sg13g2_FILL8
XSTDFILL97_1912 VDD VSS sg13g2_FILL8
XSTDFILL97_1920 VDD VSS sg13g2_FILL8
XSTDFILL97_1928 VDD VSS sg13g2_FILL8
XSTDFILL97_1936 VDD VSS sg13g2_FILL8
XSTDFILL97_1944 VDD VSS sg13g2_FILL8
XSTDFILL97_1952 VDD VSS sg13g2_FILL8
XSTDFILL97_1960 VDD VSS sg13g2_FILL8
XSTDFILL97_1968 VDD VSS sg13g2_FILL8
XSTDFILL97_1976 VDD VSS sg13g2_FILL8
XSTDFILL97_1984 VDD VSS sg13g2_FILL8
XSTDFILL97_1992 VDD VSS sg13g2_FILL8
XSTDFILL97_2000 VDD VSS sg13g2_FILL8
XSTDFILL97_2008 VDD VSS sg13g2_FILL8
XSTDFILL97_2016 VDD VSS sg13g2_FILL8
XSTDFILL97_2024 VDD VSS sg13g2_FILL8
XSTDFILL97_2032 VDD VSS sg13g2_FILL8
XSTDFILL97_2040 VDD VSS sg13g2_FILL8
XSTDFILL97_2048 VDD VSS sg13g2_FILL8
XSTDFILL97_2056 VDD VSS sg13g2_FILL8
XSTDFILL97_2064 VDD VSS sg13g2_FILL8
XSTDFILL97_2072 VDD VSS sg13g2_FILL8
XSTDFILL97_2080 VDD VSS sg13g2_FILL8
XSTDFILL97_2088 VDD VSS sg13g2_FILL8
XSTDFILL97_2096 VDD VSS sg13g2_FILL8
XSTDFILL97_2104 VDD VSS sg13g2_FILL8
XSTDFILL97_2112 VDD VSS sg13g2_FILL8
XSTDFILL97_2120 VDD VSS sg13g2_FILL8
XSTDFILL97_2128 VDD VSS sg13g2_FILL8
XSTDFILL97_2136 VDD VSS sg13g2_FILL8
XSTDFILL97_2144 VDD VSS sg13g2_FILL8
XSTDFILL97_2152 VDD VSS sg13g2_FILL2
XSTDFILL98_0 VDD VSS sg13g2_FILL8
XSTDFILL98_8 VDD VSS sg13g2_FILL8
XSTDFILL98_16 VDD VSS sg13g2_FILL8
XSTDFILL98_24 VDD VSS sg13g2_FILL8
XSTDFILL98_32 VDD VSS sg13g2_FILL8
XSTDFILL98_40 VDD VSS sg13g2_FILL8
XSTDFILL98_48 VDD VSS sg13g2_FILL8
XSTDFILL98_56 VDD VSS sg13g2_FILL8
XSTDFILL98_64 VDD VSS sg13g2_FILL8
XSTDFILL98_72 VDD VSS sg13g2_FILL8
XSTDFILL98_80 VDD VSS sg13g2_FILL8
XSTDFILL98_88 VDD VSS sg13g2_FILL8
XSTDFILL98_96 VDD VSS sg13g2_FILL8
XSTDFILL98_104 VDD VSS sg13g2_FILL8
XSTDFILL98_112 VDD VSS sg13g2_FILL8
XSTDFILL98_120 VDD VSS sg13g2_FILL8
XSTDFILL98_128 VDD VSS sg13g2_FILL8
XSTDFILL98_136 VDD VSS sg13g2_FILL8
XSTDFILL98_144 VDD VSS sg13g2_FILL8
XSTDFILL98_152 VDD VSS sg13g2_FILL8
XSTDFILL98_160 VDD VSS sg13g2_FILL8
XSTDFILL98_168 VDD VSS sg13g2_FILL8
XSTDFILL98_176 VDD VSS sg13g2_FILL8
XSTDFILL98_184 VDD VSS sg13g2_FILL8
XSTDFILL98_192 VDD VSS sg13g2_FILL8
XSTDFILL98_200 VDD VSS sg13g2_FILL8
XSTDFILL98_208 VDD VSS sg13g2_FILL8
XSTDFILL98_216 VDD VSS sg13g2_FILL8
XSTDFILL98_224 VDD VSS sg13g2_FILL8
XSTDFILL98_232 VDD VSS sg13g2_FILL8
XSTDFILL98_240 VDD VSS sg13g2_FILL8
XSTDFILL98_248 VDD VSS sg13g2_FILL8
XSTDFILL98_256 VDD VSS sg13g2_FILL8
XSTDFILL98_264 VDD VSS sg13g2_FILL8
XSTDFILL98_272 VDD VSS sg13g2_FILL8
XSTDFILL98_280 VDD VSS sg13g2_FILL8
XSTDFILL98_288 VDD VSS sg13g2_FILL8
XSTDFILL98_296 VDD VSS sg13g2_FILL8
XSTDFILL98_304 VDD VSS sg13g2_FILL8
XSTDFILL98_312 VDD VSS sg13g2_FILL8
XSTDFILL98_320 VDD VSS sg13g2_FILL8
XSTDFILL98_328 VDD VSS sg13g2_FILL8
XSTDFILL98_336 VDD VSS sg13g2_FILL8
XSTDFILL98_344 VDD VSS sg13g2_FILL8
XSTDFILL98_352 VDD VSS sg13g2_FILL8
XSTDFILL98_360 VDD VSS sg13g2_FILL8
XSTDFILL98_368 VDD VSS sg13g2_FILL8
XSTDFILL98_376 VDD VSS sg13g2_FILL8
XSTDFILL98_384 VDD VSS sg13g2_FILL8
XSTDFILL98_392 VDD VSS sg13g2_FILL8
XSTDFILL98_400 VDD VSS sg13g2_FILL8
XSTDFILL98_408 VDD VSS sg13g2_FILL8
XSTDFILL98_416 VDD VSS sg13g2_FILL8
XSTDFILL98_424 VDD VSS sg13g2_FILL8
XSTDFILL98_432 VDD VSS sg13g2_FILL8
XSTDFILL98_440 VDD VSS sg13g2_FILL8
XSTDFILL98_448 VDD VSS sg13g2_FILL8
XSTDFILL98_456 VDD VSS sg13g2_FILL8
XSTDFILL98_464 VDD VSS sg13g2_FILL8
XSTDFILL98_472 VDD VSS sg13g2_FILL8
XSTDFILL98_480 VDD VSS sg13g2_FILL8
XSTDFILL98_488 VDD VSS sg13g2_FILL8
XSTDFILL98_496 VDD VSS sg13g2_FILL8
XSTDFILL98_504 VDD VSS sg13g2_FILL8
XSTDFILL98_512 VDD VSS sg13g2_FILL8
XSTDFILL98_520 VDD VSS sg13g2_FILL8
XSTDFILL98_528 VDD VSS sg13g2_FILL8
XSTDFILL98_536 VDD VSS sg13g2_FILL8
XSTDFILL98_544 VDD VSS sg13g2_FILL8
XSTDFILL98_552 VDD VSS sg13g2_FILL8
XSTDFILL98_560 VDD VSS sg13g2_FILL8
XSTDFILL98_568 VDD VSS sg13g2_FILL8
XSTDFILL98_576 VDD VSS sg13g2_FILL8
XSTDFILL98_584 VDD VSS sg13g2_FILL8
XSTDFILL98_592 VDD VSS sg13g2_FILL8
XSTDFILL98_600 VDD VSS sg13g2_FILL8
XSTDFILL98_608 VDD VSS sg13g2_FILL8
XSTDFILL98_616 VDD VSS sg13g2_FILL8
XSTDFILL98_624 VDD VSS sg13g2_FILL8
XSTDFILL98_632 VDD VSS sg13g2_FILL8
XSTDFILL98_640 VDD VSS sg13g2_FILL8
XSTDFILL98_648 VDD VSS sg13g2_FILL8
XSTDFILL98_656 VDD VSS sg13g2_FILL8
XSTDFILL98_664 VDD VSS sg13g2_FILL8
XSTDFILL98_672 VDD VSS sg13g2_FILL8
XSTDFILL98_680 VDD VSS sg13g2_FILL8
XSTDFILL98_688 VDD VSS sg13g2_FILL8
XSTDFILL98_696 VDD VSS sg13g2_FILL8
XSTDFILL98_704 VDD VSS sg13g2_FILL8
XSTDFILL98_712 VDD VSS sg13g2_FILL8
XSTDFILL98_720 VDD VSS sg13g2_FILL8
XSTDFILL98_728 VDD VSS sg13g2_FILL8
XSTDFILL98_736 VDD VSS sg13g2_FILL8
XSTDFILL98_744 VDD VSS sg13g2_FILL8
XSTDFILL98_752 VDD VSS sg13g2_FILL8
XSTDFILL98_760 VDD VSS sg13g2_FILL8
XSTDFILL98_768 VDD VSS sg13g2_FILL8
XSTDFILL98_776 VDD VSS sg13g2_FILL8
XSTDFILL98_784 VDD VSS sg13g2_FILL8
XSTDFILL98_792 VDD VSS sg13g2_FILL8
XSTDFILL98_800 VDD VSS sg13g2_FILL8
XSTDFILL98_808 VDD VSS sg13g2_FILL8
XSTDFILL98_816 VDD VSS sg13g2_FILL8
XSTDFILL98_824 VDD VSS sg13g2_FILL8
XSTDFILL98_832 VDD VSS sg13g2_FILL8
XSTDFILL98_840 VDD VSS sg13g2_FILL8
XSTDFILL98_848 VDD VSS sg13g2_FILL8
XSTDFILL98_856 VDD VSS sg13g2_FILL8
XSTDFILL98_864 VDD VSS sg13g2_FILL8
XSTDFILL98_872 VDD VSS sg13g2_FILL8
XSTDFILL98_880 VDD VSS sg13g2_FILL8
XSTDFILL98_888 VDD VSS sg13g2_FILL8
XSTDFILL98_896 VDD VSS sg13g2_FILL8
XSTDFILL98_904 VDD VSS sg13g2_FILL8
XSTDFILL98_912 VDD VSS sg13g2_FILL8
XSTDFILL98_920 VDD VSS sg13g2_FILL8
XSTDFILL98_928 VDD VSS sg13g2_FILL8
XSTDFILL98_936 VDD VSS sg13g2_FILL8
XSTDFILL98_944 VDD VSS sg13g2_FILL8
XSTDFILL98_952 VDD VSS sg13g2_FILL8
XSTDFILL98_960 VDD VSS sg13g2_FILL8
XSTDFILL98_968 VDD VSS sg13g2_FILL8
XSTDFILL98_976 VDD VSS sg13g2_FILL8
XSTDFILL98_984 VDD VSS sg13g2_FILL8
XSTDFILL98_992 VDD VSS sg13g2_FILL8
XSTDFILL98_1000 VDD VSS sg13g2_FILL8
XSTDFILL98_1008 VDD VSS sg13g2_FILL8
XSTDFILL98_1016 VDD VSS sg13g2_FILL8
XSTDFILL98_1024 VDD VSS sg13g2_FILL8
XSTDFILL98_1032 VDD VSS sg13g2_FILL8
XSTDFILL98_1040 VDD VSS sg13g2_FILL8
XSTDFILL98_1048 VDD VSS sg13g2_FILL8
XSTDFILL98_1056 VDD VSS sg13g2_FILL8
XSTDFILL98_1064 VDD VSS sg13g2_FILL8
XSTDFILL98_1072 VDD VSS sg13g2_FILL8
XSTDFILL98_1080 VDD VSS sg13g2_FILL8
XSTDFILL98_1088 VDD VSS sg13g2_FILL8
XSTDFILL98_1096 VDD VSS sg13g2_FILL8
XSTDFILL98_1104 VDD VSS sg13g2_FILL8
XSTDFILL98_1112 VDD VSS sg13g2_FILL8
XSTDFILL98_1120 VDD VSS sg13g2_FILL8
XSTDFILL98_1128 VDD VSS sg13g2_FILL8
XSTDFILL98_1136 VDD VSS sg13g2_FILL8
XSTDFILL98_1144 VDD VSS sg13g2_FILL8
XSTDFILL98_1152 VDD VSS sg13g2_FILL8
XSTDFILL98_1160 VDD VSS sg13g2_FILL8
XSTDFILL98_1168 VDD VSS sg13g2_FILL8
XSTDFILL98_1176 VDD VSS sg13g2_FILL8
XSTDFILL98_1184 VDD VSS sg13g2_FILL8
XSTDFILL98_1192 VDD VSS sg13g2_FILL8
XSTDFILL98_1200 VDD VSS sg13g2_FILL8
XSTDFILL98_1208 VDD VSS sg13g2_FILL8
XSTDFILL98_1216 VDD VSS sg13g2_FILL8
XSTDFILL98_1224 VDD VSS sg13g2_FILL8
XSTDFILL98_1232 VDD VSS sg13g2_FILL8
XSTDFILL98_1240 VDD VSS sg13g2_FILL8
XSTDFILL98_1248 VDD VSS sg13g2_FILL8
XSTDFILL98_1256 VDD VSS sg13g2_FILL8
XSTDFILL98_1264 VDD VSS sg13g2_FILL8
XSTDFILL98_1272 VDD VSS sg13g2_FILL8
XSTDFILL98_1280 VDD VSS sg13g2_FILL8
XSTDFILL98_1288 VDD VSS sg13g2_FILL8
XSTDFILL98_1296 VDD VSS sg13g2_FILL8
XSTDFILL98_1304 VDD VSS sg13g2_FILL8
XSTDFILL98_1312 VDD VSS sg13g2_FILL8
XSTDFILL98_1320 VDD VSS sg13g2_FILL8
XSTDFILL98_1328 VDD VSS sg13g2_FILL8
XSTDFILL98_1336 VDD VSS sg13g2_FILL8
XSTDFILL98_1344 VDD VSS sg13g2_FILL8
XSTDFILL98_1352 VDD VSS sg13g2_FILL8
XSTDFILL98_1360 VDD VSS sg13g2_FILL8
XSTDFILL98_1368 VDD VSS sg13g2_FILL8
XSTDFILL98_1376 VDD VSS sg13g2_FILL8
XSTDFILL98_1384 VDD VSS sg13g2_FILL8
XSTDFILL98_1392 VDD VSS sg13g2_FILL8
XSTDFILL98_1400 VDD VSS sg13g2_FILL8
XSTDFILL98_1408 VDD VSS sg13g2_FILL8
XSTDFILL98_1416 VDD VSS sg13g2_FILL8
XSTDFILL98_1424 VDD VSS sg13g2_FILL8
XSTDFILL98_1432 VDD VSS sg13g2_FILL8
XSTDFILL98_1440 VDD VSS sg13g2_FILL8
XSTDFILL98_1448 VDD VSS sg13g2_FILL8
XSTDFILL98_1456 VDD VSS sg13g2_FILL8
XSTDFILL98_1464 VDD VSS sg13g2_FILL8
XSTDFILL98_1472 VDD VSS sg13g2_FILL8
XSTDFILL98_1480 VDD VSS sg13g2_FILL8
XSTDFILL98_1488 VDD VSS sg13g2_FILL8
XSTDFILL98_1496 VDD VSS sg13g2_FILL8
XSTDFILL98_1504 VDD VSS sg13g2_FILL8
XSTDFILL98_1512 VDD VSS sg13g2_FILL8
XSTDFILL98_1520 VDD VSS sg13g2_FILL8
XSTDFILL98_1528 VDD VSS sg13g2_FILL8
XSTDFILL98_1536 VDD VSS sg13g2_FILL8
XSTDFILL98_1544 VDD VSS sg13g2_FILL8
XSTDFILL98_1552 VDD VSS sg13g2_FILL8
XSTDFILL98_1560 VDD VSS sg13g2_FILL8
XSTDFILL98_1568 VDD VSS sg13g2_FILL8
XSTDFILL98_1576 VDD VSS sg13g2_FILL8
XSTDFILL98_1584 VDD VSS sg13g2_FILL8
XSTDFILL98_1592 VDD VSS sg13g2_FILL8
XSTDFILL98_1600 VDD VSS sg13g2_FILL8
XSTDFILL98_1608 VDD VSS sg13g2_FILL8
XSTDFILL98_1616 VDD VSS sg13g2_FILL8
XSTDFILL98_1624 VDD VSS sg13g2_FILL8
XSTDFILL98_1632 VDD VSS sg13g2_FILL8
XSTDFILL98_1640 VDD VSS sg13g2_FILL8
XSTDFILL98_1648 VDD VSS sg13g2_FILL8
XSTDFILL98_1656 VDD VSS sg13g2_FILL8
XSTDFILL98_1664 VDD VSS sg13g2_FILL8
XSTDFILL98_1672 VDD VSS sg13g2_FILL8
XSTDFILL98_1680 VDD VSS sg13g2_FILL8
XSTDFILL98_1688 VDD VSS sg13g2_FILL8
XSTDFILL98_1696 VDD VSS sg13g2_FILL8
XSTDFILL98_1704 VDD VSS sg13g2_FILL8
XSTDFILL98_1712 VDD VSS sg13g2_FILL8
XSTDFILL98_1720 VDD VSS sg13g2_FILL8
XSTDFILL98_1728 VDD VSS sg13g2_FILL8
XSTDFILL98_1736 VDD VSS sg13g2_FILL8
XSTDFILL98_1744 VDD VSS sg13g2_FILL8
XSTDFILL98_1752 VDD VSS sg13g2_FILL8
XSTDFILL98_1760 VDD VSS sg13g2_FILL8
XSTDFILL98_1768 VDD VSS sg13g2_FILL8
XSTDFILL98_1776 VDD VSS sg13g2_FILL8
XSTDFILL98_1784 VDD VSS sg13g2_FILL8
XSTDFILL98_1792 VDD VSS sg13g2_FILL8
XSTDFILL98_1800 VDD VSS sg13g2_FILL8
XSTDFILL98_1808 VDD VSS sg13g2_FILL8
XSTDFILL98_1816 VDD VSS sg13g2_FILL8
XSTDFILL98_1824 VDD VSS sg13g2_FILL8
XSTDFILL98_1832 VDD VSS sg13g2_FILL8
XSTDFILL98_1840 VDD VSS sg13g2_FILL8
XSTDFILL98_1848 VDD VSS sg13g2_FILL8
XSTDFILL98_1856 VDD VSS sg13g2_FILL8
XSTDFILL98_1864 VDD VSS sg13g2_FILL8
XSTDFILL98_1872 VDD VSS sg13g2_FILL8
XSTDFILL98_1880 VDD VSS sg13g2_FILL8
XSTDFILL98_1888 VDD VSS sg13g2_FILL8
XSTDFILL98_1896 VDD VSS sg13g2_FILL8
XSTDFILL98_1904 VDD VSS sg13g2_FILL8
XSTDFILL98_1912 VDD VSS sg13g2_FILL8
XSTDFILL98_1920 VDD VSS sg13g2_FILL8
XSTDFILL98_1928 VDD VSS sg13g2_FILL8
XSTDFILL98_1936 VDD VSS sg13g2_FILL8
XSTDFILL98_1944 VDD VSS sg13g2_FILL8
XSTDFILL98_1952 VDD VSS sg13g2_FILL8
XSTDFILL98_1960 VDD VSS sg13g2_FILL8
XSTDFILL98_1968 VDD VSS sg13g2_FILL8
XSTDFILL98_1976 VDD VSS sg13g2_FILL8
XSTDFILL98_1984 VDD VSS sg13g2_FILL8
XSTDFILL98_1992 VDD VSS sg13g2_FILL8
XSTDFILL98_2000 VDD VSS sg13g2_FILL8
XSTDFILL98_2008 VDD VSS sg13g2_FILL8
XSTDFILL98_2016 VDD VSS sg13g2_FILL8
XSTDFILL98_2024 VDD VSS sg13g2_FILL8
XSTDFILL98_2032 VDD VSS sg13g2_FILL8
XSTDFILL98_2040 VDD VSS sg13g2_FILL8
XSTDFILL98_2048 VDD VSS sg13g2_FILL8
XSTDFILL98_2056 VDD VSS sg13g2_FILL8
XSTDFILL98_2064 VDD VSS sg13g2_FILL8
XSTDFILL98_2072 VDD VSS sg13g2_FILL8
XSTDFILL98_2080 VDD VSS sg13g2_FILL8
XSTDFILL98_2088 VDD VSS sg13g2_FILL8
XSTDFILL98_2096 VDD VSS sg13g2_FILL8
XSTDFILL98_2104 VDD VSS sg13g2_FILL8
XSTDFILL98_2112 VDD VSS sg13g2_FILL8
XSTDFILL98_2120 VDD VSS sg13g2_FILL8
XSTDFILL98_2128 VDD VSS sg13g2_FILL8
XSTDFILL98_2136 VDD VSS sg13g2_FILL8
XSTDFILL98_2144 VDD VSS sg13g2_FILL8
XSTDFILL98_2152 VDD VSS sg13g2_FILL2
XSTDFILL99_0 VDD VSS sg13g2_FILL8
XSTDFILL99_8 VDD VSS sg13g2_FILL8
XSTDFILL99_16 VDD VSS sg13g2_FILL8
XSTDFILL99_24 VDD VSS sg13g2_FILL8
XSTDFILL99_32 VDD VSS sg13g2_FILL8
XSTDFILL99_40 VDD VSS sg13g2_FILL8
XSTDFILL99_48 VDD VSS sg13g2_FILL8
XSTDFILL99_56 VDD VSS sg13g2_FILL8
XSTDFILL99_64 VDD VSS sg13g2_FILL8
XSTDFILL99_72 VDD VSS sg13g2_FILL8
XSTDFILL99_80 VDD VSS sg13g2_FILL8
XSTDFILL99_88 VDD VSS sg13g2_FILL8
XSTDFILL99_96 VDD VSS sg13g2_FILL8
XSTDFILL99_104 VDD VSS sg13g2_FILL8
XSTDFILL99_112 VDD VSS sg13g2_FILL8
XSTDFILL99_120 VDD VSS sg13g2_FILL8
XSTDFILL99_128 VDD VSS sg13g2_FILL8
XSTDFILL99_136 VDD VSS sg13g2_FILL8
XSTDFILL99_144 VDD VSS sg13g2_FILL8
XSTDFILL99_152 VDD VSS sg13g2_FILL8
XSTDFILL99_160 VDD VSS sg13g2_FILL8
XSTDFILL99_168 VDD VSS sg13g2_FILL8
XSTDFILL99_176 VDD VSS sg13g2_FILL8
XSTDFILL99_184 VDD VSS sg13g2_FILL8
XSTDFILL99_192 VDD VSS sg13g2_FILL8
XSTDFILL99_200 VDD VSS sg13g2_FILL8
XSTDFILL99_208 VDD VSS sg13g2_FILL8
XSTDFILL99_216 VDD VSS sg13g2_FILL8
XSTDFILL99_224 VDD VSS sg13g2_FILL8
XSTDFILL99_232 VDD VSS sg13g2_FILL8
XSTDFILL99_240 VDD VSS sg13g2_FILL8
XSTDFILL99_248 VDD VSS sg13g2_FILL8
XSTDFILL99_256 VDD VSS sg13g2_FILL8
XSTDFILL99_264 VDD VSS sg13g2_FILL8
XSTDFILL99_272 VDD VSS sg13g2_FILL8
XSTDFILL99_280 VDD VSS sg13g2_FILL8
XSTDFILL99_288 VDD VSS sg13g2_FILL8
XSTDFILL99_296 VDD VSS sg13g2_FILL8
XSTDFILL99_304 VDD VSS sg13g2_FILL8
XSTDFILL99_312 VDD VSS sg13g2_FILL8
XSTDFILL99_320 VDD VSS sg13g2_FILL8
XSTDFILL99_328 VDD VSS sg13g2_FILL8
XSTDFILL99_336 VDD VSS sg13g2_FILL8
XSTDFILL99_344 VDD VSS sg13g2_FILL8
XSTDFILL99_352 VDD VSS sg13g2_FILL8
XSTDFILL99_360 VDD VSS sg13g2_FILL8
XSTDFILL99_368 VDD VSS sg13g2_FILL8
XSTDFILL99_376 VDD VSS sg13g2_FILL8
XSTDFILL99_384 VDD VSS sg13g2_FILL8
XSTDFILL99_392 VDD VSS sg13g2_FILL8
XSTDFILL99_400 VDD VSS sg13g2_FILL8
XSTDFILL99_408 VDD VSS sg13g2_FILL8
XSTDFILL99_416 VDD VSS sg13g2_FILL8
XSTDFILL99_424 VDD VSS sg13g2_FILL8
XSTDFILL99_432 VDD VSS sg13g2_FILL8
XSTDFILL99_440 VDD VSS sg13g2_FILL8
XSTDFILL99_448 VDD VSS sg13g2_FILL8
XSTDFILL99_456 VDD VSS sg13g2_FILL8
XSTDFILL99_464 VDD VSS sg13g2_FILL8
XSTDFILL99_472 VDD VSS sg13g2_FILL8
XSTDFILL99_480 VDD VSS sg13g2_FILL8
XSTDFILL99_488 VDD VSS sg13g2_FILL8
XSTDFILL99_496 VDD VSS sg13g2_FILL8
XSTDFILL99_504 VDD VSS sg13g2_FILL8
XSTDFILL99_512 VDD VSS sg13g2_FILL8
XSTDFILL99_520 VDD VSS sg13g2_FILL8
XSTDFILL99_528 VDD VSS sg13g2_FILL8
XSTDFILL99_536 VDD VSS sg13g2_FILL8
XSTDFILL99_544 VDD VSS sg13g2_FILL8
XSTDFILL99_552 VDD VSS sg13g2_FILL8
XSTDFILL99_560 VDD VSS sg13g2_FILL8
XSTDFILL99_568 VDD VSS sg13g2_FILL8
XSTDFILL99_576 VDD VSS sg13g2_FILL8
XSTDFILL99_584 VDD VSS sg13g2_FILL8
XSTDFILL99_592 VDD VSS sg13g2_FILL8
XSTDFILL99_600 VDD VSS sg13g2_FILL8
XSTDFILL99_608 VDD VSS sg13g2_FILL8
XSTDFILL99_616 VDD VSS sg13g2_FILL8
XSTDFILL99_624 VDD VSS sg13g2_FILL8
XSTDFILL99_632 VDD VSS sg13g2_FILL8
XSTDFILL99_640 VDD VSS sg13g2_FILL8
XSTDFILL99_648 VDD VSS sg13g2_FILL8
XSTDFILL99_656 VDD VSS sg13g2_FILL8
XSTDFILL99_664 VDD VSS sg13g2_FILL8
XSTDFILL99_672 VDD VSS sg13g2_FILL8
XSTDFILL99_680 VDD VSS sg13g2_FILL8
XSTDFILL99_688 VDD VSS sg13g2_FILL8
XSTDFILL99_696 VDD VSS sg13g2_FILL8
XSTDFILL99_704 VDD VSS sg13g2_FILL8
XSTDFILL99_712 VDD VSS sg13g2_FILL8
XSTDFILL99_720 VDD VSS sg13g2_FILL8
XSTDFILL99_728 VDD VSS sg13g2_FILL8
XSTDFILL99_736 VDD VSS sg13g2_FILL8
XSTDFILL99_744 VDD VSS sg13g2_FILL8
XSTDFILL99_752 VDD VSS sg13g2_FILL8
XSTDFILL99_760 VDD VSS sg13g2_FILL8
XSTDFILL99_768 VDD VSS sg13g2_FILL8
XSTDFILL99_776 VDD VSS sg13g2_FILL8
XSTDFILL99_784 VDD VSS sg13g2_FILL8
XSTDFILL99_792 VDD VSS sg13g2_FILL8
XSTDFILL99_800 VDD VSS sg13g2_FILL8
XSTDFILL99_808 VDD VSS sg13g2_FILL8
XSTDFILL99_816 VDD VSS sg13g2_FILL8
XSTDFILL99_824 VDD VSS sg13g2_FILL8
XSTDFILL99_832 VDD VSS sg13g2_FILL8
XSTDFILL99_840 VDD VSS sg13g2_FILL8
XSTDFILL99_848 VDD VSS sg13g2_FILL8
XSTDFILL99_856 VDD VSS sg13g2_FILL8
XSTDFILL99_864 VDD VSS sg13g2_FILL8
XSTDFILL99_872 VDD VSS sg13g2_FILL8
XSTDFILL99_880 VDD VSS sg13g2_FILL8
XSTDFILL99_888 VDD VSS sg13g2_FILL8
XSTDFILL99_896 VDD VSS sg13g2_FILL8
XSTDFILL99_904 VDD VSS sg13g2_FILL8
XSTDFILL99_912 VDD VSS sg13g2_FILL8
XSTDFILL99_920 VDD VSS sg13g2_FILL8
XSTDFILL99_928 VDD VSS sg13g2_FILL8
XSTDFILL99_936 VDD VSS sg13g2_FILL8
XSTDFILL99_944 VDD VSS sg13g2_FILL8
XSTDFILL99_952 VDD VSS sg13g2_FILL8
XSTDFILL99_960 VDD VSS sg13g2_FILL8
XSTDFILL99_968 VDD VSS sg13g2_FILL8
XSTDFILL99_976 VDD VSS sg13g2_FILL8
XSTDFILL99_984 VDD VSS sg13g2_FILL8
XSTDFILL99_992 VDD VSS sg13g2_FILL8
XSTDFILL99_1000 VDD VSS sg13g2_FILL8
XSTDFILL99_1008 VDD VSS sg13g2_FILL8
XSTDFILL99_1016 VDD VSS sg13g2_FILL8
XSTDFILL99_1024 VDD VSS sg13g2_FILL8
XSTDFILL99_1032 VDD VSS sg13g2_FILL8
XSTDFILL99_1040 VDD VSS sg13g2_FILL8
XSTDFILL99_1048 VDD VSS sg13g2_FILL8
XSTDFILL99_1056 VDD VSS sg13g2_FILL8
XSTDFILL99_1064 VDD VSS sg13g2_FILL8
XSTDFILL99_1072 VDD VSS sg13g2_FILL8
XSTDFILL99_1080 VDD VSS sg13g2_FILL8
XSTDFILL99_1088 VDD VSS sg13g2_FILL8
XSTDFILL99_1096 VDD VSS sg13g2_FILL8
XSTDFILL99_1104 VDD VSS sg13g2_FILL8
XSTDFILL99_1112 VDD VSS sg13g2_FILL8
XSTDFILL99_1120 VDD VSS sg13g2_FILL8
XSTDFILL99_1128 VDD VSS sg13g2_FILL8
XSTDFILL99_1136 VDD VSS sg13g2_FILL8
XSTDFILL99_1144 VDD VSS sg13g2_FILL8
XSTDFILL99_1152 VDD VSS sg13g2_FILL8
XSTDFILL99_1160 VDD VSS sg13g2_FILL8
XSTDFILL99_1168 VDD VSS sg13g2_FILL8
XSTDFILL99_1176 VDD VSS sg13g2_FILL8
XSTDFILL99_1184 VDD VSS sg13g2_FILL8
XSTDFILL99_1192 VDD VSS sg13g2_FILL8
XSTDFILL99_1200 VDD VSS sg13g2_FILL8
XSTDFILL99_1208 VDD VSS sg13g2_FILL8
XSTDFILL99_1216 VDD VSS sg13g2_FILL8
XSTDFILL99_1224 VDD VSS sg13g2_FILL8
XSTDFILL99_1232 VDD VSS sg13g2_FILL8
XSTDFILL99_1240 VDD VSS sg13g2_FILL8
XSTDFILL99_1248 VDD VSS sg13g2_FILL8
XSTDFILL99_1256 VDD VSS sg13g2_FILL8
XSTDFILL99_1264 VDD VSS sg13g2_FILL8
XSTDFILL99_1272 VDD VSS sg13g2_FILL8
XSTDFILL99_1280 VDD VSS sg13g2_FILL8
XSTDFILL99_1288 VDD VSS sg13g2_FILL8
XSTDFILL99_1296 VDD VSS sg13g2_FILL8
XSTDFILL99_1304 VDD VSS sg13g2_FILL8
XSTDFILL99_1312 VDD VSS sg13g2_FILL8
XSTDFILL99_1320 VDD VSS sg13g2_FILL8
XSTDFILL99_1328 VDD VSS sg13g2_FILL8
XSTDFILL99_1336 VDD VSS sg13g2_FILL8
XSTDFILL99_1344 VDD VSS sg13g2_FILL8
XSTDFILL99_1352 VDD VSS sg13g2_FILL8
XSTDFILL99_1360 VDD VSS sg13g2_FILL8
XSTDFILL99_1368 VDD VSS sg13g2_FILL8
XSTDFILL99_1376 VDD VSS sg13g2_FILL8
XSTDFILL99_1384 VDD VSS sg13g2_FILL8
XSTDFILL99_1392 VDD VSS sg13g2_FILL8
XSTDFILL99_1400 VDD VSS sg13g2_FILL8
XSTDFILL99_1408 VDD VSS sg13g2_FILL8
XSTDFILL99_1416 VDD VSS sg13g2_FILL8
XSTDFILL99_1424 VDD VSS sg13g2_FILL8
XSTDFILL99_1432 VDD VSS sg13g2_FILL8
XSTDFILL99_1440 VDD VSS sg13g2_FILL8
XSTDFILL99_1448 VDD VSS sg13g2_FILL8
XSTDFILL99_1456 VDD VSS sg13g2_FILL8
XSTDFILL99_1464 VDD VSS sg13g2_FILL8
XSTDFILL99_1472 VDD VSS sg13g2_FILL8
XSTDFILL99_1480 VDD VSS sg13g2_FILL8
XSTDFILL99_1488 VDD VSS sg13g2_FILL8
XSTDFILL99_1496 VDD VSS sg13g2_FILL8
XSTDFILL99_1504 VDD VSS sg13g2_FILL8
XSTDFILL99_1512 VDD VSS sg13g2_FILL8
XSTDFILL99_1520 VDD VSS sg13g2_FILL8
XSTDFILL99_1528 VDD VSS sg13g2_FILL8
XSTDFILL99_1536 VDD VSS sg13g2_FILL8
XSTDFILL99_1544 VDD VSS sg13g2_FILL8
XSTDFILL99_1552 VDD VSS sg13g2_FILL8
XSTDFILL99_1560 VDD VSS sg13g2_FILL8
XSTDFILL99_1568 VDD VSS sg13g2_FILL8
XSTDFILL99_1576 VDD VSS sg13g2_FILL8
XSTDFILL99_1584 VDD VSS sg13g2_FILL8
XSTDFILL99_1592 VDD VSS sg13g2_FILL8
XSTDFILL99_1600 VDD VSS sg13g2_FILL8
XSTDFILL99_1608 VDD VSS sg13g2_FILL8
XSTDFILL99_1616 VDD VSS sg13g2_FILL8
XSTDFILL99_1624 VDD VSS sg13g2_FILL8
XSTDFILL99_1632 VDD VSS sg13g2_FILL8
XSTDFILL99_1640 VDD VSS sg13g2_FILL8
XSTDFILL99_1648 VDD VSS sg13g2_FILL8
XSTDFILL99_1656 VDD VSS sg13g2_FILL8
XSTDFILL99_1664 VDD VSS sg13g2_FILL8
XSTDFILL99_1672 VDD VSS sg13g2_FILL8
XSTDFILL99_1680 VDD VSS sg13g2_FILL8
XSTDFILL99_1688 VDD VSS sg13g2_FILL8
XSTDFILL99_1696 VDD VSS sg13g2_FILL8
XSTDFILL99_1704 VDD VSS sg13g2_FILL8
XSTDFILL99_1712 VDD VSS sg13g2_FILL8
XSTDFILL99_1720 VDD VSS sg13g2_FILL8
XSTDFILL99_1728 VDD VSS sg13g2_FILL8
XSTDFILL99_1736 VDD VSS sg13g2_FILL8
XSTDFILL99_1744 VDD VSS sg13g2_FILL8
XSTDFILL99_1752 VDD VSS sg13g2_FILL8
XSTDFILL99_1760 VDD VSS sg13g2_FILL8
XSTDFILL99_1768 VDD VSS sg13g2_FILL8
XSTDFILL99_1776 VDD VSS sg13g2_FILL8
XSTDFILL99_1784 VDD VSS sg13g2_FILL8
XSTDFILL99_1792 VDD VSS sg13g2_FILL8
XSTDFILL99_1800 VDD VSS sg13g2_FILL8
XSTDFILL99_1808 VDD VSS sg13g2_FILL8
XSTDFILL99_1816 VDD VSS sg13g2_FILL8
XSTDFILL99_1824 VDD VSS sg13g2_FILL8
XSTDFILL99_1832 VDD VSS sg13g2_FILL8
XSTDFILL99_1840 VDD VSS sg13g2_FILL8
XSTDFILL99_1848 VDD VSS sg13g2_FILL8
XSTDFILL99_1856 VDD VSS sg13g2_FILL8
XSTDFILL99_1864 VDD VSS sg13g2_FILL8
XSTDFILL99_1872 VDD VSS sg13g2_FILL8
XSTDFILL99_1880 VDD VSS sg13g2_FILL8
XSTDFILL99_1888 VDD VSS sg13g2_FILL8
XSTDFILL99_1896 VDD VSS sg13g2_FILL8
XSTDFILL99_1904 VDD VSS sg13g2_FILL8
XSTDFILL99_1912 VDD VSS sg13g2_FILL8
XSTDFILL99_1920 VDD VSS sg13g2_FILL8
XSTDFILL99_1928 VDD VSS sg13g2_FILL8
XSTDFILL99_1936 VDD VSS sg13g2_FILL8
XSTDFILL99_1944 VDD VSS sg13g2_FILL8
XSTDFILL99_1952 VDD VSS sg13g2_FILL8
XSTDFILL99_1960 VDD VSS sg13g2_FILL8
XSTDFILL99_1968 VDD VSS sg13g2_FILL8
XSTDFILL99_1976 VDD VSS sg13g2_FILL8
XSTDFILL99_1984 VDD VSS sg13g2_FILL8
XSTDFILL99_1992 VDD VSS sg13g2_FILL8
XSTDFILL99_2000 VDD VSS sg13g2_FILL8
XSTDFILL99_2008 VDD VSS sg13g2_FILL8
XSTDFILL99_2016 VDD VSS sg13g2_FILL8
XSTDFILL99_2024 VDD VSS sg13g2_FILL8
XSTDFILL99_2032 VDD VSS sg13g2_FILL8
XSTDFILL99_2040 VDD VSS sg13g2_FILL8
XSTDFILL99_2048 VDD VSS sg13g2_FILL8
XSTDFILL99_2056 VDD VSS sg13g2_FILL8
XSTDFILL99_2064 VDD VSS sg13g2_FILL8
XSTDFILL99_2072 VDD VSS sg13g2_FILL8
XSTDFILL99_2080 VDD VSS sg13g2_FILL8
XSTDFILL99_2088 VDD VSS sg13g2_FILL8
XSTDFILL99_2096 VDD VSS sg13g2_FILL8
XSTDFILL99_2104 VDD VSS sg13g2_FILL8
XSTDFILL99_2112 VDD VSS sg13g2_FILL8
XSTDFILL99_2120 VDD VSS sg13g2_FILL8
XSTDFILL99_2128 VDD VSS sg13g2_FILL8
XSTDFILL99_2136 VDD VSS sg13g2_FILL8
XSTDFILL99_2144 VDD VSS sg13g2_FILL8
XSTDFILL99_2152 VDD VSS sg13g2_FILL2
XSTDFILL101_0 VDD VSS sg13g2_FILL8
XSTDFILL101_8 VDD VSS sg13g2_FILL8
XSTDFILL101_16 VDD VSS sg13g2_FILL8
XSTDFILL101_24 VDD VSS sg13g2_FILL8
XSTDFILL101_32 VDD VSS sg13g2_FILL8
XSTDFILL101_40 VDD VSS sg13g2_FILL8
XSTDFILL101_48 VDD VSS sg13g2_FILL8
XSTDFILL101_56 VDD VSS sg13g2_FILL8
XSTDFILL101_64 VDD VSS sg13g2_FILL8
XSTDFILL101_72 VDD VSS sg13g2_FILL8
XSTDFILL101_80 VDD VSS sg13g2_FILL8
XSTDFILL101_88 VDD VSS sg13g2_FILL8
XSTDFILL101_96 VDD VSS sg13g2_FILL8
XSTDFILL101_104 VDD VSS sg13g2_FILL8
XSTDFILL101_112 VDD VSS sg13g2_FILL8
XSTDFILL101_120 VDD VSS sg13g2_FILL8
XSTDFILL101_128 VDD VSS sg13g2_FILL8
XSTDFILL101_136 VDD VSS sg13g2_FILL8
XSTDFILL101_144 VDD VSS sg13g2_FILL8
XSTDFILL101_152 VDD VSS sg13g2_FILL8
XSTDFILL101_160 VDD VSS sg13g2_FILL8
XSTDFILL101_168 VDD VSS sg13g2_FILL8
XSTDFILL101_176 VDD VSS sg13g2_FILL8
XSTDFILL101_184 VDD VSS sg13g2_FILL8
XSTDFILL101_192 VDD VSS sg13g2_FILL8
XSTDFILL101_200 VDD VSS sg13g2_FILL8
XSTDFILL101_208 VDD VSS sg13g2_FILL8
XSTDFILL101_216 VDD VSS sg13g2_FILL8
XSTDFILL101_224 VDD VSS sg13g2_FILL8
XSTDFILL101_232 VDD VSS sg13g2_FILL8
XSTDFILL101_240 VDD VSS sg13g2_FILL8
XSTDFILL101_248 VDD VSS sg13g2_FILL8
XSTDFILL101_256 VDD VSS sg13g2_FILL8
XSTDFILL101_264 VDD VSS sg13g2_FILL8
XSTDFILL101_272 VDD VSS sg13g2_FILL8
XSTDFILL101_280 VDD VSS sg13g2_FILL8
XSTDFILL101_288 VDD VSS sg13g2_FILL8
XSTDFILL101_296 VDD VSS sg13g2_FILL8
XSTDFILL101_304 VDD VSS sg13g2_FILL8
XSTDFILL101_312 VDD VSS sg13g2_FILL8
XSTDFILL101_320 VDD VSS sg13g2_FILL8
XSTDFILL101_328 VDD VSS sg13g2_FILL8
XSTDFILL101_336 VDD VSS sg13g2_FILL8
XSTDFILL101_344 VDD VSS sg13g2_FILL8
XSTDFILL101_352 VDD VSS sg13g2_FILL8
XSTDFILL101_360 VDD VSS sg13g2_FILL8
XSTDFILL101_368 VDD VSS sg13g2_FILL8
XSTDFILL101_376 VDD VSS sg13g2_FILL8
XSTDFILL101_384 VDD VSS sg13g2_FILL8
XSTDFILL101_392 VDD VSS sg13g2_FILL8
XSTDFILL101_400 VDD VSS sg13g2_FILL8
XSTDFILL101_408 VDD VSS sg13g2_FILL8
XSTDFILL101_416 VDD VSS sg13g2_FILL8
XSTDFILL101_424 VDD VSS sg13g2_FILL8
XSTDFILL101_432 VDD VSS sg13g2_FILL8
XSTDFILL101_440 VDD VSS sg13g2_FILL8
XSTDFILL101_448 VDD VSS sg13g2_FILL8
XSTDFILL101_456 VDD VSS sg13g2_FILL8
XSTDFILL101_464 VDD VSS sg13g2_FILL8
XSTDFILL101_472 VDD VSS sg13g2_FILL8
XSTDFILL101_480 VDD VSS sg13g2_FILL8
XSTDFILL101_488 VDD VSS sg13g2_FILL8
XSTDFILL101_496 VDD VSS sg13g2_FILL8
XSTDFILL101_504 VDD VSS sg13g2_FILL8
XSTDFILL101_512 VDD VSS sg13g2_FILL8
XSTDFILL101_520 VDD VSS sg13g2_FILL8
XSTDFILL101_528 VDD VSS sg13g2_FILL8
XSTDFILL101_536 VDD VSS sg13g2_FILL8
XSTDFILL101_544 VDD VSS sg13g2_FILL8
XSTDFILL101_552 VDD VSS sg13g2_FILL8
XSTDFILL101_560 VDD VSS sg13g2_FILL8
XSTDFILL101_568 VDD VSS sg13g2_FILL8
XSTDFILL101_576 VDD VSS sg13g2_FILL8
XSTDFILL101_584 VDD VSS sg13g2_FILL8
XSTDFILL101_592 VDD VSS sg13g2_FILL8
XSTDFILL101_600 VDD VSS sg13g2_FILL8
XSTDFILL101_608 VDD VSS sg13g2_FILL8
XSTDFILL101_616 VDD VSS sg13g2_FILL8
XSTDFILL101_624 VDD VSS sg13g2_FILL8
XSTDFILL101_632 VDD VSS sg13g2_FILL8
XSTDFILL101_640 VDD VSS sg13g2_FILL8
XSTDFILL101_648 VDD VSS sg13g2_FILL8
XSTDFILL101_656 VDD VSS sg13g2_FILL8
XSTDFILL101_664 VDD VSS sg13g2_FILL8
XSTDFILL101_672 VDD VSS sg13g2_FILL8
XSTDFILL101_680 VDD VSS sg13g2_FILL8
XSTDFILL101_688 VDD VSS sg13g2_FILL8
XSTDFILL101_696 VDD VSS sg13g2_FILL8
XSTDFILL101_704 VDD VSS sg13g2_FILL8
XSTDFILL101_712 VDD VSS sg13g2_FILL8
XSTDFILL101_720 VDD VSS sg13g2_FILL8
XSTDFILL101_728 VDD VSS sg13g2_FILL8
XSTDFILL101_736 VDD VSS sg13g2_FILL8
XSTDFILL101_744 VDD VSS sg13g2_FILL8
XSTDFILL101_752 VDD VSS sg13g2_FILL8
XSTDFILL101_760 VDD VSS sg13g2_FILL8
XSTDFILL101_768 VDD VSS sg13g2_FILL8
XSTDFILL101_776 VDD VSS sg13g2_FILL8
XSTDFILL101_784 VDD VSS sg13g2_FILL8
XSTDFILL101_792 VDD VSS sg13g2_FILL8
XSTDFILL101_800 VDD VSS sg13g2_FILL8
XSTDFILL101_808 VDD VSS sg13g2_FILL8
XSTDFILL101_816 VDD VSS sg13g2_FILL8
XSTDFILL101_824 VDD VSS sg13g2_FILL8
XSTDFILL101_832 VDD VSS sg13g2_FILL8
XSTDFILL101_840 VDD VSS sg13g2_FILL8
XSTDFILL101_848 VDD VSS sg13g2_FILL8
XSTDFILL101_856 VDD VSS sg13g2_FILL8
XSTDFILL101_864 VDD VSS sg13g2_FILL8
XSTDFILL101_872 VDD VSS sg13g2_FILL8
XSTDFILL101_880 VDD VSS sg13g2_FILL8
XSTDFILL101_888 VDD VSS sg13g2_FILL8
XSTDFILL101_896 VDD VSS sg13g2_FILL8
XSTDFILL101_904 VDD VSS sg13g2_FILL8
XSTDFILL101_912 VDD VSS sg13g2_FILL8
XSTDFILL101_920 VDD VSS sg13g2_FILL8
XSTDFILL101_928 VDD VSS sg13g2_FILL8
XSTDFILL101_936 VDD VSS sg13g2_FILL8
XSTDFILL101_944 VDD VSS sg13g2_FILL8
XSTDFILL101_952 VDD VSS sg13g2_FILL8
XSTDFILL101_960 VDD VSS sg13g2_FILL8
XSTDFILL101_968 VDD VSS sg13g2_FILL8
XSTDFILL101_976 VDD VSS sg13g2_FILL8
XSTDFILL101_984 VDD VSS sg13g2_FILL8
XSTDFILL101_992 VDD VSS sg13g2_FILL8
XSTDFILL101_1000 VDD VSS sg13g2_FILL8
XSTDFILL101_1008 VDD VSS sg13g2_FILL8
XSTDFILL101_1016 VDD VSS sg13g2_FILL8
XSTDFILL101_1024 VDD VSS sg13g2_FILL8
XSTDFILL101_1032 VDD VSS sg13g2_FILL8
XSTDFILL101_1040 VDD VSS sg13g2_FILL8
XSTDFILL101_1048 VDD VSS sg13g2_FILL8
XSTDFILL101_1056 VDD VSS sg13g2_FILL8
XSTDFILL101_1064 VDD VSS sg13g2_FILL8
XSTDFILL101_1072 VDD VSS sg13g2_FILL8
XSTDFILL101_1080 VDD VSS sg13g2_FILL8
XSTDFILL101_1088 VDD VSS sg13g2_FILL8
XSTDFILL101_1096 VDD VSS sg13g2_FILL8
XSTDFILL101_1104 VDD VSS sg13g2_FILL8
XSTDFILL101_1112 VDD VSS sg13g2_FILL8
XSTDFILL101_1120 VDD VSS sg13g2_FILL8
XSTDFILL101_1128 VDD VSS sg13g2_FILL8
XSTDFILL101_1136 VDD VSS sg13g2_FILL8
XSTDFILL101_1144 VDD VSS sg13g2_FILL8
XSTDFILL101_1152 VDD VSS sg13g2_FILL8
XSTDFILL101_1160 VDD VSS sg13g2_FILL8
XSTDFILL101_1168 VDD VSS sg13g2_FILL8
XSTDFILL101_1176 VDD VSS sg13g2_FILL8
XSTDFILL101_1184 VDD VSS sg13g2_FILL8
XSTDFILL101_1192 VDD VSS sg13g2_FILL8
XSTDFILL101_1200 VDD VSS sg13g2_FILL8
XSTDFILL101_1208 VDD VSS sg13g2_FILL8
XSTDFILL101_1216 VDD VSS sg13g2_FILL8
XSTDFILL101_1224 VDD VSS sg13g2_FILL8
XSTDFILL101_1232 VDD VSS sg13g2_FILL8
XSTDFILL101_1240 VDD VSS sg13g2_FILL8
XSTDFILL101_1248 VDD VSS sg13g2_FILL8
XSTDFILL101_1256 VDD VSS sg13g2_FILL8
XSTDFILL101_1264 VDD VSS sg13g2_FILL8
XSTDFILL101_1272 VDD VSS sg13g2_FILL8
XSTDFILL101_1280 VDD VSS sg13g2_FILL8
XSTDFILL101_1288 VDD VSS sg13g2_FILL8
XSTDFILL101_1296 VDD VSS sg13g2_FILL8
XSTDFILL101_1304 VDD VSS sg13g2_FILL8
XSTDFILL101_1312 VDD VSS sg13g2_FILL8
XSTDFILL101_1320 VDD VSS sg13g2_FILL8
XSTDFILL101_1328 VDD VSS sg13g2_FILL8
XSTDFILL101_1336 VDD VSS sg13g2_FILL8
XSTDFILL101_1344 VDD VSS sg13g2_FILL8
XSTDFILL101_1352 VDD VSS sg13g2_FILL8
XSTDFILL101_1360 VDD VSS sg13g2_FILL8
XSTDFILL101_1368 VDD VSS sg13g2_FILL8
XSTDFILL101_1376 VDD VSS sg13g2_FILL8
XSTDFILL101_1384 VDD VSS sg13g2_FILL8
XSTDFILL101_1392 VDD VSS sg13g2_FILL8
XSTDFILL101_1400 VDD VSS sg13g2_FILL8
XSTDFILL101_1408 VDD VSS sg13g2_FILL8
XSTDFILL101_1416 VDD VSS sg13g2_FILL8
XSTDFILL101_1424 VDD VSS sg13g2_FILL8
XSTDFILL101_1432 VDD VSS sg13g2_FILL8
XSTDFILL101_1440 VDD VSS sg13g2_FILL8
XSTDFILL101_1448 VDD VSS sg13g2_FILL8
XSTDFILL101_1456 VDD VSS sg13g2_FILL8
XSTDFILL101_1464 VDD VSS sg13g2_FILL8
XSTDFILL101_1472 VDD VSS sg13g2_FILL8
XSTDFILL101_1480 VDD VSS sg13g2_FILL8
XSTDFILL101_1488 VDD VSS sg13g2_FILL8
XSTDFILL101_1496 VDD VSS sg13g2_FILL8
XSTDFILL101_1504 VDD VSS sg13g2_FILL8
XSTDFILL101_1512 VDD VSS sg13g2_FILL8
XSTDFILL101_1520 VDD VSS sg13g2_FILL8
XSTDFILL101_1528 VDD VSS sg13g2_FILL8
XSTDFILL101_1536 VDD VSS sg13g2_FILL8
XSTDFILL101_1544 VDD VSS sg13g2_FILL8
XSTDFILL101_1552 VDD VSS sg13g2_FILL8
XSTDFILL101_1560 VDD VSS sg13g2_FILL8
XSTDFILL101_1568 VDD VSS sg13g2_FILL8
XSTDFILL101_1576 VDD VSS sg13g2_FILL8
XSTDFILL101_1584 VDD VSS sg13g2_FILL8
XSTDFILL101_1592 VDD VSS sg13g2_FILL8
XSTDFILL101_1600 VDD VSS sg13g2_FILL8
XSTDFILL101_1608 VDD VSS sg13g2_FILL8
XSTDFILL101_1616 VDD VSS sg13g2_FILL8
XSTDFILL101_1624 VDD VSS sg13g2_FILL8
XSTDFILL101_1632 VDD VSS sg13g2_FILL8
XSTDFILL101_1640 VDD VSS sg13g2_FILL8
XSTDFILL101_1648 VDD VSS sg13g2_FILL8
XSTDFILL101_1656 VDD VSS sg13g2_FILL8
XSTDFILL101_1664 VDD VSS sg13g2_FILL8
XSTDFILL101_1672 VDD VSS sg13g2_FILL8
XSTDFILL101_1680 VDD VSS sg13g2_FILL8
XSTDFILL101_1688 VDD VSS sg13g2_FILL8
XSTDFILL101_1696 VDD VSS sg13g2_FILL8
XSTDFILL101_1704 VDD VSS sg13g2_FILL8
XSTDFILL101_1712 VDD VSS sg13g2_FILL8
XSTDFILL101_1720 VDD VSS sg13g2_FILL8
XSTDFILL101_1728 VDD VSS sg13g2_FILL8
XSTDFILL101_1736 VDD VSS sg13g2_FILL8
XSTDFILL101_1744 VDD VSS sg13g2_FILL8
XSTDFILL101_1752 VDD VSS sg13g2_FILL8
XSTDFILL101_1760 VDD VSS sg13g2_FILL8
XSTDFILL101_1768 VDD VSS sg13g2_FILL8
XSTDFILL101_1776 VDD VSS sg13g2_FILL8
XSTDFILL101_1784 VDD VSS sg13g2_FILL8
XSTDFILL101_1792 VDD VSS sg13g2_FILL8
XSTDFILL101_1800 VDD VSS sg13g2_FILL8
XSTDFILL101_1808 VDD VSS sg13g2_FILL8
XSTDFILL101_1816 VDD VSS sg13g2_FILL8
XSTDFILL101_1824 VDD VSS sg13g2_FILL8
XSTDFILL101_1832 VDD VSS sg13g2_FILL8
XSTDFILL101_1840 VDD VSS sg13g2_FILL8
XSTDFILL101_1848 VDD VSS sg13g2_FILL8
XSTDFILL101_1856 VDD VSS sg13g2_FILL8
XSTDFILL101_1864 VDD VSS sg13g2_FILL8
XSTDFILL101_1872 VDD VSS sg13g2_FILL8
XSTDFILL101_1880 VDD VSS sg13g2_FILL8
XSTDFILL101_1888 VDD VSS sg13g2_FILL8
XSTDFILL101_1896 VDD VSS sg13g2_FILL8
XSTDFILL101_1904 VDD VSS sg13g2_FILL8
XSTDFILL101_1912 VDD VSS sg13g2_FILL8
XSTDFILL101_1920 VDD VSS sg13g2_FILL8
XSTDFILL101_1928 VDD VSS sg13g2_FILL8
XSTDFILL101_1936 VDD VSS sg13g2_FILL8
XSTDFILL101_1944 VDD VSS sg13g2_FILL8
XSTDFILL101_1952 VDD VSS sg13g2_FILL8
XSTDFILL101_1960 VDD VSS sg13g2_FILL8
XSTDFILL101_1968 VDD VSS sg13g2_FILL8
XSTDFILL101_1976 VDD VSS sg13g2_FILL8
XSTDFILL101_1984 VDD VSS sg13g2_FILL8
XSTDFILL101_1992 VDD VSS sg13g2_FILL8
XSTDFILL101_2000 VDD VSS sg13g2_FILL8
XSTDFILL101_2008 VDD VSS sg13g2_FILL8
XSTDFILL101_2016 VDD VSS sg13g2_FILL8
XSTDFILL101_2024 VDD VSS sg13g2_FILL8
XSTDFILL101_2032 VDD VSS sg13g2_FILL8
XSTDFILL101_2040 VDD VSS sg13g2_FILL8
XSTDFILL101_2048 VDD VSS sg13g2_FILL8
XSTDFILL101_2056 VDD VSS sg13g2_FILL8
XSTDFILL101_2064 VDD VSS sg13g2_FILL8
XSTDFILL101_2072 VDD VSS sg13g2_FILL8
XSTDFILL101_2080 VDD VSS sg13g2_FILL8
XSTDFILL101_2088 VDD VSS sg13g2_FILL8
XSTDFILL101_2096 VDD VSS sg13g2_FILL8
XSTDFILL101_2104 VDD VSS sg13g2_FILL8
XSTDFILL101_2112 VDD VSS sg13g2_FILL8
XSTDFILL101_2120 VDD VSS sg13g2_FILL8
XSTDFILL101_2128 VDD VSS sg13g2_FILL8
XSTDFILL101_2136 VDD VSS sg13g2_FILL8
XSTDFILL101_2144 VDD VSS sg13g2_FILL8
XSTDFILL101_2152 VDD VSS sg13g2_FILL2
XSTDFILL102_0 VDD VSS sg13g2_FILL8
XSTDFILL102_8 VDD VSS sg13g2_FILL8
XSTDFILL102_16 VDD VSS sg13g2_FILL8
XSTDFILL102_24 VDD VSS sg13g2_FILL8
XSTDFILL102_32 VDD VSS sg13g2_FILL8
XSTDFILL102_40 VDD VSS sg13g2_FILL8
XSTDFILL102_48 VDD VSS sg13g2_FILL8
XSTDFILL102_56 VDD VSS sg13g2_FILL8
XSTDFILL102_64 VDD VSS sg13g2_FILL8
XSTDFILL102_72 VDD VSS sg13g2_FILL8
XSTDFILL102_80 VDD VSS sg13g2_FILL8
XSTDFILL102_88 VDD VSS sg13g2_FILL8
XSTDFILL102_96 VDD VSS sg13g2_FILL8
XSTDFILL102_104 VDD VSS sg13g2_FILL8
XSTDFILL102_112 VDD VSS sg13g2_FILL8
XSTDFILL102_120 VDD VSS sg13g2_FILL8
XSTDFILL102_128 VDD VSS sg13g2_FILL8
XSTDFILL102_136 VDD VSS sg13g2_FILL8
XSTDFILL102_144 VDD VSS sg13g2_FILL8
XSTDFILL102_152 VDD VSS sg13g2_FILL8
XSTDFILL102_160 VDD VSS sg13g2_FILL8
XSTDFILL102_168 VDD VSS sg13g2_FILL8
XSTDFILL102_176 VDD VSS sg13g2_FILL8
XSTDFILL102_184 VDD VSS sg13g2_FILL8
XSTDFILL102_192 VDD VSS sg13g2_FILL8
XSTDFILL102_200 VDD VSS sg13g2_FILL8
XSTDFILL102_208 VDD VSS sg13g2_FILL8
XSTDFILL102_216 VDD VSS sg13g2_FILL8
XSTDFILL102_224 VDD VSS sg13g2_FILL8
XSTDFILL102_232 VDD VSS sg13g2_FILL8
XSTDFILL102_240 VDD VSS sg13g2_FILL8
XSTDFILL102_248 VDD VSS sg13g2_FILL8
XSTDFILL102_256 VDD VSS sg13g2_FILL8
XSTDFILL102_264 VDD VSS sg13g2_FILL8
XSTDFILL102_272 VDD VSS sg13g2_FILL8
XSTDFILL102_280 VDD VSS sg13g2_FILL8
XSTDFILL102_288 VDD VSS sg13g2_FILL8
XSTDFILL102_296 VDD VSS sg13g2_FILL8
XSTDFILL102_304 VDD VSS sg13g2_FILL8
XSTDFILL102_312 VDD VSS sg13g2_FILL8
XSTDFILL102_320 VDD VSS sg13g2_FILL8
XSTDFILL102_328 VDD VSS sg13g2_FILL8
XSTDFILL102_336 VDD VSS sg13g2_FILL8
XSTDFILL102_344 VDD VSS sg13g2_FILL8
XSTDFILL102_352 VDD VSS sg13g2_FILL8
XSTDFILL102_360 VDD VSS sg13g2_FILL8
XSTDFILL102_368 VDD VSS sg13g2_FILL8
XSTDFILL102_376 VDD VSS sg13g2_FILL8
XSTDFILL102_384 VDD VSS sg13g2_FILL8
XSTDFILL102_392 VDD VSS sg13g2_FILL8
XSTDFILL102_400 VDD VSS sg13g2_FILL8
XSTDFILL102_408 VDD VSS sg13g2_FILL8
XSTDFILL102_416 VDD VSS sg13g2_FILL8
XSTDFILL102_424 VDD VSS sg13g2_FILL8
XSTDFILL102_432 VDD VSS sg13g2_FILL8
XSTDFILL102_440 VDD VSS sg13g2_FILL8
XSTDFILL102_448 VDD VSS sg13g2_FILL8
XSTDFILL102_456 VDD VSS sg13g2_FILL8
XSTDFILL102_464 VDD VSS sg13g2_FILL8
XSTDFILL102_472 VDD VSS sg13g2_FILL8
XSTDFILL102_480 VDD VSS sg13g2_FILL8
XSTDFILL102_488 VDD VSS sg13g2_FILL8
XSTDFILL102_496 VDD VSS sg13g2_FILL8
XSTDFILL102_504 VDD VSS sg13g2_FILL8
XSTDFILL102_512 VDD VSS sg13g2_FILL8
XSTDFILL102_520 VDD VSS sg13g2_FILL8
XSTDFILL102_528 VDD VSS sg13g2_FILL8
XSTDFILL102_536 VDD VSS sg13g2_FILL8
XSTDFILL102_544 VDD VSS sg13g2_FILL8
XSTDFILL102_552 VDD VSS sg13g2_FILL8
XSTDFILL102_560 VDD VSS sg13g2_FILL8
XSTDFILL102_568 VDD VSS sg13g2_FILL8
XSTDFILL102_576 VDD VSS sg13g2_FILL8
XSTDFILL102_584 VDD VSS sg13g2_FILL8
XSTDFILL102_592 VDD VSS sg13g2_FILL8
XSTDFILL102_600 VDD VSS sg13g2_FILL8
XSTDFILL102_608 VDD VSS sg13g2_FILL8
XSTDFILL102_616 VDD VSS sg13g2_FILL8
XSTDFILL102_624 VDD VSS sg13g2_FILL8
XSTDFILL102_632 VDD VSS sg13g2_FILL8
XSTDFILL102_640 VDD VSS sg13g2_FILL8
XSTDFILL102_648 VDD VSS sg13g2_FILL8
XSTDFILL102_656 VDD VSS sg13g2_FILL8
XSTDFILL102_664 VDD VSS sg13g2_FILL8
XSTDFILL102_672 VDD VSS sg13g2_FILL8
XSTDFILL102_680 VDD VSS sg13g2_FILL8
XSTDFILL102_688 VDD VSS sg13g2_FILL8
XSTDFILL102_696 VDD VSS sg13g2_FILL8
XSTDFILL102_704 VDD VSS sg13g2_FILL8
XSTDFILL102_712 VDD VSS sg13g2_FILL8
XSTDFILL102_720 VDD VSS sg13g2_FILL8
XSTDFILL102_728 VDD VSS sg13g2_FILL8
XSTDFILL102_736 VDD VSS sg13g2_FILL8
XSTDFILL102_744 VDD VSS sg13g2_FILL8
XSTDFILL102_752 VDD VSS sg13g2_FILL8
XSTDFILL102_760 VDD VSS sg13g2_FILL8
XSTDFILL102_768 VDD VSS sg13g2_FILL8
XSTDFILL102_776 VDD VSS sg13g2_FILL8
XSTDFILL102_784 VDD VSS sg13g2_FILL8
XSTDFILL102_792 VDD VSS sg13g2_FILL8
XSTDFILL102_800 VDD VSS sg13g2_FILL8
XSTDFILL102_808 VDD VSS sg13g2_FILL8
XSTDFILL102_816 VDD VSS sg13g2_FILL8
XSTDFILL102_824 VDD VSS sg13g2_FILL8
XSTDFILL102_832 VDD VSS sg13g2_FILL8
XSTDFILL102_840 VDD VSS sg13g2_FILL8
XSTDFILL102_848 VDD VSS sg13g2_FILL8
XSTDFILL102_856 VDD VSS sg13g2_FILL8
XSTDFILL102_864 VDD VSS sg13g2_FILL8
XSTDFILL102_872 VDD VSS sg13g2_FILL8
XSTDFILL102_880 VDD VSS sg13g2_FILL8
XSTDFILL102_888 VDD VSS sg13g2_FILL8
XSTDFILL102_896 VDD VSS sg13g2_FILL8
XSTDFILL102_904 VDD VSS sg13g2_FILL8
XSTDFILL102_912 VDD VSS sg13g2_FILL8
XSTDFILL102_920 VDD VSS sg13g2_FILL8
XSTDFILL102_928 VDD VSS sg13g2_FILL8
XSTDFILL102_936 VDD VSS sg13g2_FILL8
XSTDFILL102_944 VDD VSS sg13g2_FILL8
XSTDFILL102_952 VDD VSS sg13g2_FILL8
XSTDFILL102_960 VDD VSS sg13g2_FILL8
XSTDFILL102_968 VDD VSS sg13g2_FILL8
XSTDFILL102_976 VDD VSS sg13g2_FILL8
XSTDFILL102_984 VDD VSS sg13g2_FILL8
XSTDFILL102_992 VDD VSS sg13g2_FILL8
XSTDFILL102_1000 VDD VSS sg13g2_FILL8
XSTDFILL102_1008 VDD VSS sg13g2_FILL8
XSTDFILL102_1016 VDD VSS sg13g2_FILL8
XSTDFILL102_1024 VDD VSS sg13g2_FILL8
XSTDFILL102_1032 VDD VSS sg13g2_FILL8
XSTDFILL102_1040 VDD VSS sg13g2_FILL8
XSTDFILL102_1048 VDD VSS sg13g2_FILL8
XSTDFILL102_1056 VDD VSS sg13g2_FILL8
XSTDFILL102_1064 VDD VSS sg13g2_FILL8
XSTDFILL102_1072 VDD VSS sg13g2_FILL8
XSTDFILL102_1080 VDD VSS sg13g2_FILL8
XSTDFILL102_1088 VDD VSS sg13g2_FILL8
XSTDFILL102_1096 VDD VSS sg13g2_FILL8
XSTDFILL102_1104 VDD VSS sg13g2_FILL8
XSTDFILL102_1112 VDD VSS sg13g2_FILL8
XSTDFILL102_1120 VDD VSS sg13g2_FILL8
XSTDFILL102_1128 VDD VSS sg13g2_FILL8
XSTDFILL102_1136 VDD VSS sg13g2_FILL8
XSTDFILL102_1144 VDD VSS sg13g2_FILL8
XSTDFILL102_1152 VDD VSS sg13g2_FILL8
XSTDFILL102_1160 VDD VSS sg13g2_FILL8
XSTDFILL102_1168 VDD VSS sg13g2_FILL8
XSTDFILL102_1176 VDD VSS sg13g2_FILL8
XSTDFILL102_1184 VDD VSS sg13g2_FILL8
XSTDFILL102_1192 VDD VSS sg13g2_FILL8
XSTDFILL102_1200 VDD VSS sg13g2_FILL8
XSTDFILL102_1208 VDD VSS sg13g2_FILL8
XSTDFILL102_1216 VDD VSS sg13g2_FILL8
XSTDFILL102_1224 VDD VSS sg13g2_FILL8
XSTDFILL102_1232 VDD VSS sg13g2_FILL8
XSTDFILL102_1240 VDD VSS sg13g2_FILL8
XSTDFILL102_1248 VDD VSS sg13g2_FILL8
XSTDFILL102_1256 VDD VSS sg13g2_FILL8
XSTDFILL102_1264 VDD VSS sg13g2_FILL8
XSTDFILL102_1272 VDD VSS sg13g2_FILL8
XSTDFILL102_1280 VDD VSS sg13g2_FILL8
XSTDFILL102_1288 VDD VSS sg13g2_FILL8
XSTDFILL102_1296 VDD VSS sg13g2_FILL8
XSTDFILL102_1304 VDD VSS sg13g2_FILL8
XSTDFILL102_1312 VDD VSS sg13g2_FILL8
XSTDFILL102_1320 VDD VSS sg13g2_FILL8
XSTDFILL102_1328 VDD VSS sg13g2_FILL8
XSTDFILL102_1336 VDD VSS sg13g2_FILL8
XSTDFILL102_1344 VDD VSS sg13g2_FILL8
XSTDFILL102_1352 VDD VSS sg13g2_FILL8
XSTDFILL102_1360 VDD VSS sg13g2_FILL8
XSTDFILL102_1368 VDD VSS sg13g2_FILL8
XSTDFILL102_1376 VDD VSS sg13g2_FILL8
XSTDFILL102_1384 VDD VSS sg13g2_FILL8
XSTDFILL102_1392 VDD VSS sg13g2_FILL8
XSTDFILL102_1400 VDD VSS sg13g2_FILL8
XSTDFILL102_1408 VDD VSS sg13g2_FILL8
XSTDFILL102_1416 VDD VSS sg13g2_FILL8
XSTDFILL102_1424 VDD VSS sg13g2_FILL8
XSTDFILL102_1432 VDD VSS sg13g2_FILL8
XSTDFILL102_1440 VDD VSS sg13g2_FILL8
XSTDFILL102_1448 VDD VSS sg13g2_FILL8
XSTDFILL102_1456 VDD VSS sg13g2_FILL8
XSTDFILL102_1464 VDD VSS sg13g2_FILL8
XSTDFILL102_1472 VDD VSS sg13g2_FILL8
XSTDFILL102_1480 VDD VSS sg13g2_FILL8
XSTDFILL102_1488 VDD VSS sg13g2_FILL8
XSTDFILL102_1496 VDD VSS sg13g2_FILL8
XSTDFILL102_1504 VDD VSS sg13g2_FILL8
XSTDFILL102_1512 VDD VSS sg13g2_FILL8
XSTDFILL102_1520 VDD VSS sg13g2_FILL8
XSTDFILL102_1528 VDD VSS sg13g2_FILL8
XSTDFILL102_1536 VDD VSS sg13g2_FILL8
XSTDFILL102_1544 VDD VSS sg13g2_FILL8
XSTDFILL102_1552 VDD VSS sg13g2_FILL8
XSTDFILL102_1560 VDD VSS sg13g2_FILL8
XSTDFILL102_1568 VDD VSS sg13g2_FILL8
XSTDFILL102_1576 VDD VSS sg13g2_FILL8
XSTDFILL102_1584 VDD VSS sg13g2_FILL8
XSTDFILL102_1592 VDD VSS sg13g2_FILL8
XSTDFILL102_1600 VDD VSS sg13g2_FILL8
XSTDFILL102_1608 VDD VSS sg13g2_FILL8
XSTDFILL102_1616 VDD VSS sg13g2_FILL8
XSTDFILL102_1624 VDD VSS sg13g2_FILL8
XSTDFILL102_1632 VDD VSS sg13g2_FILL8
XSTDFILL102_1640 VDD VSS sg13g2_FILL8
XSTDFILL102_1648 VDD VSS sg13g2_FILL8
XSTDFILL102_1656 VDD VSS sg13g2_FILL8
XSTDFILL102_1664 VDD VSS sg13g2_FILL8
XSTDFILL102_1672 VDD VSS sg13g2_FILL8
XSTDFILL102_1680 VDD VSS sg13g2_FILL8
XSTDFILL102_1688 VDD VSS sg13g2_FILL8
XSTDFILL102_1696 VDD VSS sg13g2_FILL8
XSTDFILL102_1704 VDD VSS sg13g2_FILL8
XSTDFILL102_1712 VDD VSS sg13g2_FILL8
XSTDFILL102_1720 VDD VSS sg13g2_FILL8
XSTDFILL102_1728 VDD VSS sg13g2_FILL8
XSTDFILL102_1736 VDD VSS sg13g2_FILL8
XSTDFILL102_1744 VDD VSS sg13g2_FILL8
XSTDFILL102_1752 VDD VSS sg13g2_FILL8
XSTDFILL102_1760 VDD VSS sg13g2_FILL8
XSTDFILL102_1768 VDD VSS sg13g2_FILL8
XSTDFILL102_1776 VDD VSS sg13g2_FILL8
XSTDFILL102_1784 VDD VSS sg13g2_FILL8
XSTDFILL102_1792 VDD VSS sg13g2_FILL8
XSTDFILL102_1800 VDD VSS sg13g2_FILL8
XSTDFILL102_1808 VDD VSS sg13g2_FILL8
XSTDFILL102_1816 VDD VSS sg13g2_FILL8
XSTDFILL102_1824 VDD VSS sg13g2_FILL8
XSTDFILL102_1832 VDD VSS sg13g2_FILL8
XSTDFILL102_1840 VDD VSS sg13g2_FILL8
XSTDFILL102_1848 VDD VSS sg13g2_FILL8
XSTDFILL102_1856 VDD VSS sg13g2_FILL8
XSTDFILL102_1864 VDD VSS sg13g2_FILL8
XSTDFILL102_1872 VDD VSS sg13g2_FILL8
XSTDFILL102_1880 VDD VSS sg13g2_FILL8
XSTDFILL102_1888 VDD VSS sg13g2_FILL8
XSTDFILL102_1896 VDD VSS sg13g2_FILL8
XSTDFILL102_1904 VDD VSS sg13g2_FILL8
XSTDFILL102_1912 VDD VSS sg13g2_FILL8
XSTDFILL102_1920 VDD VSS sg13g2_FILL8
XSTDFILL102_1928 VDD VSS sg13g2_FILL8
XSTDFILL102_1936 VDD VSS sg13g2_FILL8
XSTDFILL102_1944 VDD VSS sg13g2_FILL8
XSTDFILL102_1952 VDD VSS sg13g2_FILL8
XSTDFILL102_1960 VDD VSS sg13g2_FILL8
XSTDFILL102_1968 VDD VSS sg13g2_FILL8
XSTDFILL102_1976 VDD VSS sg13g2_FILL8
XSTDFILL102_1984 VDD VSS sg13g2_FILL8
XSTDFILL102_1992 VDD VSS sg13g2_FILL8
XSTDFILL102_2000 VDD VSS sg13g2_FILL8
XSTDFILL102_2008 VDD VSS sg13g2_FILL8
XSTDFILL102_2016 VDD VSS sg13g2_FILL8
XSTDFILL102_2024 VDD VSS sg13g2_FILL8
XSTDFILL102_2032 VDD VSS sg13g2_FILL8
XSTDFILL102_2040 VDD VSS sg13g2_FILL8
XSTDFILL102_2048 VDD VSS sg13g2_FILL8
XSTDFILL102_2056 VDD VSS sg13g2_FILL8
XSTDFILL102_2064 VDD VSS sg13g2_FILL8
XSTDFILL102_2072 VDD VSS sg13g2_FILL8
XSTDFILL102_2080 VDD VSS sg13g2_FILL8
XSTDFILL102_2088 VDD VSS sg13g2_FILL8
XSTDFILL102_2096 VDD VSS sg13g2_FILL8
XSTDFILL102_2104 VDD VSS sg13g2_FILL8
XSTDFILL102_2112 VDD VSS sg13g2_FILL8
XSTDFILL102_2120 VDD VSS sg13g2_FILL8
XSTDFILL102_2128 VDD VSS sg13g2_FILL8
XSTDFILL102_2136 VDD VSS sg13g2_FILL8
XSTDFILL102_2144 VDD VSS sg13g2_FILL8
XSTDFILL102_2152 VDD VSS sg13g2_FILL2
Xseal sealring
.ENDS asicone_202508
