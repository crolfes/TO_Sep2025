* Extracted by KLayout with SG13G2 LVS runset on : 28/08/2025 21:02

.SUBCKT asicone_202508 AVDD|anode|cathode|pad|vdd
+ anode|cathode|pad|pad_adc_rst_pad anode|cathode|pad|pad_adc_clk_pad
+ anode|cathode|pad|pad_adc_result_0_pad anode|cathode|pad|pad_adc_result_1_pad
+ anode|cathode|pad|pad_adc_result_2_pad anode|cathode|pad|pad_adc_result_3_pad
+ anode|cathode|pad|pad_adc_result_4_pad anode|cathode|pad|pad_adc_valid_pad
+ anode|cathode|pad|pad_adc_sample_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply VSSIO|anode|cathode|guard|iovss
+ gate|ngate|o gate|ngate|o$1 gate|ngate|o$2 gate|ngate|o$3 gate|ngate|o$4
+ gate|ngate|o$5 gate|ngate|o$6 gate|o|pgate gate|o|pgate$1 gate|o|pgate$2
+ gate|o|pgate$3 gate|o|pgate$4 gate|o|pgate$5 gate|o|pgate$6 core|padres core
+ core$1 VDD|pad|pin1|supply|vdd RESULT[0]|c2p|core|i|q RESULT[1]|c2p|core|i|q
+ RESULT[2]|c2p|core|i|q RESULT[3]|c2p|core|i|q RESULT[4]|c2p|core|i|q
+ VALID|a3|c2p|core|i|z SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|vss
+ RST|a1|b|cdn|core|i|p2c CLK|core|i|p2c anode|cathode|pad|pad_adc_go_pad i|z z
+ zn z$1 z$2 i|z$1 z$3 z$4 i|z$2 z$5 GO|a2|core|p2c core$2 d|zn a2|zn a1|z b|zn
+ z$6 zn$1 d|z b|zn$1 a1|z$1 a1|z$2 a1|z$3 a1|b|i|q a2|a3|zn a1|b|i|q$1 a2|z
+ a1|a2|a3|z d|zn$1 a2|zn$1 a1|z$4 d|z$1 cp|z a2 VIP|core|padres z$7
+ VIN|core|padres cp|z$1 anode|cathode|pad|pad_adc_vrefp_pad d|zn$2
+ VREFH|core|padres a2$1 z$8 z$9 a2|z$1 z$10 d|z$2 a2|z$2 a2|zn$2 a1|z$5 d|zn$3
+ b|zn$2 a1|z$6 a1|z$7 a1|b|i|q$2 d|zn$4 a1|z$8 d|zn$5 a1|z$9 a2|d|zn a2|zn$3
+ i|z$3 z$11 z$12 z$13 b|q a2|i|q z$14 z$15 z$16 z$17 zn$2 d|z$3 z$18 z$19
+ a2|zn$4 d|zn$6 z$20 i|z$4 a1|b|i|q$3 a2|a3|z a1|z$10 b|zn$3 a2|z$3 a2|zn$5
+ in|pin2 a1|i|q gate|out anode|cathode|pad|pad_adc_vrefn_pad i|zn i|z$5 i|z$6
+ i|z|zn i|z$7 z$21 i|z$8 cp|z$2 i|z$9 d|zn$7 i|z$10 i|z$11 i|z|zn$1 i|z$12
+ i|zn$1 i|z$13 i|z$14 i|z|zn$2 d|zn$8 VREFL|core|padres i|z$15 i|zn$2 i|z$16
+ i|z|zn$3 i|z$17 i|z$18 i|z$19 i|z$20 i|z$21 i|z|zn$4 i|z$22 a1|i|z|zn i|z$23
+ i|zn$3 i|z|zn$5 i|z$24 i|z$25 i|z|zn$6 i|z$26 i|z$27 i|z$28 i|z$29 i|z$30
+ i|zn$4 i|zn$5 i|z$31 i|z$32 i|zn$6 i|z$33 a2|z$4 i|z$34 i|z$35 i|z$36 a1|z$11
+ i|zn$7 i|z$37 i|z|zn$7 i|z$38 i|z|zn$8 i|z$39 i|z$40 a2|i|z i|z$41 a2|z$5
+ i|z$42 i|z$43 i|z$44 i|z$45 i|z$46 i|z$47 i|zn$8 i|z$48 a1|i|q$1 i|z$49
+ i|z$50 i|z$51 i|z$52 i|z$53 i|z$54 a1|c|i|zn i|z$55 z$22 z$23 i|z$56 i|z$57
+ i|zn$9 i|zn$10 i|z$58 i|z$59 i|z$60 i|z$61 a2|b|z i|z$62 i|z$63 i|z$64 i|z$65
+ z$24 a1|c|i|zn$1 i|z$66 z$25 i|z$67 i|z$68 i|zn$11 i|z$69 i|z$70 i|z$71
+ i|z|zn$9 i|z$72 i|z$73 i|z$74 i|z$75 i|z$76 i|z$77 b|i|q i|z$78 i|z$79
+ b|i|q$1 i|z$80 i|z$81 i|z$82 i|z$83 i|z$84 i|z$85 i|z$86 a1|z$12 i|z$87
+ i|z$88 i|z$89 i|zn$12 i|z$90 i|z$91 i|z$92 b|i|q$2 i|z$93 i|z$94 i|zn$13
+ i|z$95 i|z$96 b|zn$4 cp|i|z zn$3 i|z$97 i|z$98 i|z$99 i|z$100 i|z$101 b|i|q$3
+ i|z$102 i|z$103 i|z$104 i|z$105 i|z$106 i|z$107 i|z$108 i|z$109 i|z$110
+ a2|zn$6 a1|z$13 zn$4 i|z$111 i|z$112 i|z$113 i|z$114 cp|z$3 d|zn$9 d|zn$10
+ a2|z$6 anode|cathode|pad|pad_adc_vin_pad b|zn$5 z$26 d|z$4 a2|z$7 b|zn$6
+ RD[8]|a4|z RD[9]|a4|z z$27 zn$5 gate|out$1 in|pin2$1
+ anode|cathode|pad|pad_adc_vip_pad anode|cathode|pad
+ anode|cathode|pad|pad_miso_pad gate|o|pgate$7 core|padres$1
+ DOUT_DAT|c2p|core|i|q gate|ngate|o$7 RD[1]|a2|z RD[13]|a4|zn RD[0]|a2|z i i$1
+ RD[19]|a4|z RD[35]|a2|z RD[21]|a4|z RD[45]|a4|z RD[47]|a4|z RD[3]|a2|z
+ RD[38]|a2|z RD[44]|a4|z RD[24]|a2|z RD[46]|a4|z RD[17]|a4|z RD[34]|a2|z
+ RD[40]|a4|z RD[42]|a4|z RD[37]|a2|z RD[36]|a2|z RD[43]|a4|z RD[33]|a2|z
+ RD[2]|a2|z RD[32]|a2|z RD[4]|a2|z RD[39]|a2|z RD[41]|a4|z R[13]|i|i0|q
+ R[12]|i|i0|q R[15]|i|i0|q i$2 R[8]|i|i0|q R[14]|i|i0|q R[2]|i|i0|q
+ R[5]|i|i0|q R[11]|i|i0|q R[9]|i|i0|q R[3]|i|i0|q R[4]|i|i0|q R[1]|i|i0|q
+ R[0]|i|i0|q i$3 i$4 RD[27]|a2|zn R[7]|i|i0|q RD[5]|a2|zn RD[7]|a2|zn
+ RD[31]|a2|zn RD[14]|a4|zn RD[12]|a4|zn RD[10]|a4|zn RD[18]|a4|zn RD[16]|a4|zn
+ RD[11]|a4|zn RD[20]|a4|zn RD[25]|a2|zn RD[15]|a4|zn RD[22]|a4|zn RD[29]|a2|zn
+ anode|cathode|pad|pad_mosi_pad anode|cathode|pad$1 CLK|core|i|p2c$1
+ DATA|core|i0|i1|p2c CEB|a1|core|i|p2c R[30]|i0|q R[17]|i0|q R[39]|i1|q
+ R[21]|i0|q R[43]|i0|q R[41]|i0|q R[22]|i0|q R[33]|i1|q core|padres$2
+ R[42]|i0|q R[47]|i0|q s|zn a1|zn s|zn$1 d|z$5 R[56]|i1|q d|z$6 a1|zn$1
+ a2|zn$7 a1|zn$2 a1|z$14 a1|zn$3 a2|zn$8 a2|zn$9 a2|z$8 a4|zn a2|zn$10 d|z$7
+ d|z$8 R[48]|i1|q i0|i1|q a2|zn$11 R[59]|i1|q cp|z$4 i0|i1|q$1 a2|z$9
+ a1|a3|i|i1|q a2|a3|zn$1 a1|zn$4 a3|zn a1|zn$5 RD[26]|a2|z a2|a3|z$1 a1|z$15
+ a1|zn$6 a1|zn$7 a1|i|i0|i1|q RD[28]|a2|z cp|i|z$1 core$3 a4|zn$1 a2|zn$12
+ R[51]|i1|q a1|zn$8 R[50]|i1|q a3|zn$1 s|zn$2 a1|zn$9 a4|z d|z$9 a4|zn$2
+ a3|zn$2 i1|zn a2|zn$13 a1|zn$10 a2|zn$14 a2|zn$15 a2|zn$16 a4|zn$3 i1|zn$1
+ a4|zn$4 a2|zn$17 a1|zn$11 a1|zn$12 a1|zn$13 d|z$10 R[35]|i1|q a2|z$10
+ i0|i1|q$2 a2|i|i0|i1|q a1|a3|z a3|zn$3 a1|zn$14 R[58]|i1|q d|z$11 i1|z d|z$12
+ d|z$13 d|z$14 a2|zn$18 a3|zn$4 a1|zn$15 a1|zn$16 i1|z$1 a3|zn$5 a2|zn$19
+ a2|zn$20 a3|zn$6 a3|zn$7 d|z$15 d|z$16 R[60]|i1|q i0|i1|q$3 R[55]|i1|q
+ R[53]|i1|q RD[30]|a2|z RD[23]|a4|z RD[6]|a2|zn a1|zn$17 a1|zn$18 s|z d|z$17
+ d|z$18 a2|zn$21 a4|z$1 a2|zn$22 a2|zn$23 i1|z$2 a1|zn$19 a2|zn$24 a4|zn$5
+ a2|zn$25 i1|z$3 d|z$19 R[6]|i|i0|q i0|i1|q$4 i0|i1|q$5 R[37]|i1|q d|z$20
+ a1|zn$20 R[63]|i1|q d|z$21 d|z$22 d|z$23 d|z$24 i0|i1|q$6 R[57]|i1|q
+ R[62]|i1|q i0|i1|q$7 cp|i|z$2 a1|z$16 cp|i|z$3 d|z$25 R[61]|i1|q R[54]|i1|q
+ d|z$26 i1|zn$2 d|z$27 R[52]|i1|q d|z$28 R[49]|i1|q a2|zn$26 s|z$1 R[27]|i0|q
+ d|z$29 R[34]|i1|q d|z$30 d|z$31 z$28 R[28]|i0|q d|z$32 R[31]|i0|q d|z$33
+ d|z$34 R[25]|i0|q d|z$35 a2|zn$27 d|z$36 d|z$37 i|z$115 a1|a2|a4|z s|zn$3
+ d|z$38 d|z$39 R[32]|i1|q a2|z$11 z$29 R[45]|i0|q R[38]|i1|q d|z$40 d|z$41
+ anode|cathode|pad|pad_sclk_pad anode|cathode|pad$2 s|zn$4 d|z$42 d|z$43 z$30
+ R[36]|i1|q a2|z$12 d|z$44 R[19]|i0|q d|z$45 d|z$46 d|z$47 d|z$48 a2|zn$28
+ a2|zn$29 d|z$49 R[24]|i0|q R[29]|i0|q d|z$50 d|z$51 d|z$52 d|z$53 d|z$54
+ R[10]|i|i0|q d|z$55 R[44]|i0|q R[26]|i0|q d|z$56 core|padres$3 a2|zn$30
+ a3|zn$8 d|z$57 i0|z d|z$58 a2|i|s|zn a1|a2|b|q|s a1|zn$21 b|z a2|zn$31
+ a1|i0|q i0|i1|q$8 d|z$59 R[40]|i0|q R[46]|i0|q d|z$60 d|z$61 d|z$62 d|z$63
+ R[18]|i0|q d|z$64 i0|z$1 d|z$65 cp|i|z$4 cp|i|z$5 d|z$66 cp|i|z$6 i0|i1|q$9
+ core$4 s|zn$5 s|zn$6 d|z$67 d|z$68 d|z$69 cp|i|z$7 d|z$70 R[16]|i0|q d|z$71
+ d|z$72 d|z$73 i0|z$2 R[23]|i0|q d|z$74 d|z$75 d|z$76 d|z$77 i0|i1|q$10
+ R[20]|i0|q i0|z$3 d|z$78 d|z$79 d|z$80 d|z$81 i0|z$4 i0|z$5 i0|i1|q$11
+ i0|i1|q$12 i0|i1|q$13 z$31 d|z$82 d|z$83 d|z$84 d|z$85 a1|a2|q d|z$86 z$32
+ i0|z$6 DOUT_EN|z d|s|zn d|z$87 a1|a2|q$1 d|z$88 a1|zn$22 a2|zn$32 a2|q
+ a1|a2|q$2 a1|i0|q$1 z$33 a1|i1|q a2|i|q$1 a2|z$13 d|z$89 d|z$90 d|z$91 a2|q$1
+ a4|zn$6 a1|a2|q$3 a3|zn$9 z$34 a1|i0|q$2 a2|zn$33 a1|a2|q$4 d|z$92 a2|q$2
+ a2|d|z d|z$93 d|z$94 anode|cathode|pad|pad_cs_pad anode|cathode|pad$3 d|z$95
+ a1|z$17 d|z$96 d|z$97 d|s|z a3|zn$10 a2|q$3 a1|b|d|z a2|zn$34 d|z$98
+ a1|a2|q$5 a2|i|q$2 a3|zn$11 a1|zn$23 a4|zn$7 d|z$99 a1|a2|q$6 d|z$100 a4|zn$8
+ a2|q$4 a1|a2|q$7 a2|q$5 d|z$101 a2|q$6 a2|zn$35 a2|q$7 d|z$102 d|z$103
+ d|z$104 d|z$105 a1|a2|q$8 a2|q$8 core|padres$4 d|z$106 d|z$107 d|z$108
+ a1|a2|q$9 core$5 core|padres$5 anode|cathode|pad$4 core|padres$6
+ anode|cathode|pad$5 core|padres$7 anode|cathode|pad$6 core|padres$8
+ anode|cathode|pad$7 core|padres$9 anode|cathode|pad$8 core|padres$10
+ anode|cathode|pad$9 core|padres$11 anode|cathode|pad$10 core|padres$12
+ anode|cathode|pad$11 core|padres$13 anode|cathode|pad$12 core|padres$14
+ anode|cathode|pad$13
M$1 RST|a1|b|cdn|core|i|p2c \$64423 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$2 CLK|core|i|p2c \$64425 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$3 \$63550 RESULT[0]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$4 \$63551 RESULT[0]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$5 \$63553 RESULT[1]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$6 \$63554 RESULT[1]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$7 \$63556 RESULT[2]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$8 \$63557 RESULT[2]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$9 \$63559 RESULT[3]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$10 \$63560 RESULT[3]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$11 \$63562 RESULT[4]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$12 \$63563 RESULT[4]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$13 \$63565 VALID|a3|c2p|core|i|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$14 \$63566 VALID|a3|c2p|core|i|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$15 \$63568 SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$16 \$63569 SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$17 \$89697 \$90053 \$89697 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$53 \$89698 \$90054 \$89698 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$89 \$89699 \$90055 \$89699 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$125 \$89700 \$90056 \$89700 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$161 \$89701 \$90057 \$89701 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$197 \$89702 \$90058 \$89702 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$233 \$89703 \$90059 \$89703 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$269 \$89704 \$90060 \$89704 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$305 \$89705 \$90061 \$89705 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$341 \$89706 \$90062 \$89706 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$737 VSS|anode|cathode|vss a2|zn \$92361 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$738 \$92361 a1|z d|zn VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$739 d|zn b|zn VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$740 GO|a2|core|p2c \$90574 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$741 \$94944 \$95043 \$94944 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$753 \$93030 z$6 \$93030 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$754 \$90053 zn$1 \$93030 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$755 \$90053 z$6 \$90053 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$770 \$93031 zn$1 \$90053 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$771 \$93031 z$6 \$93031 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$786 \$93032 zn$1 \$90053 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$787 \$93032 z$6 \$93032 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$789 \$94945 \$95044 \$94945 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=829.44u AS=354.5856p AD=354.5856p PS=1883.52u PD=1883.52u
M$801 \$93033 z$6 \$93033 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$802 \$90054 zn$1 \$93033 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$803 \$90054 z$6 \$90054 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$818 \$93034 zn$1 \$90054 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$819 \$93034 z$6 \$93034 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$834 \$93035 zn$1 \$90054 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$835 \$93035 z$6 \$93035 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$849 \$93036 z$6 \$93036 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$850 \$90055 zn$1 \$93036 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$851 \$90055 z$6 \$90055 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$866 \$93037 zn$1 \$90055 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$867 \$93037 z$6 \$93037 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$882 \$93038 zn$1 \$90055 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$883 \$93038 z$6 \$93038 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$897 \$93039 z$6 \$93039 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$898 \$90056 zn$1 \$93039 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$899 \$90056 z$6 \$90056 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$914 \$93040 zn$1 \$90056 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$915 \$93040 z$6 \$93040 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$930 \$93041 zn$1 \$90056 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$931 \$93041 z$6 \$93041 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$945 \$93042 z$6 \$93042 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$946 \$90057 zn$1 \$93042 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$947 \$90057 z$6 \$90057 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$962 \$93043 zn$1 \$90057 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$963 \$93043 z$6 \$93043 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$978 \$93044 zn$1 \$90057 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$979 \$93044 z$6 \$93044 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$993 \$93045 z$6 \$93045 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$994 \$90058 zn$1 \$93045 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$995 \$90058 z$6 \$90058 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1010 \$93046 zn$1 \$90058 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1011 \$93046 z$6 \$93046 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1026 \$93047 zn$1 \$90058 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1027 \$93047 z$6 \$93047 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1041 \$93048 z$6 \$93048 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1042 \$90059 zn$1 \$93048 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1043 \$90059 z$6 \$90059 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1058 \$93049 zn$1 \$90059 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1059 \$93049 z$6 \$93049 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1074 \$93050 zn$1 \$90059 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1075 \$93050 z$6 \$93050 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1089 \$93051 z$6 \$93051 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1090 \$90060 zn$1 \$93051 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1091 \$90060 z$6 \$90060 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1106 \$93052 zn$1 \$90060 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1107 \$93052 z$6 \$93052 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1122 \$93053 zn$1 \$90060 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1123 \$93053 z$6 \$93053 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1137 \$93054 z$6 \$93054 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1138 \$90061 zn$1 \$93054 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1139 \$90061 z$6 \$90061 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1154 \$93055 zn$1 \$90061 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1155 \$93055 z$6 \$93055 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1170 \$93056 zn$1 \$90061 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1171 \$93056 z$6 \$93056 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1173 \$94946 \$95045 \$94946 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$1185 \$93057 z$6 \$93057 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1186 \$90062 zn$1 \$93057 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1187 \$90062 z$6 \$90062 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1202 \$93058 zn$1 \$90062 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1203 \$93058 z$6 \$93058 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1218 \$93059 zn$1 \$90062 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1219 \$93059 z$6 \$93059 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1581 \$94578 a1|z$3 \$95725 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$1582 VSS|anode|cathode|vss a2|z \$95725 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.655u AS=0.2901875p AD=0.271825p PS=1.55u PD=1.485u
M$1583 VSS|anode|cathode|vss \$94578 d|z VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2901875p AD=0.4068p PS=1.55u PD=2.57u
M$1584 VSS|anode|cathode|vss a2|zn$1 \$96154 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$1585 \$96154 a1|z$4 d|zn$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$1586 d|zn$1 b|zn VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$1587 b|zn$1 a1|a2|a3|z \$95723 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$1588 \$95723 GO|a2|core|p2c \$95736 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$1589 \$95736 a2|a3|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$1590 a1|z$1 a1|b|i|q$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$1591 a1|z$2 a1|b|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$1592 \$100313 \$100687 \$100313 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$1604 \$98295 z$6 \$98295 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1605 \$95043 zn$1 \$98295 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1606 \$95043 z$6 \$95043 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$1621 \$98296 zn$1 \$95043 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1622 \$98296 z$6 \$98296 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1637 \$98297 zn$1 \$95043 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$1638 \$98297 z$6 \$98297 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$1652 a2 z$4 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u AS=3.2544p
+ AD=3.2544p PS=29.6u PD=29.6u
M$1653 \$95044 z$1 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=11.52u
+ AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$1654 \$95044 z$4 \$95044 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1668 \$95044 z$7 \$95044 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1669 VIP|core|padres z$3 \$95044 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=11.52u AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$1670 VIP|core|padres z$7 VIP|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1684 \$95044 z$2 \$95044 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1685 VIN|core|padres zn \$95044 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=11.52u AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$1686 VIN|core|padres z$2 VIN|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$1736 \$100314 \$100688 \$100314 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=414.72u AS=177.2928p AD=177.2928p PS=941.76u PD=941.76u
M$2024 \$100315 \$100689 \$100315 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$2036 \$98300 z$6 \$98300 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2037 \$95045 zn$1 \$98300 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2038 \$95045 z$6 \$95045 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$2053 \$98301 zn$1 \$95045 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2054 \$98301 z$6 \$98301 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2069 \$98302 zn$1 \$95045 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2070 \$98302 z$6 \$98302 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2072 \$97578 \$97512 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$2073 VSS|anode|cathode|vss cp|z \$97512 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$2074 \$99205 \$99051 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$2075 VSS|anode|cathode|vss cp|z$1 \$99051 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$2076 VSS|anode|cathode|vss \$97512 \$98777 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$2077 \$98777 d|z$1 \$97513 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.42u
+ AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$2078 \$97513 \$97578 \$98778 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$2079 VSS|anode|cathode|vss \$97579 \$98778 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$2080 VSS|anode|cathode|vss \$97513 \$97579 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$2081 \$97579 \$97578 \$98709 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$2082 \$98709 \$97512 \$98776 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$2083 VSS|anode|cathode|vss \$97580 \$98776 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$2084 VSS|anode|cathode|vss \$98709 \$97580 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$2085 \$99052 \$99205 \$99393 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$2086 \$99393 \$99054 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$2087 \$99053 \$99051 \$99382 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$2088 \$99382 \$99206 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$2089 \$99054 \$99205 \$99053 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$2090 VSS|anode|cathode|vss \$99051 \$99390 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$2091 \$99390 d|zn$1 \$99052 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$2092 VSS|anode|cathode|vss \$99052 \$99054 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$2093 VSS|anode|cathode|vss \$99053 \$99206 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$2094 b|i|q$1 \$97580 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$2095 RESULT[3]|c2p|core|i|q \$99206 VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$2456 \$102486 \$102482 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$2457 VSS|anode|cathode|vss cp|z$1 \$102482 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$2458 \$102483 \$102486 \$102749 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$2459 \$102749 \$102487 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$2460 \$102484 \$102482 \$102747 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$2461 \$102747 \$102761 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$2462 \$102487 \$102486 \$102484 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$2463 VSS|anode|cathode|vss \$102482 \$102748 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$2464 \$102748 d|zn$2 \$102483 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$2465 VSS|anode|cathode|vss \$102483 \$102487 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$2466 VSS|anode|cathode|vss \$102484 \$102761 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$2467 RESULT[0]|c2p|core|i|q \$102761 VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$2468 \$104202 z$6 \$104202 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2469 \$100687 zn$1 \$104202 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2470 \$100687 z$6 \$100687 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$2473 \$104203 zn$1 \$100687 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2474 \$104203 z$6 \$104203 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2477 \$104204 zn$1 \$100687 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2478 \$104204 z$6 \$104204 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2504 VREFH|core|padres z$7 VREFH|core|padres VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$2505 \$100688 z$3 VREFH|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$2506 \$100688 z$7 \$100688 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$2508 \$100688 z$9 \$100688 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$2509 a2 z \$100688 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$2510 a2 z$9 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u AS=1.6272p
+ AD=1.6272p PS=14.8u PD=14.8u
M$2512 \$100688 z$8 \$100688 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$2513 a2$1 z$5 \$100688 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$2514 a2$1 z$8 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$2576 \$104207 z$6 \$104207 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2577 \$100689 zn$1 \$104207 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2578 \$100689 z$6 \$100689 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$2581 \$104208 zn$1 \$100689 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2582 \$104208 z$6 \$104208 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2585 \$104209 zn$1 \$100689 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$2586 \$104209 z$6 \$104209 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$2588 VSS|anode|cathode|vss a2|z$2 \$105952 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$2589 \$105952 a1|i|q b|zn VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$2590 b|zn RST|a1|b|cdn|core|i|p2c VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$2591 \$105690 a1|z$3 \$105955 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$2592 \$105955 a2|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.655u AS=0.271825p AD=0.2901875p PS=1.485u PD=1.55u
M$2593 VSS|anode|cathode|vss \$105690 d|z$2 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2901875p AD=0.4068p PS=1.55u PD=2.57u
M$2594 VSS|anode|cathode|vss a2|zn$2 \$105953 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$2595 \$105953 a1|z$5 d|zn$3 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$2596 d|zn$3 b|zn VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$2597 \$105989 \$106438 \$105989 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$2705 \$105990 \$106439 \$105990 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=207.36u AS=88.6464p AD=88.6464p PS=470.88u PD=470.88u
M$2921 \$105991 \$106440 \$105991 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$3317 a1|z$5 RESULT[2]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$3318 b|zn$2 a1|z$7 \$108285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$3319 \$108285 a2|i|q \$108284 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$3320 \$108284 a1|a2|a3|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$3321 \$107306 \$106803 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$3322 VSS|anode|cathode|vss cp|z \$106803 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$3323 VSS|anode|cathode|vss \$106803 \$108289 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$3324 \$108289 d|z \$106804 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.42u
+ AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$3325 \$106804 \$107306 \$108288 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$3326 VSS|anode|cathode|vss \$107307 \$108288 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$3327 VSS|anode|cathode|vss \$106804 \$107307 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$3328 \$107307 \$107306 \$107993 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$3329 \$107993 \$106803 \$108292 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$3330 VSS|anode|cathode|vss \$107783 \$108292 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$3331 VSS|anode|cathode|vss \$107993 \$107783 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$3332 b|i|q \$107783 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$3333 a1|z$6 a1|b|i|q$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$3334 \$110982 \$111646 \$110982 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$3346 \$109162 z$6 \$109162 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3347 \$106438 zn$1 \$109162 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3348 \$106438 z$6 \$106438 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$3363 \$109163 zn$1 \$106438 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3364 \$109163 z$6 \$109163 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3379 \$109164 zn$1 \$106438 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3380 \$109164 z$6 \$109164 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3478 \$110983 \$111647 \$110983 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=103.68u AS=44.3232p AD=44.3232p PS=235.44u PD=235.44u
M$3491 \$106439 z$3 VREFH|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$3492 \$106439 z$7 \$106439 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$3506 \$106439 z$12 \$106439 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$3507 a2 z$11 \$106439 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$3508 a2 z$12 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.44u AS=0.8136p
+ AD=0.8136p PS=7.4u PD=7.4u
M$3522 \$106439 z$10 \$106439 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$3523 a2$1 z$13 \$106439 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$3524 a2$1 z$10 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$3526 \$110984 \$111648 \$110984 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$3574 \$110985 \$111649 \$110985 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$3766 \$110986 \$111650 \$110986 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$3778 \$109165 z$6 \$109165 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3779 \$106440 zn$1 \$109165 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3780 \$106440 z$6 \$106440 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$3795 \$109166 zn$1 \$106440 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3796 \$109166 z$6 \$109166 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3811 \$109167 zn$1 \$106440 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$3812 \$109167 z$6 \$109167 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$3814 \$110275 \$109669 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$3815 VSS|anode|cathode|vss cp|z \$109669 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$3816 VSS|anode|cathode|vss \$109669 \$111386 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$3817 \$111386 d|z$2 \$109670 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$3818 \$109670 \$110275 \$111392 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$3819 VSS|anode|cathode|vss \$109671 \$111392 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$3820 VSS|anode|cathode|vss \$109670 \$109671 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$3821 \$109671 \$110275 \$110890 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$3822 \$110890 \$109669 \$111370 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$3823 VSS|anode|cathode|vss \$110361 \$111370 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$3824 VSS|anode|cathode|vss \$110890 \$110361 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$3825 a1|z$8 RESULT[1]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$3826 \$108729 a2|d|zn d|zn$4 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$3827 d|zn$4 a1|z$9 \$108729 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$3828 \$108729 b|zn$2 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$3829 \$108730 a2|zn$3 d|zn$5 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$3830 d|zn$5 a1|z$6 \$108730 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$3831 \$108730 b|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$3832 b|q \$110361 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$3833 \$108731 i|z$3 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$3834 VSS|anode|cathode|vss \$108731 cp|z VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$4195 a1|a2|a3|z RST|a1|b|cdn|core|i|p2c VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$4196 \$111651 i|z$3 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$4197 VSS|anode|cathode|vss \$111651 cp|z$1 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$4198 \$111966 \$111445 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$4199 VSS|anode|cathode|vss cp|z$1 \$111445 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$4200 \$111446 \$111966 \$111882 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$4201 \$111882 \$111652 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$4202 \$111447 \$111445 \$111883 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$4203 \$111883 \$111967 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$4204 \$111652 \$111966 \$111447 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$4205 VSS|anode|cathode|vss \$111445 \$111968 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$4206 \$111968 d|zn \$111446 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$4207 VSS|anode|cathode|vss \$111446 \$111652 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$4208 VSS|anode|cathode|vss \$111447 \$111967 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$4209 RESULT[4]|c2p|core|i|q \$111967 VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$4210 \$114499 z$6 \$114499 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4211 \$111646 zn$1 \$114499 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4212 \$111646 z$6 \$111646 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$4215 \$114500 zn$1 \$111646 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4216 \$114500 z$6 \$114500 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4219 \$114501 zn$1 \$111646 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4220 \$114501 z$6 \$114501 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4247 \$111647 z$3 VREFH|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$4248 \$111647 z$7 \$111647 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4250 \$111647 z$14 \$111647 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4251 a2 z$15 \$111647 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$4252 a2 z$14 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p
+ AD=0.4068p PS=3.7u PD=3.7u
M$4254 \$111647 z$16 \$111647 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4255 a2$1 z$19 \$111647 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$4256 a2$1 z$16 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4259 \$111648 z$3 VREFH|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4260 \$111648 z$7 \$111648 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4262 \$111648 z$17 \$111648 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4263 a2 z$25 \$111648 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4264 a2 z$17 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p
+ AD=0.2034p PS=1.85u PD=1.85u
M$4266 \$111648 z$21 \$111648 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4267 a2$1 z$23 \$111648 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4268 a2$1 z$21 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4271 \$111649 z$3 VREFH|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4272 \$111649 z$7 \$111649 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4274 \$111649 z$18 \$111649 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4275 a2 zn$2 \$111649 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4276 a2 z$18 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p
+ AD=0.2034p PS=1.85u PD=1.85u
M$4279 a2$1 zn$2 \$111649 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4280 a2$1 z$18 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4318 \$114502 z$6 \$114502 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4319 \$111650 zn$1 \$114502 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4320 \$111650 z$6 \$111650 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$4323 \$114503 zn$1 \$111650 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4324 \$114503 z$6 \$114503 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4327 \$114504 zn$1 \$111650 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$4328 \$114504 z$6 \$114504 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$4330 \$114519 \$114505 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$4331 VSS|anode|cathode|vss cp|z \$114505 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$4332 \$114506 \$114519 \$114826 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$4333 \$114826 \$114520 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$4334 \$114507 \$114505 \$114834 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$4335 \$114834 \$114892 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$4336 \$114520 \$114519 \$114507 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$4337 VSS|anode|cathode|vss \$114505 \$114821 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$4338 \$114821 d|z$3 \$114506 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$4339 VSS|anode|cathode|vss \$114506 \$114520 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$4340 VSS|anode|cathode|vss \$114507 \$114892 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$4341 \$113285 a1|z$7 \$114140 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$4342 VSS|anode|cathode|vss a2|i|q \$114140 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.655u AS=0.2901875p AD=0.271825p PS=1.55u PD=1.485u
M$4343 VSS|anode|cathode|vss \$113285 SAMPLE|a1|c2p|core|i|z
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2901875p AD=0.4068p
+ PS=1.55u PD=2.57u
M$4344 b|i|q$3 \$114892 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$4345 \$116315 \$116455 \$116315 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4381 \$116316 \$116456 \$116316 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4417 \$116317 \$116457 \$116317 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4453 \$116318 \$116458 \$116318 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4489 \$116319 \$116459 \$116319 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4525 \$116320 \$116460 \$116320 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4561 \$116321 \$116461 \$116321 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4597 \$116322 \$116462 \$116322 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4633 \$116323 \$116463 \$116323 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$4669 \$116324 \$116464 \$116324 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$5065 \$119711 z$6 \$119711 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5066 \$116455 zn$1 \$119711 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5067 \$116455 z$6 \$116455 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5070 \$119712 zn$1 \$116455 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5071 \$119712 z$6 \$119712 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5074 \$119713 zn$1 \$116455 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5075 \$119713 z$6 \$119713 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5077 \$119714 z$6 \$119714 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5078 \$116456 zn$1 \$119714 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5079 \$116456 z$6 \$116456 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5082 \$119715 zn$1 \$116456 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5083 \$119715 z$6 \$119715 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5086 \$119716 zn$1 \$116456 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5087 \$119716 z$6 \$119716 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5089 \$119717 z$6 \$119717 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5090 \$116457 zn$1 \$119717 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5091 \$116457 z$6 \$116457 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5094 \$119718 zn$1 \$116457 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5095 \$119718 z$6 \$119718 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5098 \$119719 zn$1 \$116457 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5099 \$119719 z$6 \$119719 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5101 \$119720 z$6 \$119720 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5102 \$116458 zn$1 \$119720 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5103 \$116458 z$6 \$116458 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5106 \$119721 zn$1 \$116458 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5107 \$119721 z$6 \$119721 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5110 \$119722 zn$1 \$116458 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5111 \$119722 z$6 \$119722 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5113 \$119723 z$6 \$119723 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5114 \$116459 zn$1 \$119723 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5115 \$116459 z$6 \$116459 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5118 \$119724 zn$1 \$116459 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5119 \$119724 z$6 \$119724 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5122 \$119725 zn$1 \$116459 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5123 \$119725 z$6 \$119725 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5125 \$119726 z$6 \$119726 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5126 \$116460 zn$1 \$119726 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5127 \$116460 z$6 \$116460 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5130 \$119727 zn$1 \$116460 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5131 \$119727 z$6 \$119727 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5134 \$119728 zn$1 \$116460 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5135 \$119728 z$6 \$119728 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5137 \$119729 z$6 \$119729 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5138 \$116461 zn$1 \$119729 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5139 \$116461 z$6 \$116461 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5142 \$119730 zn$1 \$116461 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5143 \$119730 z$6 \$119730 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5146 \$119731 zn$1 \$116461 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5147 \$119731 z$6 \$119731 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5149 \$119732 z$6 \$119732 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5150 \$116462 zn$1 \$119732 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5151 \$116462 z$6 \$116462 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5154 \$119733 zn$1 \$116462 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5155 \$119733 z$6 \$119733 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5158 \$119734 zn$1 \$116462 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5159 \$119734 z$6 \$119734 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5161 \$119735 z$6 \$119735 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5162 \$116463 zn$1 \$119735 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5163 \$116463 z$6 \$116463 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5166 \$119736 zn$1 \$116463 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5167 \$119736 z$6 \$119736 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5170 \$119737 zn$1 \$116463 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5171 \$119737 z$6 \$119737 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5173 \$119738 z$6 \$119738 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5174 \$116464 zn$1 \$119738 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5175 \$116464 z$6 \$116464 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5178 \$119739 zn$1 \$116464 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5179 \$119739 z$6 \$119739 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5182 \$119740 zn$1 \$116464 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$5183 \$119740 z$6 \$119740 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$5185 \$120649 a1|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$5186 \$120650 a1|i|q \$120651 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2511p AD=0.1494p PS=1.55u PD=1.19u
M$5187 \$120651 \$120649 \$120652 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.1494p AD=0.1494p PS=1.19u PD=1.19u
M$5188 \$120652 \$120650 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.1494p AD=0.2511p PS=1.19u PD=1.55u
M$5189 VSS|anode|cathode|vss a2|i|q \$120650 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.2511p PS=1.55u PD=1.55u
M$5190 VSS|anode|cathode|vss \$120651 a2|a3|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$5191 VSS|anode|cathode|vss i|z$4 \$119240 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.36u AS=0.2511p AD=0.2034p PS=1.55u PD=1.85u
M$5192 VSS|anode|cathode|vss \$119240 i|z$3 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$5193 a2|zn$4 a1|b|i|q$3 \$120592 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5194 \$120592 a1|a2|a3|z \$120593 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5195 \$120593 a2|a3|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5196 a2|z$2 a2|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$5197 a2|z$3 \$120653 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5198 VSS|anode|cathode|vss b|i|q$2 \$120653 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5199 \$120653 a1|b|i|q$1 \$121428 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5200 \$121428 a2|zn$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5201 \$120453 a2|zn$3 d|zn$6 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5202 d|zn$6 a1|z$10 \$120453 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5203 \$120453 b|zn$3 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5204 z$20 i|z$3 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$5205 \$120654 a1|i|q \$121360 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$5206 \$121360 a2|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.655u AS=0.271825p AD=0.2901875p PS=1.485u PD=1.55u
M$5207 VSS|anode|cathode|vss \$120654 VALID|a3|c2p|core|i|z
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2901875p AD=0.4068p
+ PS=1.55u PD=2.57u
M$5208 VSS|anode|cathode|vss i|zn \$124561 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5210 VSS|anode|cathode|vss \$124561 i|z$5 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5214 \$124562 i|z|zn$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5215 VSS|anode|cathode|vss \$123895 \$124563 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5216 \$123895 \$124562 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5217 VSS|anode|cathode|vss \$124563 i|z$1 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5218 VSS|anode|cathode|vss i|z$6 \$124565 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5224 VSS|anode|cathode|vss \$124565 i|z|zn VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5240 VSS|anode|cathode|vss i|z$7 \$124568 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5246 VSS|anode|cathode|vss \$124568 z$21 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5262 VSS|anode|cathode|vss \$124622 i|z$9 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5264 VSS|anode|cathode|vss i|z$8 \$124622 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5265 \$124570 \$123896 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5266 VSS|anode|cathode|vss cp|z$2 \$123896 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5267 \$123897 \$124570 \$124444 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$5268 \$124444 \$123898 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$5269 \$123899 \$123896 \$124458 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$5270 \$124458 \$124571 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$5271 \$123898 \$124570 \$123899 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$5272 VSS|anode|cathode|vss \$123896 \$124608 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$5273 \$124608 d|zn$7 \$123897 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$5274 VSS|anode|cathode|vss \$123897 \$123898 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$5275 VSS|anode|cathode|vss \$123899 \$124571 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$5276 RESULT[1]|c2p|core|i|q \$124571 VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$5277 VSS|anode|cathode|vss i|z$2 \$126395 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5279 VSS|anode|cathode|vss \$126395 i|z$10 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5283 \$126397 i|z$10 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5284 VSS|anode|cathode|vss \$126398 \$126182 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5285 VSS|anode|cathode|vss \$126397 \$126398 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5286 VSS|anode|cathode|vss \$126182 i|z$11 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5287 VSS|anode|cathode|vss \$126830 i|z$109 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5289 VSS|anode|cathode|vss i|z$15 \$126830 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5290 \$126400 i|zn$6 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5296 VSS|anode|cathode|vss \$126400 z$7 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5312 \$126401 i|zn$2 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5318 VSS|anode|cathode|vss \$126401 i|z|zn$1 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5334 \$126403 i|z$16 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5340 VSS|anode|cathode|vss \$126403 z$15 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5356 \$126404 i|zn$8 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5357 VSS|anode|cathode|vss \$126405 \$126183 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5358 VSS|anode|cathode|vss \$126404 \$126405 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5359 VSS|anode|cathode|vss \$126183 i|z$12 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5360 i|zn$1 i|z|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5368 \$126408 i|z$13 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5369 VSS|anode|cathode|vss \$126410 \$126184 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5370 VSS|anode|cathode|vss \$126408 \$126410 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5371 VSS|anode|cathode|vss \$126184 i|z$14 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5372 \$126412 RESULT[1]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p
+ PS=9.3u PD=9.48u
M$5378 VSS|anode|cathode|vss \$126412 i|z|zn$2 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5394 \$126414 i|z|zn$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5395 VSS|anode|cathode|vss \$126415 \$126185 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5396 VSS|anode|cathode|vss \$126414 \$126415 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5397 VSS|anode|cathode|vss \$126185 i|z$81 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5398 \$126417 \$126076 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5399 VSS|anode|cathode|vss cp|z$2 \$126076 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5400 a1|b|i|q$3 \$126418 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$5401 VSS|anode|cathode|vss \$128040 i|z$75 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5403 VSS|anode|cathode|vss i|z \$128040 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5404 i|z|zn$1 i|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5412 VSS|anode|cathode|vss i|z$67 \$127585 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5418 VSS|anode|cathode|vss \$127585 z$3 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5434 \$127586 i|z$17 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5435 VSS|anode|cathode|vss \$127588 \$127589 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5436 \$127588 \$127586 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5437 VSS|anode|cathode|vss \$127589 i|z$18 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5438 VSS|anode|cathode|vss \$128041 i|z$19 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5440 VSS|anode|cathode|vss i|z$27 \$128041 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5441 VSS|anode|cathode|vss \$128043 i|z$20 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5443 VSS|anode|cathode|vss i|z$28 \$128043 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5444 VSS|anode|cathode|vss i|z$21 \$127594 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5450 VSS|anode|cathode|vss \$127594 z$12 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5466 VSS|anode|cathode|vss RESULT[4]|c2p|core|i|q \$127595
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p
+ PS=9.48u PD=9.3u
M$5472 VSS|anode|cathode|vss \$127595 i|z|zn$4 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5488 VSS|anode|cathode|vss i|z$22 \$127598 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5494 VSS|anode|cathode|vss \$127598 a1|i|z|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5510 \$127600 i|z$23 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5511 VSS|anode|cathode|vss \$127602 \$127603 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5512 \$127602 \$127600 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5513 VSS|anode|cathode|vss \$127603 i|z$32 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5514 i|zn$3 i|z|zn$5 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5522 VSS|anode|cathode|vss RESULT[2]|c2p|core|i|q \$127605
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p
+ PS=9.48u PD=9.3u
M$5528 VSS|anode|cathode|vss \$127605 i|z|zn$5 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5544 VSS|anode|cathode|vss i|z$24 \$127608 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5550 VSS|anode|cathode|vss \$127608 z$1 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5566 VSS|anode|cathode|vss \$128046 i|z$106 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5568 VSS|anode|cathode|vss i|z$29 \$128046 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5569 VSS|anode|cathode|vss \$128047 i|z$25 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5571 VSS|anode|cathode|vss i|z$12 \$128047 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5572 VSS|anode|cathode|vss \$128048 i|z$13 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5574 VSS|anode|cathode|vss i|z$30 \$128048 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5575 i|z|zn$6 i|zn$4 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5583 \$127611 i|zn$4 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5584 VSS|anode|cathode|vss \$127612 \$127613 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5585 \$127612 \$127611 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5586 VSS|anode|cathode|vss \$127613 i|z$8 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5587 i|z|zn$3 i|zn$5 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5595 \$127614 i|z$31 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$5596 VSS|anode|cathode|vss \$127614 i|z$26 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$5597 \$127616 CLK|core|i|p2c VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$5598 VSS|anode|cathode|vss \$127616 i|z$4 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$5599 VSS|anode|cathode|vss \$126076 \$127527 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$5600 \$127527 d|zn$8 \$126077 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$5601 \$126077 \$126417 \$127522 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$5602 VSS|anode|cathode|vss \$126186 \$127522 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$5603 VSS|anode|cathode|vss \$126077 \$126186 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$5604 \$126186 \$126417 \$126943 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$5605 \$126943 \$126076 \$127525 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$5606 VSS|anode|cathode|vss \$126418 \$127525 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$5607 VSS|anode|cathode|vss \$126943 \$126418 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$5608 i|zn$5 i|z|zn$3 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5616 i|zn$6 i|z|zn VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5624 VSS|anode|cathode|vss a2|z$5 \$130579 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5625 \$130579 a1|z$12 \$129460 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5626 \$129460 a1|z$12 \$130581 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5627 \$130581 a2|z$5 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5628 VSS|anode|cathode|vss \$129460 i|z$6 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5632 \$129461 i|z$38 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5633 VSS|anode|cathode|vss \$129462 \$129463 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5634 VSS|anode|cathode|vss \$129461 \$129462 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5635 VSS|anode|cathode|vss \$129463 i|z$28 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5636 VSS|anode|cathode|vss \$130202 i|z$33 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5638 VSS|anode|cathode|vss i|z$42 \$130202 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5639 VSS|anode|cathode|vss i|z$43 \$129465 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5641 VSS|anode|cathode|vss \$129465 a2|z$4 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5645 \$129467 i|z|zn$8 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5646 VSS|anode|cathode|vss \$129468 \$129469 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5647 VSS|anode|cathode|vss \$129467 \$129468 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5648 VSS|anode|cathode|vss \$129469 i|z$34 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5649 \$129471 i|z$39 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5650 VSS|anode|cathode|vss \$129472 \$129473 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5651 VSS|anode|cathode|vss \$129471 \$129472 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5652 VSS|anode|cathode|vss \$129473 i|z$35 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5653 VSS|anode|cathode|vss \$130205 i|z$36 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5655 VSS|anode|cathode|vss i|z$44 \$130205 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5656 \$129476 i|z$45 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5662 VSS|anode|cathode|vss \$129476 z$9 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5678 \$129477 i|z$46 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5684 VSS|anode|cathode|vss \$129477 z VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5700 \$129478 i|z|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=1.925u AS=0.942125p AD=0.834125p PS=5.67u PD=4.65u
M$5703 VSS|anode|cathode|vss \$129478 i|z$24 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.3904p AD=2.4984p PS=12.4u PD=13.42u
M$5711 \$129479 i|z$5 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5717 VSS|anode|cathode|vss \$129479 a1|z$11 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5733 \$129481 i|z$47 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5739 VSS|anode|cathode|vss \$129481 z$13 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5755 \$129482 i|z$25 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5756 VSS|anode|cathode|vss \$129483 \$129484 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5757 VSS|anode|cathode|vss \$129482 \$129483 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5758 VSS|anode|cathode|vss \$129484 i|z$30 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5759 i|z|zn$2 i|zn$8 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5767 \$129485 i|z$48 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$5773 VSS|anode|cathode|vss \$129485 z$14 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5789 \$129486 a2|i|z VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5790 VSS|anode|cathode|vss \$129487 \$129488 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5791 VSS|anode|cathode|vss \$129486 \$129487 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5792 VSS|anode|cathode|vss \$129488 i|z$2 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5793 \$129489 i|z$113 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5794 VSS|anode|cathode|vss \$129490 \$129491 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5795 VSS|anode|cathode|vss \$129489 \$129490 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5796 VSS|anode|cathode|vss \$129491 i|z$29 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5797 \$130446 \$130446 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$5798 i|zn$4 i|z|zn$6 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5806 i|z|zn$5 i|zn$3 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5814 i|zn$7 i|zn$2 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5822 \$129493 i|z$59 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5823 VSS|anode|cathode|vss \$129494 \$129495 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5824 VSS|anode|cathode|vss \$129493 \$129494 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$5825 VSS|anode|cathode|vss \$129495 i|z$37 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5826 VSS|anode|cathode|vss \$130212 i|z$7 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5828 VSS|anode|cathode|vss i|z$14 \$130212 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5829 \$129497 RESULT[3]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p
+ PS=9.3u PD=9.48u
M$5835 VSS|anode|cathode|vss \$129497 i|z|zn$7 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5851 a2|zn a1|i|q$1 \$130564 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5852 \$130564 a1|a2|a3|z \$130566 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5853 \$130566 a2|a3|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5854 VSS|anode|cathode|vss cp|i|z \$129355 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.36u AS=0.2511p AD=0.2034p PS=1.55u PD=1.85u
M$5855 VSS|anode|cathode|vss \$129355 cp|z$2 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$5856 a2 z$7 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u AS=0.6102p
+ AD=0.6102p PS=5.55u PD=5.55u
M$5857 a2$1 z$3 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.16u
+ AS=1.2204p AD=1.2204p PS=11.1u PD=11.1u
M$5858 a2$1 z$7 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.08u
+ AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$5868 a1|c|i|zn a2$1 \$130766 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5872 a1|c|i|zn a1|z$11 \$130766 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5876 \$130767 a2|b|z \$130766 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5880 \$130767 a1|c|i|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5884 a1|c|i|zn a2$1 \$130768 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5888 a1|c|i|zn a1|z$11 \$130768 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5892 \$130769 a2|b|z \$130768 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5896 \$130769 a1|c|i|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5900 a1|c|i|zn a2$1 \$130770 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5904 a1|c|i|zn a1|z$11 \$130770 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5908 \$130771 a2|b|z \$130770 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5912 \$130771 a1|c|i|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5916 a1|c|i|zn a2$1 \$130772 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5920 a1|c|i|zn a1|z$11 \$130772 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5924 \$130773 a2|b|z \$130772 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$5928 \$130773 a1|c|i|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$5932 VSS|anode|cathode|vss a2|b|z \$131267 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5933 \$131267 a1|c|i|zn a1|c|i|zn$1 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5934 a1|c|i|zn$1 a1|c|i|zn \$131266 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$5935 \$131266 a2|b|z VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5936 \$130774 a1|c|i|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.154925p AD=0.1105875p PS=1.73u PD=1.13u
M$5937 VSS|anode|cathode|vss \$130774 i|z$55 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1105875p AD=0.15625p PS=1.13u PD=1.73u
M$5938 VSS|anode|cathode|vss \$131123 z$22 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$5940 VSS|anode|cathode|vss i|z$55 \$131123 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5941 \$130777 i|z$33 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5942 VSS|anode|cathode|vss \$130749 \$130778 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5943 \$130749 \$130777 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5944 VSS|anode|cathode|vss \$130778 i|z$27 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5945 VSS|anode|cathode|vss i|z$40 \$130779 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5951 VSS|anode|cathode|vss \$130779 z$23 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$5967 \$130781 i|zn$11 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$5968 VSS|anode|cathode|vss \$130750 \$130782 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$5969 \$130750 \$130781 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$5970 VSS|anode|cathode|vss \$130782 i|z$56 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$5971 i|zn$8 i|z|zn$2 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$5979 VSS|anode|cathode|vss i|z$49 \$130784 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$5985 VSS|anode|cathode|vss \$130784 z$17 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6001 \$130785 i|z$51 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6002 VSS|anode|cathode|vss \$130751 \$130786 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6003 \$130751 \$130785 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6004 VSS|anode|cathode|vss \$130786 i|z$62 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6005 VSS|anode|cathode|vss i|z$24 \$130787 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6011 VSS|anode|cathode|vss \$130787 z$1 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6027 \$130788 i|z$36 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6028 VSS|anode|cathode|vss \$130752 \$130789 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6029 \$130752 \$130788 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6030 VSS|anode|cathode|vss \$130789 i|z$52 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6031 \$130790 i|z$53 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6032 VSS|anode|cathode|vss \$130754 \$130791 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6033 \$130754 \$130790 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6034 VSS|anode|cathode|vss \$130791 i|z$57 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6035 VSS|anode|cathode|vss VALID|a3|c2p|core|i|z i|zn$9 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.3032p AD=1.3032p PS=7.22u PD=7.22u
M$6039 VSS|anode|cathode|vss a2|i|z i|zn$9 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.3032p AD=1.3032p PS=7.22u PD=7.22u
M$6043 VSS|anode|cathode|vss SAMPLE|a1|c2p|core|i|z i|zn$9
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u AS=1.3032p AD=1.3032p
+ PS=7.22u PD=7.22u
M$6047 a1|i|z|zn i|zn VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=4.32u AS=1.9008p AD=1.9008p PS=10.32u PD=10.32u
M$6053 \$130755 \$130755 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6054 i|zn$10 i|z|zn$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6062 \$130795 i|z|zn$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6063 VSS|anode|cathode|vss \$130756 \$130796 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6064 \$130756 \$130795 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6065 VSS|anode|cathode|vss \$130796 i|z$42 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6066 VSS|anode|cathode|vss \$131124 i|z$58 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6068 VSS|anode|cathode|vss i|z$35 \$131124 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6069 VSS|anode|cathode|vss \$131125 i|z$59 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6071 VSS|anode|cathode|vss i|z$1 \$131125 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6072 VSS|anode|cathode|vss \$131126 i|z$48 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6074 VSS|anode|cathode|vss i|z$57 \$131126 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6075 \$130799 i|z|zn$6 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6076 VSS|anode|cathode|vss \$130757 \$130800 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6077 \$130757 \$130799 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6078 VSS|anode|cathode|vss \$130800 i|z$114 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6079 \$130801 i|z$54 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6080 VSS|anode|cathode|vss \$130759 \$130802 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6081 \$130759 \$130801 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6082 VSS|anode|cathode|vss \$130802 i|z VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6083 zn$5 \$131519 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6084 \$130803 i|z$41 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6085 VSS|anode|cathode|vss \$130760 \$130804 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6086 \$130760 \$130803 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6087 VSS|anode|cathode|vss \$130804 i|z$60 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6088 VSS|anode|cathode|vss i|zn$9 \$130806 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.925u AS=0.942125p AD=0.834125p PS=5.67u PD=4.65u
M$6091 VSS|anode|cathode|vss \$130806 i|z$22 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.3904p AD=2.4984p PS=12.4u PD=13.42u
M$6099 VSS|anode|cathode|vss \$131127 i|z$54 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6101 VSS|anode|cathode|vss i|z$37 \$131127 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6102 i|zn$2 SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p
+ PS=13.42u PD=13.42u
M$6110 VSS|anode|cathode|vss i|z$11 \$130807 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6112 VSS|anode|cathode|vss \$130807 i|z$23 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6116 VSS|anode|cathode|vss i|z$26 \$130808 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6122 VSS|anode|cathode|vss \$130808 a2|i|z VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6138 \$130809 CLK|core|i|p2c VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$6139 VSS|anode|cathode|vss \$130809 i|z$61 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$6140 \$130811 i|z$61 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$6141 VSS|anode|cathode|vss \$130811 i|z$31 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$6142 a2|z$1 \$131128 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6143 VSS|anode|cathode|vss b|q \$131128 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6144 \$131128 a1|b|i|q$2 \$131256 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6145 \$131256 a2|zn$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6146 \$130812 \$130761 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6147 VSS|anode|cathode|vss cp|z$2 \$130761 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6148 \$130762 \$130812 \$131099 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$6149 \$131099 \$130813 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$6150 \$130763 \$130761 \$131091 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$6151 \$131091 \$131129 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$6152 \$130813 \$130812 \$130763 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$6153 VSS|anode|cathode|vss \$130761 \$131098 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$6154 \$131098 d|zn$3 \$130762 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$6155 VSS|anode|cathode|vss \$130762 \$130813 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$6156 VSS|anode|cathode|vss \$130763 \$131129 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$6157 RESULT[2]|c2p|core|i|q \$131129 VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$6158 a1|c|i|zn$1 a2 \$133348 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6162 a1|c|i|zn$1 a1|z$11 \$133348 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6166 \$133211 a2|b|z \$133348 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6170 \$133211 a1|c|i|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6174 a1|c|i|zn$1 a2 \$133349 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6178 a1|c|i|zn$1 a1|z$11 \$133349 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6182 \$133212 a2|b|z \$133349 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6186 \$133212 a1|c|i|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6190 a1|c|i|zn$1 a2 \$133350 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6194 a1|c|i|zn$1 a1|z$11 \$133350 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6198 \$133213 a2|b|z \$133350 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6202 \$133213 a1|c|i|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6206 a1|c|i|zn$1 a2 \$133351 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6210 a1|c|i|zn$1 a1|z$11 \$133351 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6214 \$133214 a2|b|z \$133351 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=2.88u AS=1.3032p AD=1.1952p PS=7.22u PD=6.2u
M$6218 \$133214 a1|c|i|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6222 VSS|anode|cathode|vss a2|b|z \$133621 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6223 \$133621 a1|c|i|zn$1 a1|c|i|zn VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6224 a1|c|i|zn a1|c|i|zn$1 \$133620 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6225 \$133620 a2|b|z VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6226 VSS|anode|cathode|vss \$133160 a2|a3|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6228 VSS|anode|cathode|vss i|z$65 \$133160 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6229 VSS|anode|cathode|vss a2|z$4 \$133623 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6230 \$133623 a1|i|z|zn \$132456 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6231 \$132456 a1|i|z|zn \$133628 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6232 \$133628 a2|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6233 VSS|anode|cathode|vss \$132456 i|z$66 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6237 \$132458 i|z$74 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6243 VSS|anode|cathode|vss \$132458 z$11 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6259 \$133352 \$133352 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6260 i|z|zn$7 i|zn$10 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6268 \$132459 i|z$75 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6274 VSS|anode|cathode|vss \$132459 z$25 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6290 \$132461 i|z|zn VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.925u AS=0.942125p AD=0.834125p PS=5.67u PD=4.65u
M$6293 VSS|anode|cathode|vss \$132461 i|z$67 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.3904p AD=2.4984p PS=12.4u PD=13.42u
M$6301 \$132463 i|z|zn$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6302 VSS|anode|cathode|vss \$132464 \$132465 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6303 VSS|anode|cathode|vss \$132463 \$132464 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6304 VSS|anode|cathode|vss \$132465 i|z$63 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6305 \$132466 i|z$76 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6311 VSS|anode|cathode|vss \$132466 z$10 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6327 \$132467 i|z$58 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6333 VSS|anode|cathode|vss \$132467 z$19 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6349 VSS|anode|cathode|vss \$133164 i|z$74 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6351 VSS|anode|cathode|vss i|z$101 \$133164 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6352 \$132468 i|zn$10 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6353 VSS|anode|cathode|vss \$132469 \$132470 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6354 VSS|anode|cathode|vss \$132468 \$132469 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6355 VSS|anode|cathode|vss \$132470 i|z$68 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6356 i|zn$11 i|z|zn$8 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6364 \$133354 \$133354 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6365 \$132473 b|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6371 VSS|anode|cathode|vss \$132473 i|z|zn$8 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6387 VSS|anode|cathode|vss \$133168 i|z$69 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6389 VSS|anode|cathode|vss i|z$77 \$133168 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6390 \$132475 i|z$72 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6391 VSS|anode|cathode|vss \$132476 \$132477 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6392 VSS|anode|cathode|vss \$132475 \$132476 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6393 VSS|anode|cathode|vss \$132477 i|z$64 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6394 \$132478 i|z$69 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6395 VSS|anode|cathode|vss \$132479 \$132480 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6396 VSS|anode|cathode|vss \$132478 \$132479 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6397 VSS|anode|cathode|vss \$132480 i|z$70 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6398 VSS|anode|cathode|vss \$133170 i|z$46 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6400 VSS|anode|cathode|vss i|z$79 \$133170 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6401 \$132482 i|z$103 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6402 VSS|anode|cathode|vss \$132483 \$132484 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6403 VSS|anode|cathode|vss \$132482 \$132483 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6404 VSS|anode|cathode|vss \$132484 i|z$112 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6405 \$132485 i|z$73 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6406 VSS|anode|cathode|vss \$132486 \$132487 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6407 VSS|anode|cathode|vss \$132485 \$132486 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6408 VSS|anode|cathode|vss \$132487 i|z$71 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6409 VSS|anode|cathode|vss \$133171 i|z$16 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6411 VSS|anode|cathode|vss i|z$80 \$133171 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6412 \$132489 b|i|q$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6418 VSS|anode|cathode|vss \$132489 i|z|zn$9 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6434 \$132491 \$132446 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6435 VSS|anode|cathode|vss cp|z$1 \$132446 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6436 a1|i|q$1 \$132493 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6437 \$133781 \$133781 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6438 zn$3 \$134212 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6439 i|z|zn i|zn$6 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6447 VSS|anode|cathode|vss i|z$66 \$133929 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6453 VSS|anode|cathode|vss \$133929 a2|b|z VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6469 zn \$134213 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6470 \$133930 i|z$83 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6471 VSS|anode|cathode|vss \$133783 \$133931 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6472 \$133783 \$133930 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6473 VSS|anode|cathode|vss \$133931 i|z$86 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6474 VSS|anode|cathode|vss i|zn$7 \$133933 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.925u AS=0.942125p AD=0.834125p PS=5.67u PD=4.65u
M$6477 VSS|anode|cathode|vss \$133933 a1|z$12 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.3904p AD=2.4984p PS=12.4u PD=13.42u
M$6485 VSS|anode|cathode|vss \$133935 i|z$83 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6487 VSS|anode|cathode|vss i|z$97 \$133935 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6488 VSS|anode|cathode|vss \$133936 i|z$87 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6490 VSS|anode|cathode|vss i|z$102 \$133936 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6491 \$133938 a1|i|z|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6492 VSS|anode|cathode|vss \$133784 \$133939 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6493 \$133784 \$133938 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6494 VSS|anode|cathode|vss \$133939 i|z$43 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6495 \$132448 a1|c|i|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.154925p AD=0.1105875p PS=1.73u PD=1.13u
M$6496 VSS|anode|cathode|vss \$132448 i|z$65 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.25u AS=0.1105875p AD=0.15625p PS=1.13u PD=1.73u
M$6497 VSS|anode|cathode|vss i|z$98 \$133940 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6503 VSS|anode|cathode|vss \$133940 z$8 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6519 \$133941 i|z$84 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6520 VSS|anode|cathode|vss \$133786 \$133942 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6521 \$133786 \$133941 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6522 VSS|anode|cathode|vss \$133942 i|z$80 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6523 \$133943 i|zn$3 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6524 VSS|anode|cathode|vss \$133787 \$133944 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6525 \$133787 \$133943 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6526 VSS|anode|cathode|vss \$133944 i|z$88 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6527 VSS|anode|cathode|vss \$133946 i|z$82 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6529 VSS|anode|cathode|vss i|z$89 \$133946 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6530 i|zn$12 i|z|zn$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6538 VSS|anode|cathode|vss i|z$32 \$133949 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6540 VSS|anode|cathode|vss \$133949 a2|z$5 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.1952p AD=1.3032p PS=6.2u PD=7.22u
M$6544 i|zn a1|i|z|zn VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=4.32u AS=1.9008p AD=1.9008p PS=10.32u PD=10.32u
M$6550 VSS|anode|cathode|vss \$133950 i|z$17 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6552 VSS|anode|cathode|vss i|z$81 \$133950 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6553 \$133951 i|z$50 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6554 VSS|anode|cathode|vss \$133788 \$133952 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6555 \$133788 \$133951 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6556 VSS|anode|cathode|vss \$133952 i|z$79 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6557 VSS|anode|cathode|vss i|z$87 \$133953 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6563 VSS|anode|cathode|vss \$133953 z$16 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6579 VSS|anode|cathode|vss \$133954 i|z$39 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6581 VSS|anode|cathode|vss i|z$18 \$133954 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6582 VSS|anode|cathode|vss \$133955 i|z$41 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6584 VSS|anode|cathode|vss i|z$34 \$133955 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6585 VSS|anode|cathode|vss i|z$78 \$133956 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6591 VSS|anode|cathode|vss \$133956 z$5 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6607 VSS|anode|cathode|vss \$133957 i|z$45 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6609 VSS|anode|cathode|vss i|z$90 \$133957 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6610 VSS|anode|cathode|vss \$133959 i|z$91 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6612 VSS|anode|cathode|vss i|z$92 \$133959 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6613 VSS|anode|cathode|vss \$133962 i|z$98 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6615 VSS|anode|cathode|vss i|z$99 \$133962 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6616 VSS|anode|cathode|vss b|i|q$2 \$133964 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6622 VSS|anode|cathode|vss \$133964 i|z|zn$6 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6638 \$133965 i|z|zn$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6639 VSS|anode|cathode|vss \$133789 \$133966 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6640 \$133789 \$133965 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6641 VSS|anode|cathode|vss \$133966 i|z$89 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6642 \$133967 i|z$85 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6643 VSS|anode|cathode|vss \$133791 \$133968 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6644 \$133791 \$133967 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6645 VSS|anode|cathode|vss \$133968 i|z$93 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6646 VSS|anode|cathode|vss \$133970 i|z$49 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6648 VSS|anode|cathode|vss i|z$70 \$133970 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6649 \$133971 i|z$82 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6650 VSS|anode|cathode|vss \$133792 \$133972 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6651 \$133792 \$133971 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6652 VSS|anode|cathode|vss \$133972 i|z$94 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6653 VSS|anode|cathode|vss \$133974 i|z$85 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6655 VSS|anode|cathode|vss i|z$71 \$133974 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6656 i|z|zn$9 i|zn$13 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6664 \$133976 i|z$107 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6665 VSS|anode|cathode|vss \$133793 \$133977 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6666 \$133793 \$133976 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6667 VSS|anode|cathode|vss \$133977 i|z$100 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6668 \$133978 i|zn$12 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6669 VSS|anode|cathode|vss \$133794 \$133979 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6670 \$133794 \$133978 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6671 VSS|anode|cathode|vss \$133979 i|z$95 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6672 VSS|anode|cathode|vss \$133982 i|z$51 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6674 VSS|anode|cathode|vss i|z$96 \$133982 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6675 VSS|anode|cathode|vss \$133983 i|z$72 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6677 VSS|anode|cathode|vss i|z$95 \$133983 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6678 VSS|anode|cathode|vss \$132446 \$133732 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$6679 \$133732 d|zn$4 \$132447 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$6680 \$132447 \$132491 \$133726 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$6681 VSS|anode|cathode|vss \$132492 \$133726 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$6682 VSS|anode|cathode|vss \$132447 \$132492 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$6683 \$132492 \$132491 \$133356 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$6684 \$133356 \$132446 \$133730 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$6685 VSS|anode|cathode|vss \$132493 \$133730 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$6686 VSS|anode|cathode|vss \$133356 \$132493 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$6687 \$133804 a2|a3|zn b|zn$4 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6688 b|zn$4 RST|a1|b|cdn|core|i|p2c \$133804 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6689 \$133804 a1|b|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6690 \$133805 i|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$6691 VSS|anode|cathode|vss \$133805 cp|i|z VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$6692 \$135445 i|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6698 VSS|anode|cathode|vss \$135445 z$4 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6714 \$135446 i|z$9 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6715 VSS|anode|cathode|vss \$135447 \$135382 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6716 VSS|anode|cathode|vss \$135446 \$135447 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6717 VSS|anode|cathode|vss \$135382 i|z$97 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6718 VSS|anode|cathode|vss \$136356 i|z$50 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6720 VSS|anode|cathode|vss i|z$62 \$136356 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6721 zn$4 \$135448 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6722 \$135449 i|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6728 VSS|anode|cathode|vss \$135449 z$4 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6744 VSS|anode|cathode|vss \$136357 i|z$21 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6746 VSS|anode|cathode|vss i|z$86 \$136357 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6747 \$135450 i|z|zn$9 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6748 VSS|anode|cathode|vss \$135451 \$135383 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6749 VSS|anode|cathode|vss \$135450 \$135451 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6750 VSS|anode|cathode|vss \$135383 i|z$96 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6751 \$135452 b|i|q$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=3.85u AS=1.66825p AD=1.65025p PS=9.3u PD=9.48u
M$6757 VSS|anode|cathode|vss \$135452 i|z|zn$3 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6773 \$135453 i|z$19 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6774 VSS|anode|cathode|vss \$135454 \$135384 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6775 VSS|anode|cathode|vss \$135453 \$135454 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6776 VSS|anode|cathode|vss \$135384 i|z$105 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6777 \$135456 i|z$106 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6778 VSS|anode|cathode|vss \$135458 \$135385 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6779 VSS|anode|cathode|vss \$135456 \$135458 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6780 VSS|anode|cathode|vss \$135385 i|z$101 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6781 VSS|anode|cathode|vss \$136358 i|z$103 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6783 VSS|anode|cathode|vss i|z$56 \$136358 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6784 \$136577 \$136577 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6785 VSS|anode|cathode|vss \$136359 i|z$38 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6787 VSS|anode|cathode|vss i|z$88 \$136359 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6788 i|zn$13 i|z|zn$9 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6796 VSS|anode|cathode|vss \$136360 i|z$107 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6798 VSS|anode|cathode|vss i|z$94 \$136360 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6799 zn$2 \$135460 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6800 \$135461 i|z$108 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6801 VSS|anode|cathode|vss \$135463 \$135386 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6802 VSS|anode|cathode|vss \$135461 \$135463 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6803 VSS|anode|cathode|vss \$135386 i|z$99 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6804 \$135464 i|z$109 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6805 VSS|anode|cathode|vss \$135466 \$135387 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6806 VSS|anode|cathode|vss \$135464 \$135466 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6807 VSS|anode|cathode|vss \$135387 i|z$77 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6808 i|z|zn$4 i|zn$12 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6816 VSS|anode|cathode|vss \$136361 i|z$110 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6818 VSS|anode|cathode|vss i|z$104 \$136361 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6819 i|z|zn$8 i|zn$11 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=2.4984p AD=2.4984p PS=13.42u PD=13.42u
M$6827 VSS|anode|cathode|vss \$136362 i|z$73 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6829 VSS|anode|cathode|vss i|z$68 \$136362 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6830 VSS|anode|cathode|vss \$136363 i|z$108 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6832 VSS|anode|cathode|vss i|z$64 \$136363 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6833 \$135468 i|z$110 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6834 VSS|anode|cathode|vss \$135469 \$135388 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6835 VSS|anode|cathode|vss \$135468 \$135469 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6836 VSS|anode|cathode|vss \$135388 i|z$92 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6837 \$135470 i|z$91 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6838 VSS|anode|cathode|vss \$135471 \$135389 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6839 VSS|anode|cathode|vss \$135470 \$135471 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6840 VSS|anode|cathode|vss \$135389 i|z$90 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6841 VSS|anode|cathode|vss \$136364 i|z$84 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6843 VSS|anode|cathode|vss i|z$60 \$136364 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6844 VSS|anode|cathode|vss \$136365 i|z$40 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6846 VSS|anode|cathode|vss i|z$105 \$136365 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6847 VSS|anode|cathode|vss \$136366 i|z$76 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6849 VSS|anode|cathode|vss i|z$93 \$136366 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6850 \$135472 i|z$20 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6851 VSS|anode|cathode|vss \$135473 \$135390 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6852 VSS|anode|cathode|vss \$135472 \$135473 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6853 VSS|anode|cathode|vss \$135390 i|z$102 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6854 \$135474 i|z$111 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6855 VSS|anode|cathode|vss \$135475 \$135391 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6856 VSS|anode|cathode|vss \$135474 \$135475 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6857 VSS|anode|cathode|vss \$135391 i|z$44 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6858 VSS|anode|cathode|vss \$136367 i|z$47 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6860 VSS|anode|cathode|vss i|z$100 \$136367 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6861 \$135476 i|zn$13 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6862 VSS|anode|cathode|vss \$135477 \$135392 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6863 VSS|anode|cathode|vss \$135476 \$135477 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.267p AD=0.2712p PS=1.55u PD=2.09u
M$6864 VSS|anode|cathode|vss \$135392 i|z$104 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6865 VSS|anode|cathode|vss \$136368 i|z$78 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6867 VSS|anode|cathode|vss i|z$52 \$136368 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6868 \$135478 \$135241 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6869 VSS|anode|cathode|vss cp|z$2 \$135241 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6870 a1|b|i|q$2 \$135479 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6871 VSS|anode|cathode|vss a2|zn$6 \$136799 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6872 \$136799 a1|z$13 d|zn$2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$6873 d|zn$2 b|zn VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6874 zn$1 \$137560 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6875 \$136908 i|zn$5 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6876 VSS|anode|cathode|vss \$136862 \$136909 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6877 \$136862 \$136908 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.48u AS=0.2712p AD=0.267p PS=2.09u PD=1.55u
M$6878 VSS|anode|cathode|vss \$136909 i|z$15 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.267p AD=0.4068p PS=1.55u PD=2.57u
M$6879 VSS|anode|cathode|vss i|zn$6 \$136910 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6885 VSS|anode|cathode|vss \$136910 z$7 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6901 VSS|anode|cathode|vss i|z$67 \$136911 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=3.85u AS=1.587975p AD=1.730525p PS=9.48u PD=9.3u
M$6907 VSS|anode|cathode|vss \$136911 z$3 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=11.52u AS=4.7808p AD=4.8888p PS=24.8u PD=25.82u
M$6923 VSS|anode|cathode|vss \$136912 i|z$113 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6925 VSS|anode|cathode|vss i|z$114 \$136912 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6926 VSS|anode|cathode|vss \$136915 i|z$53 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6928 VSS|anode|cathode|vss i|z$112 \$136915 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6929 VSS|anode|cathode|vss \$136916 i|z$111 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=1.44u AS=0.7056p AD=0.5976p PS=4.12u PD=3.1u
M$6931 VSS|anode|cathode|vss i|z$63 \$136916 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6932 \$136917 \$136863 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6933 VSS|anode|cathode|vss cp|i|z \$136863 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6934 \$136864 \$136917 \$137532 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$6935 \$137532 \$136918 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$6936 \$136865 \$136863 \$137518 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$6937 \$137518 \$136919 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$6938 \$136918 \$136917 \$136865 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$6939 VSS|anode|cathode|vss \$136863 \$137527 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$6940 \$137527 d|zn$9 \$136864 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$6941 VSS|anode|cathode|vss \$136864 \$136918 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$6942 VSS|anode|cathode|vss \$136865 \$136919 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$6943 VSS|anode|cathode|vss \$135241 \$136814 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$6944 \$136814 d|zn$6 \$135242 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$6945 \$135242 \$135478 \$136816 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$6946 VSS|anode|cathode|vss \$135393 \$136816 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$6947 VSS|anode|cathode|vss \$135242 \$135393 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$6948 \$135393 \$135478 \$136579 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$6949 \$136579 \$135241 \$136792 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$6950 VSS|anode|cathode|vss \$135479 \$136792 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$6951 VSS|anode|cathode|vss \$136579 \$135479 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$6952 a1|b|i|q$1 \$136919 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6953 \$136920 \$136866 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$6954 VSS|anode|cathode|vss cp|z$3 \$136866 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$6955 \$136867 \$136920 \$137507 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$6956 \$137507 \$136921 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$6957 \$136868 \$136866 \$137497 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$6958 \$137497 \$136922 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$6959 \$136921 \$136920 \$136868 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$6960 VSS|anode|cathode|vss \$136866 \$137505 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$6961 \$137505 d|zn$10 \$136867 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$6962 VSS|anode|cathode|vss \$136867 \$136921 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$6963 VSS|anode|cathode|vss \$136868 \$136922 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$6964 a1|b|i|q \$136922 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$6965 \$140500 \$140555 \$140500 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7001 \$140501 \$140556 \$140501 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7037 \$140502 \$140557 \$140502 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7073 \$140503 \$140558 \$140503 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7109 \$140504 \$140559 \$140504 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7145 \$140505 \$140560 \$140505 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7181 \$140506 \$140561 \$140506 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7217 \$140507 \$140562 \$140507 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7253 \$140508 \$140563 \$140508 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7289 \$140509 \$140564 \$140509 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7325 \$140565 a1|z$3 \$140949 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$7326 \$140949 a2|z$6 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.655u AS=0.271825p AD=0.2901875p PS=1.485u PD=1.55u
M$7327 VSS|anode|cathode|vss \$140565 d|z$1 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2901875p AD=0.4068p PS=1.55u PD=2.57u
M$7328 a2|zn$6 a1|b|i|q$2 \$139980 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$7329 \$139980 a1|a2|a3|z \$139955 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$7330 \$139955 a2|a3|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$7691 \$142237 \$141920 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$7692 VSS|anode|cathode|vss cp|z$3 \$141920 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$7693 a2|i|q \$142239 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$7694 a2|z \$142241 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$7695 VSS|anode|cathode|vss b|i|q \$142241 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$7696 \$142241 a1|b|i|q \$143472 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$7697 \$143472 a2|zn$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$7698 \$143729 z$26 \$143729 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7699 \$140555 zn$3 \$143729 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7700 \$140555 z$26 \$140555 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7703 \$143730 zn$3 \$140555 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7704 \$143730 z$26 \$143730 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7707 \$143731 zn$3 \$140555 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7708 \$143731 z$26 \$143731 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7710 \$143732 z$26 \$143732 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7711 \$140556 zn$3 \$143732 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7712 \$140556 z$26 \$140556 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7715 \$143733 zn$3 \$140556 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7716 \$143733 z$26 \$143733 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7719 \$143734 zn$3 \$140556 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7720 \$143734 z$26 \$143734 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7722 \$143735 z$26 \$143735 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7723 \$140557 zn$3 \$143735 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7724 \$140557 z$26 \$140557 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7727 \$143736 zn$3 \$140557 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7728 \$143736 z$26 \$143736 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7731 \$143737 zn$3 \$140557 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7732 \$143737 z$26 \$143737 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7734 \$143738 z$26 \$143738 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7735 \$140558 zn$3 \$143738 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7736 \$140558 z$26 \$140558 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7739 \$143739 zn$3 \$140558 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7740 \$143739 z$26 \$143739 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7743 \$143740 zn$3 \$140558 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7744 \$143740 z$26 \$143740 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7746 \$143741 z$26 \$143741 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7747 \$140559 zn$3 \$143741 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7748 \$140559 z$26 \$140559 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7751 \$143742 zn$3 \$140559 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7752 \$143742 z$26 \$143742 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7755 \$143743 zn$3 \$140559 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7756 \$143743 z$26 \$143743 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7758 \$143744 z$26 \$143744 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7759 \$140560 zn$3 \$143744 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7760 \$140560 z$26 \$140560 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7763 \$143745 zn$3 \$140560 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7764 \$143745 z$26 \$143745 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7767 \$143746 zn$3 \$140560 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7768 \$143746 z$26 \$143746 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7770 \$143747 z$26 \$143747 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7771 \$140561 zn$3 \$143747 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7772 \$140561 z$26 \$140561 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7775 \$143748 zn$3 \$140561 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7776 \$143748 z$26 \$143748 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7779 \$143749 zn$3 \$140561 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7780 \$143749 z$26 \$143749 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7782 \$143750 z$26 \$143750 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7783 \$140562 zn$3 \$143750 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7784 \$140562 z$26 \$140562 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7787 \$143751 zn$3 \$140562 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7788 \$143751 z$26 \$143751 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7791 \$143752 zn$3 \$140562 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7792 \$143752 z$26 \$143752 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7794 \$143753 z$26 \$143753 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7795 \$140563 zn$3 \$143753 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7796 \$140563 z$26 \$140563 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7799 \$143754 zn$3 \$140563 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7800 \$143754 z$26 \$143754 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7803 \$143755 zn$3 \$140563 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7804 \$143755 z$26 \$143755 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7806 \$143756 z$26 \$143756 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7807 \$140564 zn$3 \$143756 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7808 \$140564 z$26 \$140564 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$7811 \$143757 zn$3 \$140564 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7812 \$143757 z$26 \$143757 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7815 \$143758 zn$3 \$140564 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$7816 \$143758 z$26 \$143758 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$7818 VSS|anode|cathode|vss \$141920 \$143476 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$7819 \$143476 d|zn$5 \$141921 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$7820 \$141921 \$142237 \$143474 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$7821 VSS|anode|cathode|vss \$142238 \$143474 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$7822 VSS|anode|cathode|vss \$141921 \$142238 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$7823 \$142238 \$142237 \$143400 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$7824 \$143400 \$141920 \$143475 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$7825 VSS|anode|cathode|vss \$142239 \$143475 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$7826 VSS|anode|cathode|vss \$143400 \$142239 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$7827 \$143688 a2|a3|zn b|zn$5 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$7828 b|zn$5 RST|a1|b|cdn|core|i|p2c \$143688 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$7829 \$143688 a1|b|i|q$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$7830 \$145966 \$146281 \$145966 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$7866 \$145967 \$146282 \$145967 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=829.44u AS=354.5856p AD=354.5856p PS=1883.52u PD=1883.52u
M$7902 \$145968 \$146283 \$145968 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=414.72u AS=177.2928p AD=177.2928p PS=941.76u PD=941.76u
M$7938 \$145969 \$146284 \$145969 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=103.68u AS=44.3232p AD=44.3232p PS=235.44u PD=235.44u
M$7974 \$145970 \$146285 \$145970 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$8010 \$145971 \$146286 \$145971 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$8154 \$145972 \$146287 \$145972 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$8550 \$145714 \$144911 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$8551 VSS|anode|cathode|vss cp|z$3 \$144911 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$8552 VSS|anode|cathode|vss \$144911 \$146838 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$8553 \$146838 d|z$4 \$144913 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$8554 \$144913 \$145714 \$146837 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$8555 VSS|anode|cathode|vss \$144914 \$146837 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.1659p AD=0.10375p PS=1.3u PD=1.08u
M$8556 VSS|anode|cathode|vss \$144913 \$144914 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$8557 \$144914 \$145714 \$146288 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$8558 \$146288 \$144911 \$146840 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$8559 VSS|anode|cathode|vss \$146170 \$146840 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.236525p AD=0.10375p PS=1.55u PD=1.08u
M$8560 VSS|anode|cathode|vss \$146288 \$146170 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$8561 a1|z$3 \$146994 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$8562 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$146994
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p
+ PS=1.55u PD=1.55u
M$8563 \$146994 a1|i|q \$147186 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$8564 \$147186 a2|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$8565 \$146995 a1|z$3 \$147184 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$8566 \$147184 a2|z$7 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.655u AS=0.271825p AD=0.2901875p PS=1.485u PD=1.55u
M$8567 VSS|anode|cathode|vss \$146995 d|z$3 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2901875p AD=0.4068p PS=1.55u PD=2.57u
M$8568 b|i|q$2 \$146170 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$8569 \$146996 cp|i|z VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.36u AS=0.2034p AD=0.2511p PS=1.85u PD=1.55u
M$8570 VSS|anode|cathode|vss \$146996 cp|z$3 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2511p AD=0.4068p PS=1.55u PD=2.57u
M$8571 \$149147 z$26 \$149147 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8572 \$146281 zn$3 \$149147 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8573 \$146281 z$26 \$146281 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$8576 \$149148 zn$3 \$146281 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8577 \$149148 z$26 \$149148 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8580 \$149149 zn$3 \$146281 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8581 \$149149 z$26 \$149149 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8583 a2$1 z$4 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8584 \$146282 z$1 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=11.52u
+ AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$8585 \$146282 z$4 \$146282 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8587 \$146282 z$7 \$146282 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8588 VIN|core|padres z$3 \$146282 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=11.52u AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$8589 VIN|core|padres z$7 VIN|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8591 \$146282 z$27 \$146282 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8592 VIP|core|padres zn$5 \$146282 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=11.52u AS=6.5088p AD=6.5088p PS=59.2u PD=59.2u
M$8593 VIP|core|padres z$27 VIP|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8595 VREFL|core|padres z$7 VREFL|core|padres VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8596 \$146283 z$3 VREFL|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=5.76u AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8597 \$146283 z$7 \$146283 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$8599 \$146283 z$9 \$146283 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$8600 a2$1 z \$146283 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8601 a2$1 z$9 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$8603 \$146283 z$8 \$146283 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$8604 a2 z$5 \$146283 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=5.76u
+ AS=3.2544p AD=3.2544p PS=29.6u PD=29.6u
M$8605 a2 z$8 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u AS=1.6272p
+ AD=1.6272p PS=14.8u PD=14.8u
M$8608 \$146284 z$3 VREFL|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$8609 \$146284 z$7 \$146284 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8611 \$146284 z$14 \$146284 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8612 a2$1 z$15 \$146284 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$8613 a2$1 z$14 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8615 \$146284 z$16 \$146284 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8616 a2 z$19 \$146284 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$8617 a2 z$16 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p
+ AD=0.4068p PS=3.7u PD=3.7u
M$8620 \$146285 z$3 VREFL|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8621 \$146285 z$7 \$146285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8623 \$146285 z$17 \$146285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8624 a2$1 z$25 \$146285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8625 a2$1 z$17 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8627 \$146285 z$21 \$146285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8628 a2 z$23 \$146285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8629 a2 z$21 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p
+ AD=0.2034p PS=1.85u PD=1.85u
M$8632 \$146286 z$3 VREFL|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8633 \$146286 z$7 \$146286 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8635 \$146286 z$24 \$146286 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8636 a2$1 zn$4 \$146286 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8637 a2$1 z$24 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u
+ AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8640 a2 zn$4 \$146286 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u
+ AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8641 a2 z$24 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.36u AS=0.2034p
+ AD=0.2034p PS=1.85u PD=1.85u
M$8679 \$149150 z$26 \$149150 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8680 \$146287 zn$3 \$149150 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8681 \$146287 z$26 \$146287 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$8684 \$149151 zn$3 \$146287 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8685 \$149151 z$26 \$149151 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8688 \$149152 zn$3 \$146287 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$8689 \$149152 z$26 \$149152 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$8691 a2|z$6 \$150022 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$8692 VSS|anode|cathode|vss b|i|q$1 \$150022 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$8693 \$150022 a1|i|q$1 \$150057 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$8694 \$150057 a2|zn$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$8695 \$149644 a2|zn$3 d|zn$9 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$8696 d|zn$9 a1|z$9 \$149644 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$8697 \$149644 b|zn$6 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$8698 \$151000 \$151285 \$151000 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$8806 \$151001 \$151286 \$151001 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=207.36u AS=88.6464p AD=88.6464p PS=470.88u PD=470.88u
M$9022 \$151002 \$151287 \$151002 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$9418 \$151288 a1|z$3 \$152559 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.655u AS=0.370075p AD=0.271825p PS=2.44u PD=1.485u
M$9419 VSS|anode|cathode|vss a2|z$3 \$152559 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.655u AS=0.2901875p AD=0.271825p PS=1.55u PD=1.485u
M$9420 VSS|anode|cathode|vss \$151288 d|z$4 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2901875p AD=0.4068p PS=1.55u PD=2.57u
M$9421 \$152828 a2|a3|zn b|zn$6 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$9422 b|zn$6 RST|a1|b|cdn|core|i|p2c \$152828 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9423 \$152828 a1|b|i|q$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$9424 \$154109 z$26 \$154109 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9425 \$151285 zn$3 \$154109 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9426 \$151285 z$26 \$151285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$9429 \$154110 zn$3 \$151285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9430 \$154110 z$26 \$154110 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9433 \$154111 zn$3 \$151285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9434 \$154111 z$26 \$154111 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9461 \$151286 z$3 VREFL|core|padres VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=2.88u AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$9462 \$151286 z$7 \$151286 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$9464 \$151286 z$12 \$151286 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$9465 a2$1 z$11 \$151286 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$9466 a2$1 z$12 a2$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.44u
+ AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$9468 \$151286 z$10 \$151286 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.44u AS=0.8136p AD=0.8136p PS=7.4u PD=7.4u
M$9469 a2 z$13 \$151286 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.88u
+ AS=1.6272p AD=1.6272p PS=14.8u PD=14.8u
M$9470 a2 z$10 a2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=1.44u AS=0.8136p
+ AD=0.8136p PS=7.4u PD=7.4u
M$9532 \$154112 z$26 \$154112 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9533 \$151287 zn$3 \$154112 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9534 \$151287 z$26 \$151287 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$9537 \$154113 zn$3 \$151287 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9538 \$154113 z$26 \$154113 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9541 \$154114 zn$3 \$151287 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$9542 \$154114 z$26 \$154114 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$9544 a1|z$13 RESULT[0]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$9545 a2|z$7 \$155837 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$9546 VSS|anode|cathode|vss b|i|q$3 \$155837 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9547 \$155837 a1|b|i|q$3 \$155910 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9548 \$155910 a2|zn$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$9549 \$155370 a2|zn$3 d|zn$10 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$9550 d|zn$10 a1|z$1 \$155370 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$9551 \$155370 b|zn$4 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$9552 a1|z RESULT[4]|c2p|core|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$9553 VSS|anode|cathode|vss VALID|a3|c2p|core|i|z \$155838
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p
+ PS=2.27u PD=1.83u
M$9554 VSS|anode|cathode|vss \$155838 RD[8]|a4|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$9555 VSS|anode|cathode|vss SAMPLE|a1|c2p|core|i|z \$155840
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p
+ PS=2.27u PD=1.83u
M$9556 VSS|anode|cathode|vss \$155840 RD[9]|a4|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$9557 \$155911 \$156793 \$155911 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$9881 \$155912 \$156794 \$155912 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$10277 a2|zn$1 a1|b|i|q$1 \$158502 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$10278 \$158502 a1|a2|a3|z \$158501 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$10279 \$158501 a2|a3|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$10280 \$159940 z$26 \$159940 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10281 \$156793 zn$3 \$159940 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10282 \$156793 z$26 \$156793 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$10285 \$159941 zn$3 \$156793 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10286 \$159941 z$26 \$159941 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10289 \$159942 zn$3 \$156793 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10290 \$159942 z$26 \$159942 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10388 \$159943 z$26 \$159943 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10389 \$156794 zn$3 \$159943 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10390 \$156794 z$26 \$156794 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$10393 \$159944 zn$3 \$156794 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10394 \$159944 z$26 \$159944 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10397 \$159945 zn$3 \$156794 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$10398 \$159945 z$26 \$159945 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$10400 \$159264 \$158745 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$10401 VSS|anode|cathode|vss cp|z$3 \$158745 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$10402 \$158746 \$159264 \$159266 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.151775p AD=0.10375p PS=1.25u PD=1.08u
M$10403 \$159266 \$158998 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.1659p PS=1.08u PD=1.3u
M$10404 \$158747 \$158745 \$159267 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.25u AS=0.1418875p AD=0.10375p PS=1.215u PD=1.08u
M$10405 \$159267 \$159265 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.25u AS=0.10375p AD=0.236525p PS=1.08u PD=1.55u
M$10406 \$158998 \$159264 \$158747 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.385u AS=0.1837875p AD=0.1418875p PS=1.3u PD=1.215u
M$10407 VSS|anode|cathode|vss \$158745 \$159268 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.42u AS=0.2373p AD=0.1743p PS=1.97u PD=1.25u
M$10408 \$159268 a2|d|zn \$158746 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.42u AS=0.1743p AD=0.151775p PS=1.25u PD=1.25u
M$10409 VSS|anode|cathode|vss \$158746 \$158998 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.47u AS=0.1659p AD=0.1837875p PS=1.3u PD=1.3u
M$10410 VSS|anode|cathode|vss \$158747 \$159265 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.236525p AD=0.4068p PS=1.55u PD=2.57u
M$10411 a2|zn$2 a1|b|i|q \$161717 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$10412 \$161717 a1|a2|a3|z \$161718 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$10413 \$161718 a2|a3|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$10414 a1|i|q \$159265 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$10415 \$161605 \$162307 \$161605 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$10739 \$161606 \$162308 \$161606 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11135 VSS|anode|cathode|vss a2|zn$4 \$162440 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$11136 \$162440 a1|z$8 d|zn$7 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$11137 d|zn$7 b|zn VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$11138 VSS|anode|cathode|vss a2|a3|zn a2|d|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$11139 a2|d|zn RST|a1|b|cdn|core|i|p2c VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p
+ PS=1.55u PD=2.57u
M$11140 \$165672 z$26 \$165672 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11141 \$162307 zn$3 \$165672 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11142 \$162307 z$26 \$162307 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$11145 \$165673 zn$3 \$162307 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11146 \$165673 z$26 \$165673 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11149 \$165674 zn$3 \$162307 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11150 \$165674 z$26 \$165674 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11248 \$165675 z$26 \$165675 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11249 \$162308 zn$3 \$165675 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11250 \$162308 z$26 \$162308 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$11253 \$165676 zn$3 \$162308 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11254 \$165676 z$26 \$165676 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11257 \$165677 zn$3 \$162308 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11258 \$165677 z$26 \$165677 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11260 \$164985 a2|zn$3 d|zn$8 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$11261 d|zn$8 a1|z$2 \$164985 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$11262 \$164985 b|zn$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$11263 a2|zn$3 a1|i|q \$165503 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$11264 \$165503 a2|z$2 \$165502 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$11265 \$165502 a1|a2|a3|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$11266 \$165678 a2|a3|zn b|zn$3 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$11267 b|zn$3 RST|a1|b|cdn|core|i|p2c \$165678 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.2988p PS=1.55u PD=1.55u
M$11268 \$165678 a1|b|i|q$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p PS=1.55u PD=2.57u
M$11269 a1|z$7 a1|i|q VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$11270 \$167430 \$168095 \$167430 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11306 \$167431 \$168096 \$167431 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11342 \$167432 \$168097 \$167432 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11378 \$167433 \$168098 \$167433 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11414 \$167434 \$168099 \$167434 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11450 \$167435 \$168100 \$167435 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11486 \$167436 \$168101 \$167436 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11522 \$167437 \$168102 \$167437 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11558 \$167438 \$168103 \$167438 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11594 \$167439 \$168104 \$167439 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=51.84u AS=22.1616p AD=22.1616p PS=117.72u PD=117.72u
M$11990 \$170779 z$26 \$170779 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11991 \$168095 zn$3 \$170779 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11992 \$168095 z$26 \$168095 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$11995 \$170780 zn$3 \$168095 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$11996 \$170780 z$26 \$170780 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$11999 \$170781 zn$3 \$168095 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12000 \$170781 z$26 \$170781 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12002 \$170782 z$26 \$170782 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12003 \$168096 zn$3 \$170782 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12004 \$168096 z$26 \$168096 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12007 \$170783 zn$3 \$168096 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12008 \$170783 z$26 \$170783 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12011 \$170784 zn$3 \$168096 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12012 \$170784 z$26 \$170784 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12014 \$170785 z$26 \$170785 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12015 \$168097 zn$3 \$170785 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12016 \$168097 z$26 \$168097 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12019 \$170786 zn$3 \$168097 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12020 \$170786 z$26 \$170786 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12023 \$170787 zn$3 \$168097 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12024 \$170787 z$26 \$170787 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12026 \$170788 z$26 \$170788 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12027 \$168098 zn$3 \$170788 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12028 \$168098 z$26 \$168098 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12031 \$170789 zn$3 \$168098 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12032 \$170789 z$26 \$170789 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12035 \$170790 zn$3 \$168098 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12036 \$170790 z$26 \$170790 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12038 \$170791 z$26 \$170791 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12039 \$168099 zn$3 \$170791 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12040 \$168099 z$26 \$168099 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12043 \$170792 zn$3 \$168099 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12044 \$170792 z$26 \$170792 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12047 \$170793 zn$3 \$168099 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12048 \$170793 z$26 \$170793 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12050 \$170794 z$26 \$170794 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12051 \$168100 zn$3 \$170794 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12052 \$168100 z$26 \$168100 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12055 \$170795 zn$3 \$168100 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12056 \$170795 z$26 \$170795 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12059 \$170796 zn$3 \$168100 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12060 \$170796 z$26 \$170796 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12062 \$170797 z$26 \$170797 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12063 \$168101 zn$3 \$170797 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12064 \$168101 z$26 \$168101 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12067 \$170798 zn$3 \$168101 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12068 \$170798 z$26 \$170798 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12071 \$170799 zn$3 \$168101 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12072 \$170799 z$26 \$170799 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12074 \$170800 z$26 \$170800 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12075 \$168102 zn$3 \$170800 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12076 \$168102 z$26 \$168102 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12079 \$170801 zn$3 \$168102 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12080 \$170801 z$26 \$170801 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12083 \$170802 zn$3 \$168102 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12084 \$170802 z$26 \$170802 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12086 \$170803 z$26 \$170803 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12087 \$168103 zn$3 \$170803 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12088 \$168103 z$26 \$168103 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12091 \$170804 zn$3 \$168103 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12092 \$170804 z$26 \$170804 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12095 \$170805 zn$3 \$168103 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12096 \$170805 z$26 \$170805 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12098 \$170806 z$26 \$170806 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12099 \$168104 zn$3 \$170806 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12100 \$168104 z$26 \$168104 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=1.08u AS=0.6102p AD=0.6102p PS=5.55u PD=5.55u
M$12103 \$170807 zn$3 \$168104 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12104 \$170807 z$26 \$170807 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12107 \$170808 zn$3 \$168104 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.72u AS=0.4068p AD=0.4068p PS=3.7u PD=3.7u
M$12108 \$170808 z$26 \$170808 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.36u AS=0.2034p AD=0.2034p PS=1.85u PD=1.85u
M$12110 a1|z$9 a1|i|q$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$12111 a1|z$10 a1|b|i|q$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p PS=2.57u PD=2.57u
M$12112 VSS|anode|cathode|vss a2|a3|z a2|zn$5 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.2988p PS=2.57u PD=1.55u
M$12113 a2|zn$5 RST|a1|b|cdn|core|i|p2c VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.2988p AD=0.4068p
+ PS=1.55u PD=2.57u
M$12114 a1|z$4 RESULT[3]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.72u AS=0.4068p AD=0.4068p
+ PS=2.57u PD=2.57u
M$12115 \$200626 DOUT_DAT|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$12116 \$202259 DOUT_DAT|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$12117 VSS|anode|cathode|vss \$212052 RD[6]|a2|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12118 VSS|anode|cathode|vss i \$211248 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12119 VSS|anode|cathode|vss \$211248 RD[1]|a2|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12120 VSS|anode|cathode|vss \$212053 RD[13]|a4|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12121 VSS|anode|cathode|vss i$1 \$211251 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12122 VSS|anode|cathode|vss \$211251 RD[0]|a2|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12123 \$211252 \$211252 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12124 \$211253 \$211253 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12125 VSS|anode|cathode|vss \$213964 RD[5]|a2|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12126 VSS|anode|cathode|vss \$213965 RD[7]|a2|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12127 VSS|anode|cathode|vss R[13]|i|i0|q \$213461 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12128 VSS|anode|cathode|vss \$213461 RD[45]|a4|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12129 VSS|anode|cathode|vss R[15]|i|i0|q \$213462 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12130 VSS|anode|cathode|vss \$213462 RD[47]|a4|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12131 VSS|anode|cathode|vss i$2 \$213463 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12132 VSS|anode|cathode|vss \$213463 RD[3]|a2|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12133 VSS|anode|cathode|vss R[6]|i|i0|q \$213464 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12134 VSS|anode|cathode|vss \$213464 RD[38]|a2|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12135 VSS|anode|cathode|vss \$213970 RD[31]|a2|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12136 VSS|anode|cathode|vss \$215219 \$215219 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12137 VSS|anode|cathode|vss \$215220 \$215220 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12138 VSS|anode|cathode|vss R[12]|i|i0|q \$213466 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12139 VSS|anode|cathode|vss \$213466 RD[44]|a4|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12140 VSS|anode|cathode|vss \$215221 \$215221 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12141 VSS|anode|cathode|vss \$215222 \$215222 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12142 RD[46]|a4|z \$213468 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12143 VSS|anode|cathode|vss R[14]|i|i0|q \$213468 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12144 VSS|anode|cathode|vss \$213974 RD[14]|a4|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12145 VSS|anode|cathode|vss R[2]|i|i0|q \$213469 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12146 VSS|anode|cathode|vss \$213469 RD[34]|a2|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12147 \$215224 \$215224 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12148 VSS|anode|cathode|vss R[8]|i|i0|q \$213470 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12149 VSS|anode|cathode|vss \$213470 RD[40]|a4|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12150 RD[12]|a4|zn \$213978 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12151 RD[10]|a4|zn \$213979 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12152 RD[42]|a4|z \$213471 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12153 VSS|anode|cathode|vss R[10]|i|i0|q \$213471 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12154 RD[37]|a2|z \$213472 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12155 VSS|anode|cathode|vss R[5]|i|i0|q \$213472 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12156 RD[41]|a4|z \$213473 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12157 VSS|anode|cathode|vss R[9]|i|i0|q \$213473 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12158 RD[35]|a2|z \$213474 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12159 VSS|anode|cathode|vss R[3]|i|i0|q \$213474 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12160 RD[36]|a2|z \$213475 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12161 VSS|anode|cathode|vss R[4]|i|i0|q \$213475 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12162 VSS|anode|cathode|vss R[11]|i|i0|q \$213476 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12163 VSS|anode|cathode|vss \$213476 RD[43]|a4|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12164 RD[18]|a4|zn \$213984 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12165 VSS|anode|cathode|vss \$213985 RD[16]|a4|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12166 RD[33]|a2|z \$213477 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12167 VSS|anode|cathode|vss R[1]|i|i0|q \$213477 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12168 VSS|anode|cathode|vss \$213987 RD[11]|a4|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12169 VSS|anode|cathode|vss \$213988 RD[20]|a4|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12170 RD[25]|a2|zn \$213989 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12171 RD[2]|a2|z \$213478 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12172 VSS|anode|cathode|vss i$3 \$213478 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12173 VSS|anode|cathode|vss R[0]|i|i0|q \$213479 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12174 VSS|anode|cathode|vss \$213479 RD[32]|a2|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12175 \$215232 \$215232 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12176 RD[4]|a2|z \$213480 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12177 VSS|anode|cathode|vss i$4 \$213480 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12178 RD[15]|a4|zn \$213993 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12179 RD[39]|a2|z \$213481 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12180 VSS|anode|cathode|vss R[7]|i|i0|q \$213481 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12181 RD[27]|a2|zn \$213995 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12182 RD[22]|a4|zn \$213996 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12183 RD[29]|a2|zn \$213997 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12184 VSS|anode|cathode|vss cp|z$4 \$230012 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12185 VSS|anode|cathode|vss \$230012 \$229341 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12186 \$230013 \$229341 \$230052 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12187 \$230052 \$230014 \$230053 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12188 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$230053
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12189 \$229342 \$230012 \$230015 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12190 VSS|anode|cathode|vss \$230012 \$230114 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12191 \$230114 d|z$8 \$230013 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12192 VSS|anode|cathode|vss \$230013 \$230014 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12193 \$230014 \$229341 \$229342 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12194 VSS|anode|cathode|vss \$230016 \$230015 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12195 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$230113
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12196 \$230113 \$229342 \$230016 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12197 VSS|anode|cathode|vss \$230016 R[51]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12198 \$230017 s|zn \$230018 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12199 \$230019 \$229344 \$230017 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12200 VSS|anode|cathode|vss i0|i1|q \$230019 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12201 VSS|anode|cathode|vss R[48]|i1|q \$230018 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12202 VSS|anode|cathode|vss s|zn \$229344 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12203 VSS|anode|cathode|vss \$230017 d|z$5 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12204 \$230021 s|zn$1 \$230022 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12205 \$230023 \$229345 \$230021 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12206 VSS|anode|cathode|vss i0|i1|q \$230023 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12207 VSS|anode|cathode|vss R[56]|i1|q \$230022 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12208 VSS|anode|cathode|vss s|zn$1 \$229345 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12209 VSS|anode|cathode|vss \$230021 d|z$6 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12210 \$230026 s|zn \$230027 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12211 \$230028 \$229346 \$230026 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12212 VSS|anode|cathode|vss i0|i1|q$1 \$230028 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12213 VSS|anode|cathode|vss R[51]|i1|q \$230027 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12214 VSS|anode|cathode|vss s|zn \$229346 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12215 VSS|anode|cathode|vss \$230026 d|z$8 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12216 \$229347 a1|a3|i|i1|q \$230111 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12217 \$230111 a2|z$9 \$230112 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12218 \$230112 a1|i|i0|i1|q a4|zn$1 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12219 VSS|anode|cathode|vss RD[45]|a4|z \$229347 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12220 \$229348 RD[38]|a2|z \$230109 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12221 \$230109 a1|a3|i|i1|q a1|zn$1 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12222 VSS|anode|cathode|vss a2|a3|zn$1 \$229348 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12223 \$229349 RD[1]|a2|z \$230110 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12224 \$230110 a1|a3|z a2|zn$7 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12225 VSS|anode|cathode|vss a2|a3|zn$1 \$229349 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12226 \$229350 a3|zn \$230106 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12227 \$230106 a2|zn$13 \$230107 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12228 \$230107 a1|zn$4 a2|zn$12 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12229 VSS|anode|cathode|vss a4|zn$1 \$229350 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12230 VSS|anode|cathode|vss a2|zn$11 \$230108 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12231 \$230108 a1|zn$5 a1|zn$2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12232 VSS|anode|cathode|vss a2|zn$7 \$230103 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12233 \$230103 a1|zn$10 \$230032 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12234 VSS|anode|cathode|vss \$230032 a1|z$14 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12235 \$229351 RD[37]|a2|z \$230104 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12236 \$230104 a1|a3|i|i1|q a3|zn VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12237 VSS|anode|cathode|vss a2|a3|zn$1 \$229351 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12238 \$229353 RD[26]|a2|z \$230105 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12239 \$230105 a1|a3|z a1|zn$3 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12240 VSS|anode|cathode|vss a2|a3|z$1 \$229353 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12241 \$229354 a1|a3|z \$230099 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12242 \$230099 a2|i|i0|i1|q \$230100 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12243 \$230100 a1|z$15 a2|zn$8 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12244 VSS|anode|cathode|vss RD[18]|a4|zn \$229354 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12245 VSS|anode|cathode|vss a2|zn$20 \$230101 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12246 \$230101 a1|zn$6 a1|zn$8 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12247 VSS|anode|cathode|vss a2|zn$9 \$230102 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12248 \$230102 a1|zn$7 \$230037 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12249 VSS|anode|cathode|vss \$230037 a2|z$8 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12250 \$229355 RD[34]|a2|z \$230097 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12251 \$230097 a1|a3|i|i1|q a1|zn$6 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12252 VSS|anode|cathode|vss a2|a3|zn$1 \$229355 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12253 \$229356 a1|a3|i|i1|q \$230098 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12254 \$230098 a2|z$9 \$230095 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12255 \$230095 a1|i|i0|i1|q a4|zn VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12256 VSS|anode|cathode|vss RD[43]|a4|z \$229356 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12257 \$229357 RD[28]|a2|z \$230096 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12258 \$230096 a1|a3|z a2|zn$10 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12259 VSS|anode|cathode|vss a2|a3|z$1 \$229357 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12260 \$229358 a1|a3|z \$230092 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12261 \$230092 a2|z$9 \$230091 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12262 \$230091 a1|i|i0|i1|q a1|zn VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12263 VSS|anode|cathode|vss RD[15]|a4|zn \$229358 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12264 \$229359 a1|a3|z \$230093 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12265 \$230093 a2|z$9 \$230094 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12266 \$230094 a1|i|i0|i1|q a2|zn$9 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12267 VSS|anode|cathode|vss RD[9]|a4|z \$229359 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12268 \$230041 s|zn$1 \$230042 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12269 \$230043 \$229361 \$230041 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12270 VSS|anode|cathode|vss i0|i1|q$1 \$230043 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12271 VSS|anode|cathode|vss R[59]|i1|q \$230042 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12272 VSS|anode|cathode|vss s|zn$1 \$229361 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12273 VSS|anode|cathode|vss \$230041 d|z$7 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12274 VSS|anode|cathode|vss cp|i|z$1 \$230045 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12275 VSS|anode|cathode|vss \$230045 \$229362 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12276 \$230046 \$229362 \$230050 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12277 \$230050 \$230047 \$230051 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12278 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$230051
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12279 \$229363 \$230045 \$230048 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12280 VSS|anode|cathode|vss \$230045 \$230090 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12281 \$230090 d|z$7 \$230046 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12282 VSS|anode|cathode|vss \$230046 \$230047 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12283 \$230047 \$229362 \$229363 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12284 VSS|anode|cathode|vss \$230049 \$230048 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12285 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$230089
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12286 \$230089 \$229363 \$230049 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12287 VSS|anode|cathode|vss \$230049 R[59]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12288 DATA|core|i0|i1|p2c \$231093 VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p
+ PS=6.18u PD=6.18u
M$12289 \$231704 s|zn$2 \$231703 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12290 \$231704 R[35]|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12291 VSS|anode|cathode|vss i0|i1|q$1 \$231705 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12292 \$231705 \$231480 \$231703 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12293 VSS|anode|cathode|vss s|zn$2 \$231480 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12294 VSS|anode|cathode|vss \$231703 d|z$9 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12295 VSS|anode|cathode|vss \$232244 \$233376 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12296 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$233408
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12297 \$233408 \$231711 \$232244 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12298 VSS|anode|cathode|vss \$232244 R[48]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12299 VSS|anode|cathode|vss \$232246 \$233377 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12300 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$233419
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12301 \$233419 \$231716 \$232246 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12302 VSS|anode|cathode|vss \$232246 R[56]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12303 \$233378 a1|a3|i|i1|q \$233415 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12304 \$233415 a2|z$9 \$233426 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12305 \$233426 a1|i|i0|i1|q a4|zn$2 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12306 \$233378 RD[42]|a4|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12307 \$233379 a1|a3|i|i1|q \$233423 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12308 \$233423 a2|z$9 \$233421 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12309 \$233421 a1|i|i0|i1|q a3|zn$2 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12310 \$233379 RD[41]|a4|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12311 \$233380 a3|zn$3 \$233430 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12312 \$233430 a2|z$10 \$233429 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12313 \$233429 a1|zn$9 i1|zn VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12314 \$233380 a4|z VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12315 \$233381 a1|a3|z \$233436 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12316 \$233436 a2|i|i0|i1|q \$233435 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12317 \$233435 a1|z$15 a2|zn$13 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12318 \$233381 RD[21]|a4|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12319 \$233382 a1|a3|z \$233432 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12320 \$233432 a2|i|i0|i1|q \$233431 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12321 \$233431 a1|z$15 a1|zn$10 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12322 \$233382 RD[17]|a4|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12323 \$233383 a1|a3|z \$233433 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12324 \$233433 a2|z$9 \$233434 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12325 \$233434 a1|i|i0|i1|q a1|zn$5 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12326 \$233383 RD[13]|a4|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12327 \$233384 a1|a3|z \$233427 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12328 \$233427 a2|i|i0|i1|q \$233428 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12329 \$233428 a1|z$15 a2|zn$14 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12330 \$233384 RD[19]|a4|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12331 \$233385 a3|zn$5 \$233422 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12332 \$233422 a2|zn$14 \$233420 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12333 \$233420 a1|zn$14 a2|zn$15 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12334 \$233385 a4|zn VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12335 \$233386 a3|zn$7 \$233424 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12336 \$233424 a2|zn$8 \$233425 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12337 \$233425 a1|zn$3 a2|zn$16 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12338 \$233386 a4|zn$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12339 \$233387 a1|a3|i|i1|q \$233417 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12340 \$233417 a2|z$9 \$233418 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12341 \$233418 a1|i|i0|i1|q a4|zn$3 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12342 \$233387 RD[44]|a4|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12343 \$233388 a3|zn$2 \$233411 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12344 \$233411 a2|z$8 \$233412 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12345 \$233412 a1|z$14 i1|zn$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12346 \$233388 a4|zn$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12347 \$233389 RD[25]|a2|zn \$233416 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12348 \$233416 a1|a3|z a4|zn$4 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12349 \$233389 a2|a3|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12350 \$233390 a3|zn$1 \$233407 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12351 \$233407 a2|zn$10 \$233409 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12352 \$233409 a1|zn$13 a2|zn$17 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12353 \$233390 a4|zn$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12354 \$233391 a1|a3|z \$233400 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12355 \$233400 a2|z$9 \$233401 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12356 \$233401 a1|i|i0|i1|q a1|zn$11 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12357 \$233391 RD[11]|a4|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12358 \$233392 a1|a3|z \$233405 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12359 \$233405 a2|z$9 \$233406 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12360 \$233406 a1|i|i0|i1|q a1|zn$12 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12361 \$233392 RD[8]|a4|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12362 \$233393 RD[4]|a2|z \$233399 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12363 \$233399 a1|a3|z a1|zn$13 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12364 \$233393 a2|a3|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12365 \$231733 s|zn$1 \$231732 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12366 \$231733 R[58]|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12367 VSS|anode|cathode|vss i0|i1|q$2 \$231734 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12368 \$231734 \$231484 \$231732 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12369 VSS|anode|cathode|vss s|zn$1 \$231484 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12370 VSS|anode|cathode|vss \$231732 d|z$10 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12371 VSS|anode|cathode|vss \$232250 \$233394 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12372 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$233396
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12373 \$233396 \$231740 \$232250 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12374 VSS|anode|cathode|vss \$232250 R[50]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12375 \$231707 cp|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12376 VSS|anode|cathode|vss \$231707 \$231708 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12377 VSS|anode|cathode|vss \$231707 \$233404 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12378 \$233404 d|z$5 \$231709 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12379 \$231709 \$231708 \$233403 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12380 \$233403 \$232243 \$233402 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12381 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$233402
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12382 \$232243 \$231709 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12383 \$232243 \$231708 \$231711 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12384 \$231711 \$231707 \$233376 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12385 \$231712 cp|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12386 VSS|anode|cathode|vss \$231712 \$231713 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12387 VSS|anode|cathode|vss \$231712 \$233414 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12388 \$233414 d|z$6 \$231714 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12389 \$231714 \$231713 \$233413 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12390 \$233413 \$232245 \$233410 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12391 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$233410
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12392 \$232245 \$231714 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12393 \$232245 \$231713 \$231716 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12394 \$231716 \$231712 \$233377 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12395 \$231736 cp|i|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12396 VSS|anode|cathode|vss \$231736 \$231737 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12397 VSS|anode|cathode|vss \$231736 \$233397 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12398 \$233397 d|z$11 \$231738 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12399 \$231738 \$231737 \$233398 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12400 \$233398 \$232249 \$233395 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12401 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$233395
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12402 \$232249 \$231738 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12403 \$232249 \$231737 \$231740 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12404 \$231740 \$231736 \$233394 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12405 VSS|anode|cathode|vss cp|z$4 \$233645 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12406 VSS|anode|cathode|vss \$233645 \$233646 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12407 \$233647 \$233646 \$234235 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12408 \$234235 \$233648 \$234234 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12409 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$234234
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12410 \$233649 \$233645 \$233650 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12411 VSS|anode|cathode|vss \$233645 \$234237 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12412 \$234237 d|z$16 \$233647 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12413 VSS|anode|cathode|vss \$233647 \$233648 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12414 \$233648 \$233646 \$233649 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12415 VSS|anode|cathode|vss \$233651 \$233650 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12416 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$234240
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12417 \$234240 \$233649 \$233651 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12418 VSS|anode|cathode|vss \$233651 R[53]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12419 \$233652 s|zn$1 \$233653 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12420 \$233654 \$233655 \$233652 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12421 VSS|anode|cathode|vss i0|i1|q$3 \$233654 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12422 VSS|anode|cathode|vss R[60]|i1|q \$233653 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12423 VSS|anode|cathode|vss s|zn$1 \$233655 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12424 VSS|anode|cathode|vss \$233652 d|z$12 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12425 \$233657 s|zn \$233658 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12426 \$233659 \$233660 \$233657 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12427 VSS|anode|cathode|vss i0|i1|q$4 \$233659 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12428 VSS|anode|cathode|vss R[55]|i1|q \$233658 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12429 VSS|anode|cathode|vss s|zn \$233660 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12430 VSS|anode|cathode|vss \$233657 d|z$13 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12431 \$233662 s|z \$233663 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12432 \$233664 \$233665 \$233662 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12433 VSS|anode|cathode|vss R[2]|i|i0|q \$233664 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12434 VSS|anode|cathode|vss i0|i1|q$2 \$233663 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12435 VSS|anode|cathode|vss s|z \$233665 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12436 VSS|anode|cathode|vss \$233662 d|z$14 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12437 \$233667 s|zn \$233668 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12438 \$233669 \$233670 \$233667 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12439 VSS|anode|cathode|vss i0|i1|q$5 \$233669 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12440 VSS|anode|cathode|vss R[53]|i1|q \$233668 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12441 VSS|anode|cathode|vss s|zn \$233670 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12442 VSS|anode|cathode|vss \$233667 d|z$16 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12443 \$233671 a1|a3|i|i1|q \$234254 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12444 \$234254 a2|z$9 \$234253 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12445 \$234253 a1|i|i0|i1|q a2|zn$18 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12446 VSS|anode|cathode|vss RD[47]|a4|z \$233671 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12447 \$233673 RD[30]|a2|z \$234252 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12448 \$234252 a1|a3|z a3|zn$4 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12449 VSS|anode|cathode|vss a2|a3|z$1 \$233673 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12450 \$233675 a1|a3|z \$234250 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12451 \$234250 a2|i|i0|i1|q \$234251 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12452 \$234251 a1|z$15 a1|zn$15 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12453 VSS|anode|cathode|vss RD[23]|a4|z \$233675 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12454 \$233677 RD[6]|a2|zn \$234249 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12455 \$234249 a1|a3|z a1|zn$16 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12456 VSS|anode|cathode|vss a2|a3|zn$1 \$233677 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12457 VSS|anode|cathode|vss a1|zn$2 \$233679 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12458 VSS|anode|cathode|vss a2|zn$12 \$233679 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.374525p AD=0.263525p PS=2.205u PD=1.465u
M$12459 VSS|anode|cathode|vss \$233679 i1|z$1 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.374525p AD=0.358775p PS=2.205u PD=2.4u
M$12460 \$233681 RD[35]|a2|z \$234248 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12461 \$234248 a1|a3|i|i1|q a3|zn$5 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12462 VSS|anode|cathode|vss a2|a3|zn$1 \$233681 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12463 \$233683 RD[0]|a2|z \$234247 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12464 \$234247 a1|a3|z a2|zn$19 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12465 VSS|anode|cathode|vss a2|a3|zn$1 \$233683 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12466 \$233685 a1|a3|z \$234245 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12467 \$234245 a2|z$9 \$234246 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12468 \$234246 a1|i|i0|i1|q a2|zn$20 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12469 VSS|anode|cathode|vss RD[10]|a4|zn \$233685 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12470 \$233687 RD[33]|a2|z \$234244 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12471 \$234244 a1|a3|i|i1|q a1|zn$7 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12472 VSS|anode|cathode|vss a2|a3|zn$1 \$233687 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12473 VSS|anode|cathode|vss a1|zn$8 \$233688 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12474 VSS|anode|cathode|vss a2|zn$16 \$233688 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.374525p AD=0.263525p PS=2.205u PD=1.465u
M$12475 VSS|anode|cathode|vss \$233688 i1|z VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.374525p AD=0.358775p PS=2.205u PD=2.4u
M$12476 \$233689 RD[29]|a2|zn \$234243 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12477 \$234243 a1|a3|z a2|zn$11 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12478 VSS|anode|cathode|vss a2|a3|z$1 \$233689 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12479 \$233690 a1|a3|z \$234241 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12480 \$234241 a2|i|i0|i1|q \$234242 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12481 \$234242 a1|z$15 a3|zn$6 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12482 VSS|anode|cathode|vss RD[16]|a4|zn \$233690 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12483 \$233692 RD[2]|a2|z \$234236 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12484 \$234236 a1|a3|z a3|zn$7 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12485 VSS|anode|cathode|vss a2|a3|zn$1 \$233692 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12486 \$233694 a3|zn$6 \$234238 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12487 \$234238 a2|zn$19 \$234239 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12488 \$234239 a1|zn$12 a1|zn$17 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12489 VSS|anode|cathode|vss a4|zn$5 \$233694 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12490 VSS|anode|cathode|vss a2|zn$24 \$234233 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12491 \$234233 a1|zn$19 a1|zn$18 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12492 \$233695 s|zn \$233696 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12493 \$233697 \$233698 \$233695 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12494 VSS|anode|cathode|vss i0|i1|q$2 \$233697 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12495 VSS|anode|cathode|vss R[50]|i1|q \$233696 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12496 VSS|anode|cathode|vss s|zn \$233698 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12497 VSS|anode|cathode|vss \$233695 d|z$11 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12498 \$233699 s|z \$233700 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12499 \$233701 \$233702 \$233699 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12500 VSS|anode|cathode|vss R[7]|i|i0|q \$233701 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12501 VSS|anode|cathode|vss i0|i1|q$4 \$233700 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12502 VSS|anode|cathode|vss s|z \$233702 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12503 VSS|anode|cathode|vss \$233699 d|z$15 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12504 VSS|anode|cathode|vss cp|i|z$1 \$233704 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12505 VSS|anode|cathode|vss \$233704 \$233705 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12506 \$233706 \$233705 \$234228 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12507 \$234228 \$233707 \$234229 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12508 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$234229
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12509 \$233708 \$233704 \$233709 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12510 VSS|anode|cathode|vss \$233704 \$234227 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12511 \$234227 d|z$10 \$233706 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12512 VSS|anode|cathode|vss \$233706 \$233707 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12513 \$233707 \$233705 \$233708 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12514 VSS|anode|cathode|vss \$233710 \$233709 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12515 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$234226
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12516 \$234226 \$233708 \$233710 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12517 VSS|anode|cathode|vss \$233710 R[58]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12518 \$235865 s|zn$2 \$235807 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12519 \$235865 R[37]|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12520 VSS|anode|cathode|vss i0|i1|q$5 \$235866 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12521 \$235866 \$235806 \$235807 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12522 VSS|anode|cathode|vss s|zn$2 \$235806 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12523 VSS|anode|cathode|vss \$235807 d|z$17 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12524 VSS|anode|cathode|vss \$236644 \$237596 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12525 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$237791
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12526 \$237791 \$235811 \$236644 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12527 VSS|anode|cathode|vss \$236644 R[55]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12528 VSS|anode|cathode|vss \$236645 \$237597 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12529 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$237787
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12530 \$237787 \$235815 \$236645 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12531 VSS|anode|cathode|vss \$236645 R[2]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12532 \$235870 s|z \$235818 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12533 \$235870 i0|i1|q$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12534 VSS|anode|cathode|vss R[6]|i|i0|q \$235871 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12535 \$235871 \$235816 \$235818 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12536 VSS|anode|cathode|vss s|z \$235816 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12537 VSS|anode|cathode|vss \$235818 d|z$18 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12538 \$237598 a1|a3|i|i1|q \$237785 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12539 \$237785 a2|z$9 \$237786 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12540 \$237786 a1|i|i0|i1|q a2|zn$21 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12541 \$237598 RD[46]|a4|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12542 a4|z$1 \$235874 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12543 \$237599 a1|a3|z \$237783 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12544 \$237783 a2|z$9 \$237784 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12545 \$237784 a1|i|i0|i1|q a2|zn$22 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12546 \$237599 RD[14]|a4|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12547 \$237600 a1|a3|z \$237780 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12548 \$237780 a2|i|i0|i1|q \$237781 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12549 \$237781 a1|z$15 a2|zn$23 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12550 \$237600 RD[22]|a4|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12551 VSS|anode|cathode|vss \$236646 \$237601 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12552 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$237775
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12553 \$237775 \$235822 \$236646 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12554 VSS|anode|cathode|vss \$236646 R[5]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12555 \$237602 RD[3]|a2|z \$237776 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12556 \$237776 a1|a3|z a1|zn$14 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12557 \$237602 a2|a3|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12558 \$237603 a1|a3|z \$237773 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12559 \$237773 a2|z$9 \$237774 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12560 \$237774 a1|i|i0|i1|q a1|zn$19 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12561 \$237603 RD[12]|a4|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12562 \$237604 a1|a3|z \$237771 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12563 \$237771 a2|i|i0|i1|q \$237772 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12564 \$237772 a1|z$15 a2|zn$24 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12565 \$237604 RD[20]|a4|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12566 \$237605 RD[39]|a2|z \$237768 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12567 \$237768 a1|a3|i|i1|q a1|zn$9 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12568 \$237605 a2|a3|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12569 \$237606 RD[24]|a2|z \$237769 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12570 \$237769 a1|a3|z a4|zn$5 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12571 \$237606 a2|a3|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12572 \$237607 RD[27]|a2|zn \$237767 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12573 \$237767 a1|a3|z a2|zn$25 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12574 \$237607 a2|a3|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12575 \$235887 s|zn$1 \$235824 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12576 \$235887 R[63]|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12577 VSS|anode|cathode|vss i0|i1|q$4 \$235888 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12578 \$235888 \$235823 \$235824 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12579 VSS|anode|cathode|vss s|zn$1 \$235823 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12580 VSS|anode|cathode|vss \$235824 d|z$19 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12581 VSS|anode|cathode|vss \$236647 \$237608 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12582 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$237761
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12583 \$237761 \$235828 \$236647 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12584 VSS|anode|cathode|vss \$236647 R[7]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12585 \$235808 cp|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12586 VSS|anode|cathode|vss \$235808 \$235809 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12587 VSS|anode|cathode|vss \$235808 \$237796 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12588 \$237796 d|z$13 \$235868 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12589 \$235868 \$235809 \$237797 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12590 \$237797 \$236600 \$237798 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12591 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$237798
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12592 \$236600 \$235868 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12593 \$236600 \$235809 \$235811 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12594 \$235811 \$235808 \$237596 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12595 \$235812 cp|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12596 VSS|anode|cathode|vss \$235812 \$235813 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12597 VSS|anode|cathode|vss \$235812 \$237794 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12598 \$237794 d|z$14 \$235869 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12599 \$235869 \$235813 \$237789 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12600 \$237789 \$236601 \$237790 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12601 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$237790
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12602 \$236601 \$235869 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12603 \$236601 \$235813 \$235815 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12604 \$235815 \$235812 \$237597 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12605 VSS|anode|cathode|vss a2|zn$22 \$237782 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12606 \$237782 a1|zn$1 \$235874 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12607 \$235819 cp|i|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12608 VSS|anode|cathode|vss \$235819 \$235820 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12609 VSS|anode|cathode|vss \$235819 \$237777 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12610 \$237777 d|z$20 \$235878 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12611 \$235878 \$235820 \$237778 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12612 \$237778 \$236603 \$237779 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12613 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$237779
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12614 \$236603 \$235878 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12615 \$236603 \$235820 \$235822 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12616 \$235822 \$235819 \$237601 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12617 VSS|anode|cathode|vss a1|zn$18 \$235879 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12618 \$235879 a2|zn$17 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.263525p AD=0.374525p PS=1.465u PD=2.205u
M$12619 VSS|anode|cathode|vss \$235879 i1|z$2 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.374525p AD=0.358775p PS=2.205u PD=2.4u
M$12620 VSS|anode|cathode|vss a1|zn$20 \$235885 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12621 \$235885 a2|zn$15 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.263525p AD=0.374525p PS=1.465u PD=2.205u
M$12622 VSS|anode|cathode|vss \$235885 i1|z$3 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.374525p AD=0.358775p PS=2.205u PD=2.4u
M$12623 \$235825 cp|i|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12624 VSS|anode|cathode|vss \$235825 \$235826 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12625 VSS|anode|cathode|vss \$235825 \$237763 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12626 \$237763 d|z$15 \$235890 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12627 \$235890 \$235826 \$237764 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12628 \$237764 \$236605 \$237765 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12629 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$237765
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12630 \$236605 \$235890 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12631 \$236605 \$235826 \$235828 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12632 \$235828 \$235825 \$237608 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12633 VSS|anode|cathode|vss cp|z$4 \$237816 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12634 VSS|anode|cathode|vss \$237816 \$237799 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12635 \$237817 \$237799 \$238561 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12636 \$238561 \$237818 \$238560 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12637 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$238560
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12638 \$237800 \$237816 \$237819 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12639 VSS|anode|cathode|vss \$237816 \$238563 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12640 \$238563 d|z$12 \$237817 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12641 VSS|anode|cathode|vss \$237817 \$237818 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12642 \$237818 \$237799 \$237800 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12643 VSS|anode|cathode|vss \$237820 \$237819 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12644 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$238565
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12645 \$238565 \$237800 \$237820 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12646 VSS|anode|cathode|vss \$237820 R[60]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12647 \$237821 s|zn$1 \$237822 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12648 \$237823 \$237801 \$237821 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12649 VSS|anode|cathode|vss i0|i1|q$6 \$237823 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12650 VSS|anode|cathode|vss R[57]|i1|q \$237822 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12651 VSS|anode|cathode|vss s|zn$1 \$237801 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12652 VSS|anode|cathode|vss \$237821 d|z$21 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12653 \$237825 s|zn$1 \$237826 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12654 \$237827 \$237802 \$237825 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12655 VSS|anode|cathode|vss i0|i1|q$7 \$237827 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12656 VSS|anode|cathode|vss R[62]|i1|q \$237826 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12657 VSS|anode|cathode|vss s|zn$1 \$237802 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12658 VSS|anode|cathode|vss \$237825 d|z$22 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12659 VSS|anode|cathode|vss cp|i|z$2 \$237829 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12660 VSS|anode|cathode|vss \$237829 \$237803 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12661 \$237830 \$237803 \$238591 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12662 \$238591 \$237831 \$238592 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12663 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$238592
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12664 \$237804 \$237829 \$237832 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12665 VSS|anode|cathode|vss \$237829 \$238586 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12666 \$238586 d|z$18 \$237830 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12667 VSS|anode|cathode|vss \$237830 \$237831 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12668 \$237831 \$237803 \$237804 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12669 VSS|anode|cathode|vss \$237833 \$237832 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12670 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$238597
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12671 \$238597 \$237804 \$237833 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12672 VSS|anode|cathode|vss \$237833 R[6]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12673 \$237805 a3|zn$4 \$238605 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12674 \$238605 a2|zn$21 \$238604 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12675 \$238604 a1|z$16 i1|zn$2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12676 VSS|anode|cathode|vss a4|z$1 \$237805 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12677 VSS|anode|cathode|vss a2|zn$23 \$238608 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12678 \$238608 a1|zn$16 \$237834 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12679 VSS|anode|cathode|vss \$237834 a1|z$16 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12680 \$237835 s|z \$237836 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12681 \$237837 \$237806 \$237835 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12682 VSS|anode|cathode|vss R[5]|i|i0|q \$237837 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12683 VSS|anode|cathode|vss i0|i1|q$5 \$237836 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12684 VSS|anode|cathode|vss s|z \$237806 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12685 VSS|anode|cathode|vss \$237835 d|z$20 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12686 VSS|anode|cathode|vss cp|i|z$3 \$237838 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12687 VSS|anode|cathode|vss \$237838 \$237807 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12688 \$237839 \$237807 \$238619 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12689 \$238619 \$237840 \$238618 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12690 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$238618
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12691 \$237808 \$237838 \$237841 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12692 VSS|anode|cathode|vss \$237838 \$238613 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12693 \$238613 d|z$25 \$237839 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12694 VSS|anode|cathode|vss \$237839 \$237840 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12695 \$237840 \$237807 \$237808 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12696 VSS|anode|cathode|vss \$237842 \$237841 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12697 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$238616
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12698 \$238616 \$237808 \$237842 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12699 VSS|anode|cathode|vss \$237842 R[0]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12700 \$237843 s|zn$1 \$237844 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12701 \$237845 \$237809 \$237843 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12702 VSS|anode|cathode|vss i0|i1|q$5 \$237845 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12703 VSS|anode|cathode|vss R[61]|i1|q \$237844 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12704 VSS|anode|cathode|vss s|zn$1 \$237809 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12705 VSS|anode|cathode|vss \$237843 d|z$23 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12706 \$237847 s|zn \$237848 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12707 \$237849 \$237810 \$237847 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12708 VSS|anode|cathode|vss i0|i1|q$7 \$237849 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12709 VSS|anode|cathode|vss R[54]|i1|q \$237848 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12710 VSS|anode|cathode|vss s|zn \$237810 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12711 VSS|anode|cathode|vss \$237847 d|z$24 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12712 \$237811 a1|a2|a4|z \$238609 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12713 \$238609 a1|a3|i|i1|q s|zn$1 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12714 VSS|anode|cathode|vss a2|a3|z$1 \$237811 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12715 VSS|anode|cathode|vss cp|i|z$1 \$237851 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12716 VSS|anode|cathode|vss \$237851 \$237812 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12717 \$237852 \$237812 \$238602 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12718 \$238602 \$237853 \$238603 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12719 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$238603
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12720 \$237813 \$237851 \$237854 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12721 VSS|anode|cathode|vss \$237851 \$238598 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12722 \$238598 d|z$26 \$237852 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12723 VSS|anode|cathode|vss \$237852 \$237853 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12724 \$237853 \$237812 \$237813 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12725 VSS|anode|cathode|vss \$237855 \$237854 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12726 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$238596
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12727 \$238596 \$237813 \$237855 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12728 VSS|anode|cathode|vss \$237855 R[4]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12729 VSS|anode|cathode|vss cp|i|z$1 \$237856 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12730 VSS|anode|cathode|vss \$237856 \$237814 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12731 \$237857 \$237814 \$238593 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12732 \$238593 \$237858 \$238585 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12733 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$238585
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12734 \$237815 \$237856 \$237859 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12735 VSS|anode|cathode|vss \$237856 \$238590 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12736 \$238590 d|z$19 \$237857 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12737 VSS|anode|cathode|vss \$237857 \$237858 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12738 \$237858 \$237814 \$237815 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12739 VSS|anode|cathode|vss \$237860 \$237859 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12740 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$238588
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12741 \$238588 \$237815 \$237860 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12742 VSS|anode|cathode|vss \$237860 R[63]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12743 VSS|anode|cathode|vss \$240877 \$241578 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12744 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242118
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12745 \$242118 \$240238 \$240877 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12746 VSS|anode|cathode|vss \$240877 R[57]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12747 VSS|anode|cathode|vss \$240878 \$241579 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12748 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242131
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12749 \$242131 \$240242 \$240878 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12750 VSS|anode|cathode|vss \$240878 R[62]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12751 \$240303 s|zn \$240243 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12752 \$240303 R[52]|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12753 VSS|anode|cathode|vss i0|i1|q$3 \$240304 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12754 \$240304 \$240244 \$240243 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12755 VSS|anode|cathode|vss s|zn \$240244 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12756 VSS|anode|cathode|vss \$240243 d|z$27 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12757 VSS|anode|cathode|vss \$240880 \$241580 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12758 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242140
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12759 \$242140 \$240248 \$240880 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12760 VSS|anode|cathode|vss \$240880 R[52]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12761 a2|a3|z$1 \$240308 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12762 a2|z$10 \$240309 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12763 a4|z \$240310 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12764 \$240311 s|z \$240249 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12765 \$240311 i0|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12766 VSS|anode|cathode|vss R[0]|i|i0|q \$240312 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12767 \$240312 \$240250 \$240249 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12768 VSS|anode|cathode|vss s|z \$240250 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12769 VSS|anode|cathode|vss \$240249 d|z$25 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12770 VSS|anode|cathode|vss \$240881 \$241581 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12771 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242141
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12772 \$242141 \$240254 \$240881 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12773 VSS|anode|cathode|vss \$240881 R[61]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12774 VSS|anode|cathode|vss \$240882 \$241582 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12775 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242134
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12776 \$242134 \$240258 \$240882 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12777 VSS|anode|cathode|vss \$240882 R[54]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12778 VSS|anode|cathode|vss a2|zn$25 \$242132 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12779 \$242132 a1|zn$11 a1|zn$20 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12780 \$240315 s|zn \$240259 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12781 \$240315 R[49]|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12782 VSS|anode|cathode|vss i0|i1|q$6 \$240316 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12783 \$240316 \$240260 \$240259 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12784 VSS|anode|cathode|vss s|zn \$240260 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12785 VSS|anode|cathode|vss \$240259 d|z$28 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12786 VSS|anode|cathode|vss \$240883 \$241583 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12787 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242125
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12788 \$242125 \$240264 \$240883 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12789 VSS|anode|cathode|vss \$240883 R[49]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12790 \$240235 cp|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12791 VSS|anode|cathode|vss \$240235 \$240236 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12792 VSS|anode|cathode|vss \$240235 \$242113 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12793 \$242113 d|z$21 \$240301 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12794 \$240301 \$240236 \$242115 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12795 \$242115 \$240571 \$242114 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12796 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242114
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12797 \$240571 \$240301 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12798 \$240571 \$240236 \$240238 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12799 \$240238 \$240235 \$241578 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12800 \$240239 cp|i|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12801 VSS|anode|cathode|vss \$240239 \$240240 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12802 VSS|anode|cathode|vss \$240239 \$242120 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12803 \$242120 d|z$22 \$240302 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12804 \$240302 \$240240 \$242127 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12805 \$242127 \$240572 \$242126 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12806 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242126
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12807 \$240572 \$240302 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12808 \$240572 \$240240 \$240242 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12809 \$240242 \$240239 \$241579 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12810 \$240245 cp|i|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12811 VSS|anode|cathode|vss \$240245 \$240246 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12812 VSS|anode|cathode|vss \$240245 \$242133 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12813 \$242133 d|z$27 \$240306 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12814 \$240306 \$240246 \$242139 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12815 \$242139 \$240573 \$242138 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12816 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242138
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12817 \$240573 \$240306 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12818 \$240573 \$240246 \$240248 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12819 \$240248 \$240245 \$241580 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12820 VSS|anode|cathode|vss a2|i|i0|i1|q \$242145 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12821 \$242145 a1|i|i0|i1|q \$240308 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12822 VSS|anode|cathode|vss a2|zn$26 \$242142 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12823 \$242142 a1|zn$15 \$240309 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12824 VSS|anode|cathode|vss a2|zn$18 \$242146 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$12825 \$242146 a1|zn \$240310 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$12826 \$240251 cp|i|z$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12827 VSS|anode|cathode|vss \$240251 \$240252 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12828 VSS|anode|cathode|vss \$240251 \$242147 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12829 \$242147 d|z$23 \$240313 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12830 \$240313 \$240252 \$242143 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12831 \$242143 \$240574 \$242144 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12832 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242144
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12833 \$240574 \$240313 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12834 \$240574 \$240252 \$240254 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12835 \$240254 \$240251 \$241581 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12836 \$240255 cp|i|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12837 VSS|anode|cathode|vss \$240255 \$240256 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12838 VSS|anode|cathode|vss \$240255 \$242135 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12839 \$242135 d|z$24 \$240314 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12840 \$240314 \$240256 \$242136 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12841 \$242136 \$240575 \$242137 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12842 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242137
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12843 \$240575 \$240314 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12844 \$240575 \$240256 \$240258 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12845 \$240258 \$240255 \$241582 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12846 \$240261 cp|i|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$12847 VSS|anode|cathode|vss \$240261 \$240262 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12848 VSS|anode|cathode|vss \$240261 \$242128 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12849 \$242128 d|z$28 \$240318 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12850 \$240318 \$240262 \$242129 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12851 \$242129 \$240576 \$242130 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12852 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242130
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12853 \$240576 \$240318 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$12854 \$240576 \$240262 \$240264 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12855 \$240264 \$240261 \$241583 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12856 VSS|anode|cathode|vss cp|z$4 \$242202 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12857 VSS|anode|cathode|vss \$242202 \$242148 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12858 \$242203 \$242148 \$242744 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12859 \$242744 \$242204 \$242743 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12860 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242743
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12861 \$242149 \$242202 \$242205 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12862 VSS|anode|cathode|vss \$242202 \$242746 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12863 \$242746 d|z$9 \$242203 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12864 VSS|anode|cathode|vss \$242203 \$242204 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12865 \$242204 \$242148 \$242149 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12866 VSS|anode|cathode|vss \$242206 \$242205 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12867 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242751
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12868 \$242751 \$242149 \$242206 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12869 VSS|anode|cathode|vss \$242206 R[35]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12870 VSS|anode|cathode|vss cp|i|z$2 \$242207 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12871 VSS|anode|cathode|vss \$242207 \$242150 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12872 \$242209 \$242150 \$242773 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12873 \$242773 \$242210 \$242771 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12874 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242771
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12875 \$242151 \$242207 \$242211 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12876 VSS|anode|cathode|vss \$242207 \$242760 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12877 \$242760 d|z$29 \$242209 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12878 VSS|anode|cathode|vss \$242209 \$242210 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12879 \$242210 \$242150 \$242151 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12880 VSS|anode|cathode|vss \$242212 \$242211 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12881 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242784
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12882 \$242784 \$242151 \$242212 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12883 VSS|anode|cathode|vss \$242212 R[34]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12884 \$242214 s|z$1 \$242215 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12885 \$242216 \$242152 \$242214 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12886 VSS|anode|cathode|vss R[30]|i0|q \$242216 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12887 VSS|anode|cathode|vss i0|i1|q$7 \$242215 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12888 VSS|anode|cathode|vss s|z$1 \$242152 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12889 VSS|anode|cathode|vss \$242214 d|z$30 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12890 \$242218 s|z$1 \$242219 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12891 \$242220 \$243746 \$242218 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12892 VSS|anode|cathode|vss R[27]|i0|q \$242220 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12893 VSS|anode|cathode|vss i0|i1|q$1 \$242219 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12894 VSS|anode|cathode|vss s|z$1 \$243746 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12895 VSS|anode|cathode|vss \$242218 d|z$31 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12896 z$28 cp|i|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$12897 \$242155 RD[36]|a2|z \$242788 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12898 \$242788 a1|a3|i|i1|q a3|zn$1 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12899 VSS|anode|cathode|vss a2|a3|zn$1 \$242155 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12900 \$242223 s|z$1 \$242224 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12901 \$242226 \$242156 \$242223 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12902 VSS|anode|cathode|vss R[28]|i0|q \$242226 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12903 VSS|anode|cathode|vss i0|i1|q$3 \$242224 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12904 VSS|anode|cathode|vss s|z$1 \$242156 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12905 VSS|anode|cathode|vss \$242223 d|z$32 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12906 VSS|anode|cathode|vss i|z$115 \$242228 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12907 VSS|anode|cathode|vss \$242228 cp|i|z$2 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12908 \$242229 s|z$1 \$242230 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12909 \$242232 \$242157 \$242229 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12910 VSS|anode|cathode|vss R[31]|i0|q \$242232 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12911 VSS|anode|cathode|vss i0|i1|q$4 \$242230 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12912 VSS|anode|cathode|vss s|z$1 \$242157 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12913 VSS|anode|cathode|vss \$242229 d|z$33 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12914 VSS|anode|cathode|vss cp|i|z$3 \$242234 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12915 VSS|anode|cathode|vss \$242234 \$242158 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12916 \$242236 \$242158 \$242802 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12917 \$242802 \$242237 \$242800 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12918 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242800
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12919 \$242159 \$242234 \$242238 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12920 VSS|anode|cathode|vss \$242234 \$242803 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12921 \$242803 d|z$34 \$242236 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12922 VSS|anode|cathode|vss \$242236 \$242237 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12923 \$242237 \$242158 \$242159 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12924 VSS|anode|cathode|vss \$242239 \$242238 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12925 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242806
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12926 \$242806 \$242159 \$242239 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12927 VSS|anode|cathode|vss \$242239 R[39]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12928 \$242240 s|z$1 \$242241 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12929 \$242243 \$242160 \$242240 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12930 VSS|anode|cathode|vss R[25]|i0|q \$242243 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12931 VSS|anode|cathode|vss i0|i1|q$6 \$242241 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12932 VSS|anode|cathode|vss s|z$1 \$242160 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12933 VSS|anode|cathode|vss \$242240 d|z$35 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12934 \$242161 a1|a3|i|i1|q \$242810 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12935 \$242810 a2|i|i0|i1|q \$242804 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$12936 \$242804 a1|z$15 s|zn VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u
+ AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12937 VSS|anode|cathode|vss a1|a2|a4|z \$242161 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12938 \$242162 a1|a2|a4|z \$242808 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12939 \$242808 a1|a3|i|i1|q s|zn$2 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12940 VSS|anode|cathode|vss a2|a3|zn$1 \$242162 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12941 \$242245 s|z \$242246 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12942 \$242247 \$242163 \$242245 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12943 VSS|anode|cathode|vss R[4]|i|i0|q \$242247 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12944 VSS|anode|cathode|vss i0|i1|q$3 \$242246 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12945 VSS|anode|cathode|vss s|z \$242163 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12946 VSS|anode|cathode|vss \$242245 d|z$26 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12947 \$242164 RD[32]|a2|z \$242796 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12948 \$242796 a1|a3|i|i1|q a2|zn$27 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12949 VSS|anode|cathode|vss a2|a3|zn$1 \$242164 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12950 \$242249 s|z \$242250 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$12951 \$242251 \$243748 \$242249 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12952 VSS|anode|cathode|vss R[1]|i|i0|q \$242251 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12953 VSS|anode|cathode|vss i0|i1|q$6 \$242250 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$12954 VSS|anode|cathode|vss s|z \$243748 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12955 VSS|anode|cathode|vss \$242249 d|z$36 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12956 VSS|anode|cathode|vss cp|i|z$1 \$242253 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12957 VSS|anode|cathode|vss \$242253 \$242165 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$12958 \$242255 \$242165 \$242792 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$12959 \$242792 \$242256 \$242783 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$12960 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242783
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$12961 \$242166 \$242253 \$242257 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$12962 VSS|anode|cathode|vss \$242253 \$242789 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$12963 \$242789 d|z$37 \$242255 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$12964 VSS|anode|cathode|vss \$242255 \$242256 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$12965 \$242256 \$242165 \$242166 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$12966 VSS|anode|cathode|vss \$242258 \$242257 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12967 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$242770
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12968 \$242770 \$242166 \$242258 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12969 VSS|anode|cathode|vss \$242258 R[3]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12970 \$244563 s|zn$2 \$244529 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12971 \$244563 R[38]|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12972 VSS|anode|cathode|vss i0|i1|q$7 \$244564 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12973 \$244564 \$244530 \$244529 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12974 VSS|anode|cathode|vss s|zn$2 \$244530 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12975 VSS|anode|cathode|vss \$244529 d|z$38 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12976 \$244566 s|zn$3 \$244531 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$12977 \$244566 i0|i1|q$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$12978 VSS|anode|cathode|vss R[45]|i0|q \$244567 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$12979 \$244567 \$244532 \$244531 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$12980 VSS|anode|cathode|vss s|zn$3 \$244532 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12981 VSS|anode|cathode|vss \$244531 d|z$39 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$12982 cp|z$4 \$244534 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$12983 VSS|anode|cathode|vss i|z$115 \$244534 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$12984 VSS|anode|cathode|vss \$245494 \$245926 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12985 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246295
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12986 \$246295 \$244538 \$245494 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12987 VSS|anode|cathode|vss \$245494 R[30]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12988 VSS|anode|cathode|vss \$245495 \$245927 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12989 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246303
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12990 \$246303 \$244542 \$245495 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12991 VSS|anode|cathode|vss \$245495 R[27]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12992 \$245928 RD[31]|a2|zn \$246302 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$12993 \$246302 a1|a3|z a3|zn$3 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12994 \$245928 a2|a3|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$12995 VSS|anode|cathode|vss \$245496 \$245929 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$12996 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246320
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$12997 \$246320 \$244546 \$245496 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$12998 VSS|anode|cathode|vss \$245496 R[31]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$12999 VSS|anode|cathode|vss \$245497 \$245930 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13000 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246329
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13001 \$246329 \$244550 \$245497 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13002 VSS|anode|cathode|vss \$245497 R[32]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13003 VSS|anode|cathode|vss \$245498 \$245931 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13004 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246327
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13005 \$246327 \$244554 \$245498 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13006 VSS|anode|cathode|vss \$245498 R[25]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13007 a2|z$11 \$244575 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13008 VSS|anode|cathode|vss \$245499 \$245932 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13009 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246298
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13010 \$246298 \$244558 \$245499 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13011 VSS|anode|cathode|vss \$245499 R[33]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13012 z$29 cp|i|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$13013 VSS|anode|cathode|vss \$245500 \$245933 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13014 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246274
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13015 \$246274 \$244562 \$245500 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13016 VSS|anode|cathode|vss \$245500 R[1]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13017 \$244535 cp|i|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13018 VSS|anode|cathode|vss \$244535 \$244536 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13019 VSS|anode|cathode|vss \$244535 \$246285 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13020 \$246285 d|z$30 \$244569 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13021 \$244569 \$244536 \$246281 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13022 \$246281 \$244833 \$246279 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13023 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246279
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13024 \$244833 \$244569 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13025 \$244833 \$244536 \$244538 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13026 \$244538 \$244535 \$245926 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13027 \$244539 cp|i|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13028 VSS|anode|cathode|vss \$244539 \$244540 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13029 VSS|anode|cathode|vss \$244539 \$246299 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13030 \$246299 d|z$31 \$244570 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13031 \$244570 \$244540 \$246297 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13032 \$246297 \$244834 \$246296 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13033 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246296
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13034 \$244834 \$244570 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13035 \$244834 \$244540 \$244542 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13036 \$244542 \$244539 \$245927 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13037 \$244543 cp|i|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13038 VSS|anode|cathode|vss \$244543 \$244544 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13039 VSS|anode|cathode|vss \$244543 \$246306 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13040 \$246306 d|z$33 \$244571 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13041 \$244571 \$244544 \$246314 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13042 \$246314 \$244835 \$246313 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13043 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246313
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13044 \$244835 \$244571 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13045 \$244835 \$244544 \$244546 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13046 \$244546 \$244543 \$245929 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13047 \$244547 cp|i|z$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13048 VSS|anode|cathode|vss \$244547 \$244548 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13049 VSS|anode|cathode|vss \$244547 \$246316 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13050 \$246316 d|z$40 \$244572 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13051 \$244572 \$244548 \$246324 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13052 \$246324 \$244836 \$246323 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13053 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246323
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13054 \$244836 \$244572 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13055 \$244836 \$244548 \$244550 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13056 \$244550 \$244547 \$245930 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13057 \$244551 cp|i|z$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13058 VSS|anode|cathode|vss \$244551 \$244552 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13059 VSS|anode|cathode|vss \$244551 \$246332 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13060 \$246332 d|z$35 \$244574 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13061 \$244574 \$244552 \$246333 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13062 \$246333 \$244837 \$246331 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13063 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246331
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13064 \$244837 \$244574 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13065 \$244837 \$244552 \$244554 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13066 \$244554 \$244551 \$245931 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13067 VSS|anode|cathode|vss a2|a3|zn$1 \$246330 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13068 \$246330 a1|a3|z \$244575 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13069 \$244555 cp|i|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13070 VSS|anode|cathode|vss \$244555 \$244556 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13071 VSS|anode|cathode|vss \$244555 \$246325 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13072 \$246325 d|z$41 \$244577 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13073 \$244577 \$244556 \$246309 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13074 \$246309 \$244838 \$246310 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13075 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246310
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13076 \$244838 \$244577 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13077 \$244838 \$244556 \$244558 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13078 \$244558 \$244555 \$245932 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13079 \$244559 cp|i|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13080 VSS|anode|cathode|vss \$244559 \$244560 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13081 VSS|anode|cathode|vss \$244559 \$246289 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13082 \$246289 d|z$36 \$244579 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13083 \$244579 \$244560 \$246292 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13084 \$246292 \$244839 \$246294 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13085 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$246294
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13086 \$244839 \$244579 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13087 \$244839 \$244560 \$244562 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13088 \$244562 \$244559 \$245933 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13089 VSS|anode|cathode|vss cp|z$4 \$246601 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13090 VSS|anode|cathode|vss \$246601 \$246550 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13091 \$246602 \$246550 \$247066 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13092 \$247066 \$246603 \$247065 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13093 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$247065
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13094 \$246551 \$246601 \$246604 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13095 VSS|anode|cathode|vss \$246601 \$247063 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13096 \$247063 d|z$17 \$246602 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13097 VSS|anode|cathode|vss \$246602 \$246603 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13098 \$246603 \$246550 \$246551 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13099 VSS|anode|cathode|vss \$246605 \$246604 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13100 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$247174
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13101 \$247174 \$246551 \$246605 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13102 VSS|anode|cathode|vss \$246605 R[37]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13103 \$246606 s|zn$2 \$246607 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13104 \$246608 \$246552 \$246606 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13105 VSS|anode|cathode|vss i0|i1|q$2 \$246608 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13106 VSS|anode|cathode|vss R[34]|i1|q \$246607 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13107 VSS|anode|cathode|vss s|zn$2 \$246552 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13108 VSS|anode|cathode|vss \$246606 d|z$29 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13109 \$246609 s|zn$4 \$246610 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13110 \$246611 \$246554 \$246609 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13111 VSS|anode|cathode|vss R[12]|i|i0|q \$246611 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13112 VSS|anode|cathode|vss i0|i1|q$3 \$246610 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13113 VSS|anode|cathode|vss s|zn$4 \$246554 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13114 VSS|anode|cathode|vss \$246609 d|z$42 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13115 \$246555 RD[5]|a2|zn \$247170 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13116 \$247170 a1|a3|z a1|zn$4 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13117 VSS|anode|cathode|vss a2|a3|zn$1 \$246555 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13118 \$246613 s|zn$4 \$246614 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13119 \$246615 \$246556 \$246613 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13120 VSS|anode|cathode|vss R[11]|i|i0|q \$246615 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13121 VSS|anode|cathode|vss i0|i1|q$1 \$246614 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13122 VSS|anode|cathode|vss s|zn$4 \$246556 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13123 VSS|anode|cathode|vss \$246613 d|z$43 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13124 VSS|anode|cathode|vss cp|i|z$2 \$246617 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13125 VSS|anode|cathode|vss \$246617 \$246557 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13126 \$246618 \$246557 \$247068 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13127 \$247068 \$246619 \$247067 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13128 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$247067
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13129 \$246558 \$246617 \$246620 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13130 VSS|anode|cathode|vss \$246617 \$247069 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13131 \$247069 d|z$32 \$246618 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13132 VSS|anode|cathode|vss \$246618 \$246619 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13133 \$246619 \$246557 \$246558 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13134 VSS|anode|cathode|vss \$246621 \$246620 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13135 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$247169
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13136 \$247169 \$246558 \$246621 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13137 VSS|anode|cathode|vss \$246621 R[28]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13138 VSS|anode|cathode|vss a1|i|i0|i1|q a2|a3|zn$1 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13139 a2|a3|zn$1 a2|i|i0|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13140 \$246622 s|zn$2 \$246623 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13141 \$246624 \$246559 \$246622 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13142 VSS|anode|cathode|vss i0|i1|q$4 \$246624 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13143 VSS|anode|cathode|vss R[39]|i1|q \$246623 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13144 VSS|anode|cathode|vss s|zn$2 \$246559 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13145 VSS|anode|cathode|vss \$246622 d|z$34 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13146 \$246625 s|zn$2 \$246626 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13147 \$246627 \$246560 \$246625 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13148 VSS|anode|cathode|vss i0|i1|q \$246627 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13149 VSS|anode|cathode|vss R[32]|i1|q \$246626 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13150 VSS|anode|cathode|vss s|zn$2 \$246560 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13151 VSS|anode|cathode|vss \$246625 d|z$40 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13152 z$30 cp|i|z$3 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$13153 VSS|anode|cathode|vss i|z$115 \$246629 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13154 VSS|anode|cathode|vss \$246629 cp|i|z$3 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13155 VSS|anode|cathode|vss a2|a3|z$1 \$247167 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13156 \$247167 a1|a3|z \$246631 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13157 VSS|anode|cathode|vss \$246631 a2|z$12 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13158 VSS|anode|cathode|vss a2|z$12 \$247166 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13159 \$247166 a1|a2|a4|z \$246633 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13160 VSS|anode|cathode|vss \$246633 s|z$1 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13161 \$246634 s|zn$2 \$246635 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13162 \$246636 \$246561 \$246634 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13163 VSS|anode|cathode|vss i0|i1|q$3 \$246636 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13164 VSS|anode|cathode|vss R[36]|i1|q \$246635 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13165 VSS|anode|cathode|vss s|zn$2 \$246561 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13166 VSS|anode|cathode|vss \$246634 d|z$44 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13167 VSS|anode|cathode|vss cp|i|z$3 \$246638 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13168 VSS|anode|cathode|vss \$246638 \$246562 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13169 \$246639 \$246562 \$247073 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13170 \$247073 \$246640 \$247072 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13171 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$247072
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13172 \$246563 \$246638 \$246641 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13173 VSS|anode|cathode|vss \$246638 \$247071 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13174 \$247071 d|z$44 \$246639 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13175 VSS|anode|cathode|vss \$246639 \$246640 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13176 \$246640 \$246562 \$246563 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13177 VSS|anode|cathode|vss \$246642 \$246641 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13178 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$247165
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13179 \$247165 \$246563 \$246642 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13180 VSS|anode|cathode|vss \$246642 R[36]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13181 \$246643 s|z \$246644 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13182 \$246645 \$246564 \$246643 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13183 VSS|anode|cathode|vss R[3]|i|i0|q \$246645 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13184 VSS|anode|cathode|vss i0|i1|q$1 \$246644 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13185 VSS|anode|cathode|vss s|z \$246564 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13186 VSS|anode|cathode|vss \$246643 d|z$37 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13187 VSS|anode|cathode|vss i|z$115 \$246646 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13188 VSS|anode|cathode|vss \$246646 cp|i|z$1 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13189 VSS|anode|cathode|vss \$249190 \$250309 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13190 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$250598
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13191 \$250598 \$249104 \$249190 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13192 VSS|anode|cathode|vss \$249190 R[38]|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13193 \$249106 s|zn$4 \$249105 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13194 \$249106 i0|i1|q$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13195 VSS|anode|cathode|vss R[15]|i|i0|q \$249107 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13196 \$249107 \$249094 \$249105 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13197 VSS|anode|cathode|vss s|zn$4 \$249094 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13198 VSS|anode|cathode|vss \$249105 d|z$45 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13199 VSS|anode|cathode|vss \$249192 \$250310 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13200 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$250602
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13201 \$250602 \$249113 \$249192 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13202 VSS|anode|cathode|vss \$249192 R[15]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13203 VSS|anode|cathode|vss \$249194 \$250311 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13204 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$250609
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13205 \$250609 \$249118 \$249194 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13206 VSS|anode|cathode|vss \$249194 R[11]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13207 a1|z$15 a1|i|i0|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$13208 \$249120 s|z$1 \$249119 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13209 \$249120 i0|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13210 VSS|anode|cathode|vss R[24]|i0|q \$249121 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13211 \$249121 \$249095 \$249119 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13212 VSS|anode|cathode|vss s|z$1 \$249095 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13213 VSS|anode|cathode|vss \$249119 d|z$46 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13214 \$249124 s|zn$4 \$249123 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13215 \$249124 i0|i1|q$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13216 VSS|anode|cathode|vss R[14]|i|i0|q \$249125 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13217 \$249125 \$249096 \$249123 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13218 VSS|anode|cathode|vss s|zn$4 \$249096 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13219 VSS|anode|cathode|vss \$249123 d|z$47 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13220 \$249128 s|z$1 \$249127 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13221 \$249128 i0|i1|q$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13222 VSS|anode|cathode|vss R[29]|i0|q \$249129 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13223 \$249129 \$249097 \$249127 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13224 VSS|anode|cathode|vss s|z$1 \$249097 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13225 VSS|anode|cathode|vss \$249127 d|z$48 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13226 \$250312 a2|i|i0|i1|q \$250608 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13227 \$250608 a1|z$15 a2|zn$28 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13228 \$250312 a1|a3|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13229 \$250313 a2|z$9 \$250611 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13230 \$250611 a1|i|i0|i1|q a2|zn$29 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13231 \$250313 a1|a3|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13232 s|z \$249133 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13233 \$249135 s|zn$2 \$249134 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13234 \$249135 R[33]|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13235 VSS|anode|cathode|vss i0|i1|q$6 \$249136 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13236 \$249136 \$249098 \$249134 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13237 VSS|anode|cathode|vss s|zn$2 \$249098 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13238 VSS|anode|cathode|vss \$249134 d|z$41 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13239 \$249138 s|zn$4 \$249137 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13240 \$249138 i0|i1|q$6 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13241 VSS|anode|cathode|vss R[9]|i|i0|q \$249139 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13242 \$249139 \$249099 \$249137 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13243 VSS|anode|cathode|vss s|zn$4 \$249099 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13244 VSS|anode|cathode|vss \$249137 d|z$49 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13245 VSS|anode|cathode|vss \$249198 \$250314 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13246 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$250578
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13247 \$250578 \$249145 \$249198 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13248 VSS|anode|cathode|vss \$249198 R[9]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13249 \$249100 cp|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13250 VSS|anode|cathode|vss \$249100 \$249101 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13251 VSS|anode|cathode|vss \$249100 \$250579 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13252 \$250579 d|z$38 \$249102 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13253 \$249102 \$249101 \$250599 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13254 \$250599 \$249189 \$250600 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13255 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$250600
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13256 \$249189 \$249102 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13257 \$249189 \$249101 \$249104 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13258 \$249104 \$249100 \$250309 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13259 \$249109 cp|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13260 VSS|anode|cathode|vss \$249109 \$249110 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13261 VSS|anode|cathode|vss \$249109 \$250601 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13262 \$250601 d|z$45 \$249111 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13263 \$249111 \$249110 \$250605 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13264 \$250605 \$249191 \$250604 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13265 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$250604
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13266 \$249191 \$249111 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13267 \$249191 \$249110 \$249113 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13268 \$249113 \$249109 \$250310 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13269 \$249114 cp|i|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13270 VSS|anode|cathode|vss \$249114 \$249115 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13271 VSS|anode|cathode|vss \$249114 \$250607 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13272 \$250607 d|z$43 \$249116 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13273 \$249116 \$249115 \$250606 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13274 \$250606 \$249193 \$250610 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13275 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$250610
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13276 \$249193 \$249116 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13277 \$249193 \$249115 \$249118 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13278 \$249118 \$249114 \$250311 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13279 VSS|anode|cathode|vss a2|z$11 \$250603 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$13280 \$250603 a1|a2|a4|z \$249133 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$13281 \$249141 cp|i|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13282 VSS|anode|cathode|vss \$249141 \$249142 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13283 VSS|anode|cathode|vss \$249141 \$250589 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13284 \$250589 d|z$49 \$249143 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13285 \$249143 \$249142 \$250591 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13286 \$250591 \$249197 \$250594 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13287 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$250594
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13288 \$249197 \$249143 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13289 \$249197 \$249142 \$249145 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13290 \$249145 \$249141 \$250314 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13291 \$251079 s|zn$3 \$251080 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13292 \$251081 \$250812 \$251079 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13293 VSS|anode|cathode|vss R[42]|i0|q \$251081 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13294 VSS|anode|cathode|vss i0|i1|q$2 \$251080 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13295 VSS|anode|cathode|vss s|zn$3 \$250812 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13296 VSS|anode|cathode|vss \$251079 d|z$50 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13297 \$251083 s|zn$4 \$251084 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13298 \$251085 \$250813 \$251083 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13299 VSS|anode|cathode|vss R[13]|i|i0|q \$251085 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13300 VSS|anode|cathode|vss i0|i1|q$5 \$251084 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13301 VSS|anode|cathode|vss s|zn$4 \$250813 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13302 VSS|anode|cathode|vss \$251083 d|z$51 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13303 VSS|anode|cathode|vss cp|z$4 \$251087 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13304 VSS|anode|cathode|vss \$251087 \$250814 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13305 \$251088 \$250814 \$251137 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13306 \$251137 \$251089 \$251138 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13307 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$251138
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13308 \$250815 \$251087 \$251090 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13309 VSS|anode|cathode|vss \$251087 \$251486 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13310 \$251486 d|z$51 \$251088 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13311 VSS|anode|cathode|vss \$251088 \$251089 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13312 \$251089 \$250814 \$250815 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13313 VSS|anode|cathode|vss \$251091 \$251090 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13314 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$251488
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13315 \$251488 \$250815 \$251091 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13316 VSS|anode|cathode|vss \$251091 R[13]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13317 \$251092 s|zn$3 \$251093 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13318 \$251094 \$250816 \$251092 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13319 VSS|anode|cathode|vss R[44]|i0|q \$251094 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13320 VSS|anode|cathode|vss i0|i1|q$3 \$251093 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13321 VSS|anode|cathode|vss s|zn$3 \$250816 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13322 VSS|anode|cathode|vss \$251092 d|z$52 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13323 \$250817 RD[7]|a2|zn \$251489 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13324 \$251489 a1|a3|z a2|zn$26 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13325 VSS|anode|cathode|vss a2|a3|zn$1 \$250817 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13326 \$251096 s|zn$4 \$251097 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13327 \$251098 \$250818 \$251096 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13328 VSS|anode|cathode|vss R[8]|i|i0|q \$251098 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13329 VSS|anode|cathode|vss i0|i1|q \$251097 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13330 VSS|anode|cathode|vss s|zn$4 \$250818 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13331 VSS|anode|cathode|vss \$251096 d|z$53 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13332 a1|a3|z a1|a3|i|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$13333 a2|z$9 a2|i|i0|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$13334 \$251100 s|z$1 \$251101 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13335 \$251102 \$250819 \$251100 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13336 VSS|anode|cathode|vss R[26]|i0|q \$251102 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13337 VSS|anode|cathode|vss i0|i1|q$2 \$251101 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13338 VSS|anode|cathode|vss s|z$1 \$250819 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13339 VSS|anode|cathode|vss \$251100 d|z$54 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13340 VSS|anode|cathode|vss cp|i|z$3 \$251104 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13341 VSS|anode|cathode|vss \$251104 \$250820 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13342 \$251105 \$250820 \$251135 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13343 \$251135 \$251106 \$251136 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13344 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$251136
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13345 \$250821 \$251104 \$251107 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13346 VSS|anode|cathode|vss \$251104 \$251513 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13347 \$251513 d|z$46 \$251105 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13348 VSS|anode|cathode|vss \$251105 \$251106 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13349 \$251106 \$250820 \$250821 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13350 VSS|anode|cathode|vss \$251108 \$251107 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13351 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$251514
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13352 \$251514 \$250821 \$251108 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13353 VSS|anode|cathode|vss \$251108 R[24]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13354 VSS|anode|cathode|vss cp|i|z$3 \$251109 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13355 VSS|anode|cathode|vss \$251109 \$250822 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13356 \$251110 \$250822 \$251133 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13357 \$251133 \$251111 \$251134 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13358 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$251134
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13359 \$250823 \$251109 \$251112 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13360 VSS|anode|cathode|vss \$251109 \$251518 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13361 \$251518 d|z$48 \$251110 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13362 VSS|anode|cathode|vss \$251110 \$251111 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13363 \$251111 \$250822 \$250823 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13364 VSS|anode|cathode|vss \$251113 \$251112 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13365 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$251519
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13366 \$251519 \$250823 \$251113 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13367 VSS|anode|cathode|vss \$251113 R[29]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13368 VSS|anode|cathode|vss cp|i|z$3 \$251114 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13369 VSS|anode|cathode|vss \$251114 \$250824 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13370 \$251115 \$250824 \$251131 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13371 \$251131 \$251116 \$251132 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13372 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$251132
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13373 \$250825 \$251114 \$251117 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13374 VSS|anode|cathode|vss \$251114 \$251521 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13375 \$251521 d|z$56 \$251115 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13376 VSS|anode|cathode|vss \$251115 \$251116 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13377 \$251116 \$250824 \$250825 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13378 VSS|anode|cathode|vss \$251118 \$251117 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13379 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$251520
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13380 \$251520 \$250825 \$251118 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13381 VSS|anode|cathode|vss \$251118 R[41]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13382 \$251119 s|zn$4 \$251120 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13383 \$251121 \$250826 \$251119 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13384 VSS|anode|cathode|vss R[10]|i|i0|q \$251121 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13385 VSS|anode|cathode|vss i0|i1|q$2 \$251120 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13386 VSS|anode|cathode|vss s|zn$4 \$250826 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13387 VSS|anode|cathode|vss \$251119 d|z$55 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13388 VSS|anode|cathode|vss cp|i|z$1 \$251124 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13389 VSS|anode|cathode|vss \$251124 \$250827 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13390 \$251125 \$250827 \$251129 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13391 \$251129 \$251126 \$251130 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13392 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$251130
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13393 \$250828 \$251124 \$251127 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13394 VSS|anode|cathode|vss \$251124 \$251516 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13395 \$251516 d|z$55 \$251125 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13396 VSS|anode|cathode|vss \$251125 \$251126 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13397 \$251126 \$250827 \$250828 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13398 VSS|anode|cathode|vss \$251128 \$251127 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13399 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$251515
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13400 \$251515 \$250828 \$251128 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13401 VSS|anode|cathode|vss \$251128 R[10]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13402 VSS|anode|cathode|vss \$253477 \$254687 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13403 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$254748
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13404 \$254748 \$252804 \$253477 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13405 VSS|anode|cathode|vss \$253477 R[45]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13406 VSS|anode|cathode|vss \$253479 \$254688 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13407 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$254744
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13408 \$254744 \$252808 \$253479 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13409 VSS|anode|cathode|vss \$253479 R[12]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13410 VSS|anode|cathode|vss \$253481 \$254689 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13411 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$254740
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13412 \$254740 \$252812 \$253481 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13413 VSS|anode|cathode|vss \$253481 R[8]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13414 VSS|anode|cathode|vss \$253483 \$254690 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13415 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$254736
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13416 \$254736 \$252816 \$253483 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13417 VSS|anode|cathode|vss \$253483 R[26]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13418 VSS|anode|cathode|vss \$253485 \$254691 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13419 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$254732
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13420 \$254732 \$252820 \$253485 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13421 VSS|anode|cathode|vss \$253485 R[14]|i|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13422 \$254692 a2|z$9 \$254731 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13423 \$254731 a1|i|i0|i1|q a2|zn$30 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13424 \$254692 a1|a3|i|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13425 \$253384 s|zn$3 \$252821 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13426 \$253384 i0|i1|q$6 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13427 VSS|anode|cathode|vss R[41]|i0|q \$253385 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13428 \$253385 \$252822 \$252821 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13429 VSS|anode|cathode|vss s|zn$3 \$252822 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13430 VSS|anode|cathode|vss \$252821 d|z$56 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13431 VSS|anode|cathode|vss a1|zn$21 s|zn$3 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13432 s|zn$3 a2|zn$30 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13433 \$254693 a1|a3|i|i1|q \$254729 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13434 \$254729 a2|z$9 \$254730 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$13435 \$254730 a1|i|i0|i1|q a3|zn$8 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13436 \$254693 RD[40]|a4|z VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13437 \$253388 a1|zn$17 \$254694 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13438 \$254694 b|z VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.4015p PS=1.53u PD=2.27u
M$13439 VSS|anode|cathode|vss \$253388 d|z$57 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.4015p AD=0.3955p PS=2.27u PD=2.53u
M$13440 \$253388 a2|zn$31 \$254694 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$13441 \$253486 a1|i0|q \$254728 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13442 \$254728 a2|i|s|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.4015p PS=1.53u PD=2.27u
M$13443 VSS|anode|cathode|vss a1|a2|b|q|s \$253486 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.4015p AD=0.3955p PS=2.27u PD=2.53u
M$13444 b|z \$253486 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$13445 \$253391 a2|i|s|zn \$252823 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13446 \$253391 i0|i1|q$8 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13447 VSS|anode|cathode|vss a1|i0|q \$253392 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13448 \$253392 \$252824 \$252823 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13449 VSS|anode|cathode|vss a2|i|s|zn \$252824 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13450 VSS|anode|cathode|vss \$252823 i0|z VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13451 \$253394 a1|a2|b|q|s \$252825 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13452 \$253394 i1|zn$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13453 VSS|anode|cathode|vss i0|z \$253395 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13454 \$253395 \$252826 \$252825 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13455 VSS|anode|cathode|vss a1|a2|b|q|s \$252826 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13456 VSS|anode|cathode|vss \$252825 d|z$58 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13457 \$252801 cp|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13458 VSS|anode|cathode|vss \$252801 \$252802 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13459 VSS|anode|cathode|vss \$252801 \$254749 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13460 \$254749 d|z$39 \$253378 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13461 \$253378 \$252802 \$254750 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13462 \$254750 \$253476 \$254751 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13463 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$254751
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13464 \$253476 \$253378 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13465 \$253476 \$252802 \$252804 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13466 \$252804 \$252801 \$254687 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13467 \$252805 cp|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13468 VSS|anode|cathode|vss \$252805 \$252806 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13469 VSS|anode|cathode|vss \$252805 \$254745 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13470 \$254745 d|z$42 \$253379 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13471 \$253379 \$252806 \$254746 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13472 \$254746 \$253478 \$254747 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13473 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$254747
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13474 \$253478 \$253379 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13475 \$253478 \$252806 \$252808 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13476 \$252808 \$252805 \$254688 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13477 \$252809 cp|i|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13478 VSS|anode|cathode|vss \$252809 \$252810 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13479 VSS|anode|cathode|vss \$252809 \$254741 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13480 \$254741 d|z$53 \$253380 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13481 \$253380 \$252810 \$254742 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13482 \$254742 \$253480 \$254743 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13483 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$254743
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13484 \$253480 \$253380 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13485 \$253480 \$252810 \$252812 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13486 \$252812 \$252809 \$254689 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13487 \$252813 cp|i|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13488 VSS|anode|cathode|vss \$252813 \$252814 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13489 VSS|anode|cathode|vss \$252813 \$254737 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13490 \$254737 d|z$54 \$253381 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13491 \$253381 \$252814 \$254738 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13492 \$254738 \$253482 \$254739 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13493 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$254739
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13494 \$253482 \$253381 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13495 \$253482 \$252814 \$252816 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13496 \$252816 \$252813 \$254690 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13497 \$252817 cp|i|z$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13498 VSS|anode|cathode|vss \$252817 \$252818 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13499 VSS|anode|cathode|vss \$252817 \$254733 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13500 \$254733 d|z$47 \$253382 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13501 \$253382 \$252818 \$254734 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13502 \$254734 \$253484 \$254735 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13503 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$254735
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13504 \$253484 \$253382 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13505 \$253484 \$252818 \$252820 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13506 \$252820 \$252817 \$254691 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13507 VSS|anode|cathode|vss cp|z$4 \$255075 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13508 VSS|anode|cathode|vss \$255075 \$254828 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13509 \$255076 \$254828 \$255440 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13510 \$255440 \$255077 \$255435 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13511 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$255435
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13512 \$254829 \$255075 \$255078 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13513 VSS|anode|cathode|vss \$255075 \$255448 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13514 \$255448 d|z$50 \$255076 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13515 VSS|anode|cathode|vss \$255076 \$255077 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13516 \$255077 \$254828 \$254829 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13517 VSS|anode|cathode|vss \$255079 \$255078 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13518 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$255425
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13519 \$255425 \$254829 \$255079 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13520 VSS|anode|cathode|vss \$255079 R[42]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13521 VSS|anode|cathode|vss cp|z$4 \$255080 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13522 VSS|anode|cathode|vss \$255080 \$254830 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13523 \$255082 \$254830 \$255418 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13524 \$255418 \$255083 \$255422 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13525 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$255422
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13526 \$254831 \$255080 \$255084 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13527 VSS|anode|cathode|vss \$255080 \$255415 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13528 \$255415 d|z$59 \$255082 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13529 VSS|anode|cathode|vss \$255082 \$255083 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13530 \$255083 \$254830 \$254831 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13531 VSS|anode|cathode|vss \$255085 \$255084 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13532 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$255408
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13533 \$255408 \$254831 \$255085 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13534 VSS|anode|cathode|vss \$255085 R[40]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13535 \$255087 s|zn$3 \$255088 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13536 \$255090 \$254832 \$255087 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13537 VSS|anode|cathode|vss R[46]|i0|q \$255090 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13538 VSS|anode|cathode|vss i0|i1|q$7 \$255088 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13539 VSS|anode|cathode|vss s|zn$3 \$254832 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13540 VSS|anode|cathode|vss \$255087 d|z$60 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13541 VSS|anode|cathode|vss cp|i|z$4 \$255092 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13542 VSS|anode|cathode|vss \$255092 \$254833 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13543 \$255093 \$254833 \$255399 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13544 \$255399 \$255094 \$255386 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13545 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$255386
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13546 \$254834 \$255092 \$255095 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13547 VSS|anode|cathode|vss \$255092 \$255398 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13548 \$255398 d|z$60 \$255093 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13549 VSS|anode|cathode|vss \$255093 \$255094 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13550 \$255094 \$254833 \$254834 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13551 VSS|anode|cathode|vss \$255096 \$255095 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13552 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$255395
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13553 \$255395 \$254834 \$255096 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13554 VSS|anode|cathode|vss \$255096 R[46]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13555 VSS|anode|cathode|vss CLK|core|i|p2c$1 \$255097 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13556 VSS|anode|cathode|vss \$255097 i|z$115 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13557 \$255098 s|zn$6 \$255099 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13558 \$255100 \$254835 \$255098 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13559 VSS|anode|cathode|vss R[18]|i0|q \$255100 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13560 VSS|anode|cathode|vss i0|i1|q$2 \$255099 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13561 VSS|anode|cathode|vss s|zn$6 \$254835 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13562 VSS|anode|cathode|vss \$255098 d|z$61 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13563 \$255102 s|zn$3 \$255103 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13564 \$255104 \$254836 \$255102 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13565 VSS|anode|cathode|vss R[43]|i0|q \$255104 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13566 VSS|anode|cathode|vss i0|i1|q$1 \$255103 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13567 VSS|anode|cathode|vss s|zn$3 \$254836 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13568 VSS|anode|cathode|vss \$255102 d|z$62 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13569 \$255106 s|zn$3 \$255107 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13570 \$255108 \$254837 \$255106 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13571 VSS|anode|cathode|vss R[47]|i0|q \$255108 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13572 VSS|anode|cathode|vss i0|i1|q$4 \$255107 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13573 VSS|anode|cathode|vss s|zn$3 \$254837 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13574 VSS|anode|cathode|vss \$255106 d|z$63 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13575 VSS|anode|cathode|vss a1|zn$21 s|zn$4 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13576 s|zn$4 a2|zn$29 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13577 \$254838 a2|zn$27 \$255346 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13578 \$255346 a1|a2|b|q|s a2|zn$31 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13579 VSS|anode|cathode|vss a3|zn$8 \$254838 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13580 VSS|anode|cathode|vss cp|i|z$3 \$255110 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13581 VSS|anode|cathode|vss \$255110 \$254839 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13582 \$255111 \$254839 \$255339 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13583 \$255339 \$255112 \$255324 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13584 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$255324
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13585 \$254840 \$255110 \$255113 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13586 VSS|anode|cathode|vss \$255110 \$255336 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13587 \$255336 d|z$57 \$255111 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13588 VSS|anode|cathode|vss \$255111 \$255112 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13589 \$255112 \$254839 \$254840 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13590 VSS|anode|cathode|vss \$255114 \$255113 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13591 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$255329
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13592 \$255329 \$254840 \$255114 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13593 VSS|anode|cathode|vss \$255114 a1|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13594 VSS|anode|cathode|vss cp|i|z$1 \$255115 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13595 VSS|anode|cathode|vss \$255115 \$254841 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13596 \$255116 \$254841 \$255306 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13597 \$255306 \$255117 \$255307 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13598 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$255307
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13599 \$254842 \$255115 \$255118 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13600 VSS|anode|cathode|vss \$255115 \$255323 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13601 \$255323 d|z$58 \$255116 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13602 VSS|anode|cathode|vss \$255116 \$255117 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13603 \$255117 \$254841 \$254842 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13604 VSS|anode|cathode|vss \$255119 \$255118 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13605 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$255296
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13606 \$255296 \$254842 \$255119 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13607 VSS|anode|cathode|vss \$255119 i0|i1|q$8 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13608 VSS|anode|cathode|vss \$258009 \$258888 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13609 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258918
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13610 \$258918 \$257001 \$258009 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13611 VSS|anode|cathode|vss \$258009 i0|i1|q$7 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13612 \$257749 s|zn$3 \$257002 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13613 \$257749 i0|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13614 VSS|anode|cathode|vss R[40]|i0|q \$257750 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13615 \$257750 \$257003 \$257002 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13616 VSS|anode|cathode|vss s|zn$3 \$257003 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13617 VSS|anode|cathode|vss \$257002 d|z$59 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13618 VSS|anode|cathode|vss \$258011 \$258889 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13619 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258912
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13620 \$258912 \$257007 \$258011 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13621 VSS|anode|cathode|vss \$258011 R[44]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13622 \$257753 s|zn$5 \$257008 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13623 \$257753 a1|a3|i|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13624 VSS|anode|cathode|vss a2|i|i0|i1|q \$257754 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13625 \$257754 \$257009 \$257008 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13626 VSS|anode|cathode|vss s|zn$5 \$257009 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13627 VSS|anode|cathode|vss \$257008 d|z$64 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13628 VSS|anode|cathode|vss \$258012 \$258890 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13629 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258907
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13630 \$258907 \$257013 \$258012 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13631 VSS|anode|cathode|vss \$258012 a1|a3|i|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13632 VSS|anode|cathode|vss \$258014 \$258891 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13633 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258906
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13634 \$258906 \$257017 \$258014 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13635 VSS|anode|cathode|vss \$258014 R[18]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13636 VSS|anode|cathode|vss \$258015 \$258892 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13637 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258900
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13638 \$258900 \$257021 \$258015 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13639 VSS|anode|cathode|vss \$258015 R[43]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13640 VSS|anode|cathode|vss \$258016 \$258893 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13641 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258895
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13642 \$258895 \$257025 \$258016 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13643 VSS|anode|cathode|vss \$258016 R[47]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13644 \$257764 a2|i|s|zn \$257026 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13645 \$257764 i0|i1|q$9 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13646 VSS|anode|cathode|vss i0|i1|q$8 \$257765 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13647 \$257765 \$257027 \$257026 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13648 VSS|anode|cathode|vss a2|i|s|zn \$257027 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13649 VSS|anode|cathode|vss \$257026 i0|z$1 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13650 \$257767 a1|a2|b|q|s \$257028 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13651 \$257767 i1|z VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13652 VSS|anode|cathode|vss i0|z$1 \$257768 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13653 \$257768 \$257029 \$257028 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13654 VSS|anode|cathode|vss a1|a2|b|q|s \$257029 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13655 VSS|anode|cathode|vss \$257028 d|z$65 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13656 CLK|core|i|p2c$1 \$258894 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$13657 \$256998 cp|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13658 VSS|anode|cathode|vss \$256998 \$256999 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13659 VSS|anode|cathode|vss \$256998 \$258915 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13660 \$258915 d|z$66 \$257747 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13661 \$257747 \$256999 \$258916 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13662 \$258916 \$257748 \$258917 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13663 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258917
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13664 \$257748 \$257747 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13665 \$257748 \$256999 \$257001 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13666 \$257001 \$256998 \$258888 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13667 \$257004 cp|i|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13668 VSS|anode|cathode|vss \$257004 \$257005 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13669 VSS|anode|cathode|vss \$257004 \$258913 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13670 \$258913 d|z$52 \$257751 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13671 \$257751 \$257005 \$258914 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13672 \$258914 \$257752 \$258911 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13673 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258911
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13674 \$257752 \$257751 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13675 \$257752 \$257005 \$257007 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13676 \$257007 \$257004 \$258889 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13677 \$257010 cp|i|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13678 VSS|anode|cathode|vss \$257010 \$257011 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13679 VSS|anode|cathode|vss \$257010 \$258908 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13680 \$258908 d|z$64 \$257756 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13681 \$257756 \$257011 \$258909 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13682 \$258909 \$257757 \$258910 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13683 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258910
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13684 \$257757 \$257756 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13685 \$257757 \$257011 \$257013 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13686 \$257013 \$257010 \$258890 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13687 \$257014 cp|i|z$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13688 VSS|anode|cathode|vss \$257014 \$257015 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13689 VSS|anode|cathode|vss \$257014 \$258903 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13690 \$258903 d|z$61 \$257758 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13691 \$257758 \$257015 \$258904 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13692 \$258904 \$257759 \$258905 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13693 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258905
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13694 \$257759 \$257758 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13695 \$257759 \$257015 \$257017 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13696 \$257017 \$257014 \$258891 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13697 \$257018 cp|i|z$6 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13698 VSS|anode|cathode|vss \$257018 \$257019 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13699 VSS|anode|cathode|vss \$257018 \$258901 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13700 \$258901 d|z$62 \$257760 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13701 \$257760 \$257019 \$258902 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13702 \$258902 \$257761 \$258899 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13703 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258899
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13704 \$257761 \$257760 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13705 \$257761 \$257019 \$257021 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13706 \$257021 \$257018 \$258892 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13707 \$257022 cp|i|z$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13708 VSS|anode|cathode|vss \$257022 \$257023 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13709 VSS|anode|cathode|vss \$257022 \$258896 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13710 \$258896 d|z$63 \$257762 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13711 \$257762 \$257023 \$258897 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13712 \$258897 \$257763 \$258898 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13713 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$258898
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13714 \$257763 \$257762 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13715 \$257763 \$257023 \$257025 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13716 \$257025 \$257022 \$258893 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13717 VSS|anode|cathode|vss cp|i|z$7 \$259368 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13718 VSS|anode|cathode|vss \$259368 \$259348 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13719 \$259369 \$259348 \$259707 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13720 \$259707 \$259370 \$259708 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13721 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259708
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13722 \$259349 \$259368 \$259371 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13723 VSS|anode|cathode|vss \$259368 \$259952 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13724 \$259952 d|z$70 \$259369 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13725 VSS|anode|cathode|vss \$259369 \$259370 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13726 \$259370 \$259348 \$259349 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13727 VSS|anode|cathode|vss \$259372 \$259371 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13728 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259955
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13729 \$259955 \$259349 \$259372 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13730 VSS|anode|cathode|vss \$259372 i0|i1|q$5 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13731 \$259373 s|zn$5 \$259374 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13732 \$259375 \$259351 \$259373 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13733 VSS|anode|cathode|vss i0|i1|q$5 \$259375 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13734 VSS|anode|cathode|vss i0|i1|q$7 \$259374 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13735 VSS|anode|cathode|vss s|zn$5 \$259351 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13736 VSS|anode|cathode|vss \$259373 d|z$66 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13737 \$259376 s|zn$6 \$259377 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13738 \$259378 \$259353 \$259376 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13739 VSS|anode|cathode|vss R[16]|i0|q \$259378 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13740 VSS|anode|cathode|vss i0|i1|q \$259377 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13741 VSS|anode|cathode|vss s|zn$6 \$259353 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13742 VSS|anode|cathode|vss \$259376 d|z$67 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13743 \$259380 s|zn$6 \$259381 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13744 \$259382 \$259354 \$259380 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13745 VSS|anode|cathode|vss R[23]|i0|q \$259382 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13746 VSS|anode|cathode|vss i0|i1|q$4 \$259381 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13747 VSS|anode|cathode|vss s|zn$6 \$259354 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13748 VSS|anode|cathode|vss \$259380 d|z$68 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13749 VSS|anode|cathode|vss cp|i|z$4 \$259384 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13750 VSS|anode|cathode|vss \$259384 \$259355 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13751 \$259385 \$259355 \$259692 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13752 \$259692 \$259386 \$259693 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13753 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259693
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13754 \$259356 \$259384 \$259387 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13755 VSS|anode|cathode|vss \$259384 \$259958 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13756 \$259958 d|z$68 \$259385 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13757 VSS|anode|cathode|vss \$259385 \$259386 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13758 \$259386 \$259355 \$259356 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13759 VSS|anode|cathode|vss \$259388 \$259387 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13760 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259954
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13761 \$259954 \$259356 \$259388 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13762 VSS|anode|cathode|vss \$259388 R[23]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13763 VSS|anode|cathode|vss cp|i|z$4 \$259389 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13764 VSS|anode|cathode|vss \$259389 \$259357 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13765 \$259390 \$259357 \$259676 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13766 \$259676 \$259391 \$259677 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13767 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259677
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13768 \$259358 \$259389 \$259392 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13769 VSS|anode|cathode|vss \$259389 \$259949 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13770 \$259949 d|z$71 \$259390 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13771 VSS|anode|cathode|vss \$259390 \$259391 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13772 \$259391 \$259357 \$259358 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13773 VSS|anode|cathode|vss \$259393 \$259392 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13774 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259919
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13775 \$259919 \$259358 \$259393 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13776 VSS|anode|cathode|vss \$259393 a2|i|i0|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13777 VSS|anode|cathode|vss cp|i|z$5 \$259394 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13778 VSS|anode|cathode|vss \$259394 \$259359 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13779 \$259395 \$259359 \$259660 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13780 \$259660 \$259396 \$259661 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13781 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259661
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13782 \$259360 \$259394 \$259397 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13783 VSS|anode|cathode|vss \$259394 \$259914 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13784 \$259914 d|z$72 \$259395 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13785 VSS|anode|cathode|vss \$259395 \$259396 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13786 \$259396 \$259359 \$259360 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13787 VSS|anode|cathode|vss \$259398 \$259397 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13788 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259910
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13789 \$259910 \$259360 \$259398 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13790 VSS|anode|cathode|vss \$259398 R[21]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13791 VSS|anode|cathode|vss a1|zn$21 s|zn$6 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$13792 s|zn$6 a2|zn$28 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13793 VSS|anode|cathode|vss cp|i|z$6 \$259399 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13794 VSS|anode|cathode|vss \$259399 \$259361 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13795 \$259400 \$259361 \$259647 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13796 \$259647 \$259401 \$259649 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13797 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259649
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13798 \$259362 \$259399 \$259402 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13799 VSS|anode|cathode|vss \$259399 \$259907 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13800 \$259907 d|z$73 \$259400 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13801 VSS|anode|cathode|vss \$259400 \$259401 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13802 \$259401 \$259361 \$259362 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13803 VSS|anode|cathode|vss \$259403 \$259402 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13804 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259902
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13805 \$259902 \$259362 \$259403 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13806 VSS|anode|cathode|vss \$259403 R[22]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13807 \$259404 a1|a2|b|q|s \$259405 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13808 \$259406 \$259363 \$259404 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13809 VSS|anode|cathode|vss i0|z$2 \$259406 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13810 VSS|anode|cathode|vss i1|z$3 \$259405 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13811 VSS|anode|cathode|vss a1|a2|b|q|s \$259363 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13812 VSS|anode|cathode|vss \$259404 d|z$69 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13813 VSS|anode|cathode|vss cp|i|z$6 \$259408 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13814 VSS|anode|cathode|vss \$259408 \$259364 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13815 \$259409 \$259364 \$259625 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13816 \$259625 \$259410 \$259626 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13817 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259626
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13818 \$259365 \$259408 \$259411 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13819 VSS|anode|cathode|vss \$259408 \$259882 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13820 \$259882 d|z$65 \$259409 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13821 VSS|anode|cathode|vss \$259409 \$259410 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13822 \$259410 \$259364 \$259365 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13823 VSS|anode|cathode|vss \$259412 \$259411 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13824 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$259870
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13825 \$259870 \$259365 \$259412 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13826 VSS|anode|cathode|vss \$259412 i0|i1|q$9 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13827 \$261263 s|zn$5 \$261262 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13828 \$261263 i0|i1|q$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13829 VSS|anode|cathode|vss i0|i1|q$3 \$261264 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13830 \$261264 \$261217 \$261262 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13831 VSS|anode|cathode|vss s|zn$5 \$261217 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13832 VSS|anode|cathode|vss \$261262 d|z$70 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13833 \$261266 s|zn$5 \$261265 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13834 \$261266 i0|i1|q$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13835 VSS|anode|cathode|vss i0|i1|q$7 \$261267 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13836 \$261267 \$261218 \$261265 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13837 VSS|anode|cathode|vss s|zn$5 \$261218 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13838 VSS|anode|cathode|vss \$261265 d|z$74 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13839 VSS|anode|cathode|vss \$262081 \$263108 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13840 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263126
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13841 \$263126 \$261273 \$262081 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13842 VSS|anode|cathode|vss \$262081 i0|i1|q$4 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13843 VSS|anode|cathode|vss \$262082 \$263109 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13844 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263124
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13845 \$263124 \$261278 \$262082 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13846 VSS|anode|cathode|vss \$262082 a1|i|i0|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13847 \$261280 s|zn$5 \$261279 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13848 \$261280 a2|i|i0|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13849 VSS|anode|cathode|vss a1|i|i0|i1|q \$261281 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13850 \$261281 \$261219 \$261279 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13851 VSS|anode|cathode|vss s|zn$5 \$261219 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13852 VSS|anode|cathode|vss \$261279 d|z$71 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13853 \$261283 s|zn$6 \$261282 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13854 \$261283 i0|i1|q$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13855 VSS|anode|cathode|vss R[21]|i0|q \$261284 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13856 \$261284 \$261220 \$261282 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13857 VSS|anode|cathode|vss s|zn$6 \$261220 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13858 VSS|anode|cathode|vss \$261282 d|z$72 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13859 \$261286 s|zn$6 \$261285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13860 \$261286 i0|i1|q$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13861 VSS|anode|cathode|vss R[20]|i0|q \$261287 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13862 \$261287 \$261221 \$261285 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13863 VSS|anode|cathode|vss s|zn$6 \$261221 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13864 VSS|anode|cathode|vss \$261285 d|z$75 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13865 \$261290 s|zn$6 \$261289 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13866 \$261290 i0|i1|q$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13867 VSS|anode|cathode|vss R[19]|i0|q \$261291 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13868 \$261291 \$261222 \$261289 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13869 VSS|anode|cathode|vss s|zn$6 \$261222 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13870 VSS|anode|cathode|vss \$261289 d|z$76 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13871 \$261294 s|zn$6 \$261293 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13872 \$261294 i0|i1|q$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13873 VSS|anode|cathode|vss R[22]|i0|q \$261295 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13874 \$261295 \$261223 \$261293 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13875 VSS|anode|cathode|vss s|zn$6 \$261223 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13876 VSS|anode|cathode|vss \$261293 d|z$73 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13877 \$261297 a1|a2|b|q|s \$261296 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$13878 \$261297 i1|z$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$13879 VSS|anode|cathode|vss i0|z$3 \$261298 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13880 \$261298 \$261224 \$261296 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13881 VSS|anode|cathode|vss a1|a2|b|q|s \$261224 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13882 VSS|anode|cathode|vss \$261296 d|z$77 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13883 VSS|anode|cathode|vss \$262083 \$263110 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13884 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263113
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13885 \$263113 \$261304 \$262083 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13886 VSS|anode|cathode|vss \$262083 i0|i1|q$10 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13887 VSS|anode|cathode|vss cp|i|z$7 \$263506 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13888 VSS|anode|cathode|vss \$263506 \$263439 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13889 \$263507 \$263439 \$263779 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13890 \$263779 \$263508 \$263778 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13891 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263778
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13892 \$263440 \$263506 \$263509 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13893 VSS|anode|cathode|vss \$263506 \$263781 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13894 \$263781 d|z$81 \$263507 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13895 VSS|anode|cathode|vss \$263507 \$263508 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13896 \$263508 \$263439 \$263440 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13897 VSS|anode|cathode|vss \$263510 \$263509 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13898 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$264062
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13899 \$264062 \$263440 \$263510 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13900 VSS|anode|cathode|vss \$263510 i0|i1|q$1 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13901 VSS|anode|cathode|vss cp|i|z$7 \$263511 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13902 VSS|anode|cathode|vss \$263511 \$263441 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13903 \$261269 cp|i|z$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13904 VSS|anode|cathode|vss \$261269 \$261270 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13905 \$263512 \$263441 \$263793 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13906 \$263793 \$263513 \$263791 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13907 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263791
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13908 \$263442 \$263511 \$263514 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13909 VSS|anode|cathode|vss \$263511 \$263794 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13910 \$263794 d|z$67 \$263512 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13911 VSS|anode|cathode|vss \$263512 \$263513 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13912 \$263513 \$263441 \$263442 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13913 VSS|anode|cathode|vss \$261269 \$263125 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13914 \$263125 d|z$74 \$261271 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13915 \$261271 \$261270 \$263129 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13916 \$263129 \$261847 \$263127 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13917 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263127
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13918 \$261847 \$261271 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13919 \$261847 \$261270 \$261273 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13920 \$261273 \$261269 \$263108 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13921 VSS|anode|cathode|vss \$263515 \$263514 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13922 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$264066
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13923 \$264066 \$263442 \$263515 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13924 VSS|anode|cathode|vss \$263515 R[16]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13925 \$263516 s|zn$5 \$263517 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13926 \$263518 \$263443 \$263516 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13927 VSS|anode|cathode|vss i0|i1|q$4 \$263518 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13928 VSS|anode|cathode|vss a1|i|i0|i1|q \$263517 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13929 \$261274 cp|i|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13930 VSS|anode|cathode|vss \$261274 \$261275 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13931 VSS|anode|cathode|vss \$261274 \$263128 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13932 \$263128 d|z$78 \$261276 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13933 \$261276 \$261275 \$263131 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13934 \$263131 \$261848 \$263130 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13935 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263130
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13936 \$261848 \$261276 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$13937 \$261848 \$261275 \$261278 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13938 \$261278 \$261274 \$263109 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13939 VSS|anode|cathode|vss s|zn$5 \$263443 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13940 VSS|anode|cathode|vss \$263516 d|z$78 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13941 \$263519 a1|a2|b|q|s \$263520 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13942 \$263521 \$263444 \$263519 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13943 VSS|anode|cathode|vss i0|z$4 \$263521 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13944 VSS|anode|cathode|vss i1|zn$2 \$263520 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13945 VSS|anode|cathode|vss a1|a2|b|q|s \$263444 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13946 VSS|anode|cathode|vss \$263519 d|z$79 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13947 \$263523 a1|a2|b|q|s \$263524 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13948 \$263525 \$263445 \$263523 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13949 VSS|anode|cathode|vss i0|z$5 \$263525 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13950 VSS|anode|cathode|vss i1|z$1 \$263524 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13951 VSS|anode|cathode|vss a1|a2|b|q|s \$263445 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13952 VSS|anode|cathode|vss \$263523 d|z$80 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13953 \$263527 a2|i|s|zn \$263528 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$13954 \$263529 \$263446 \$263527 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$13955 VSS|anode|cathode|vss i0|i1|q$12 \$263529 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$13956 VSS|anode|cathode|vss i0|i1|q$11 \$263528 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$13957 VSS|anode|cathode|vss a2|i|s|zn \$263446 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$13958 VSS|anode|cathode|vss \$263527 i0|z$5 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$13959 VSS|anode|cathode|vss cp|i|z$5 \$263530 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13960 VSS|anode|cathode|vss \$263530 \$263447 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13961 \$263531 \$263447 \$263787 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13962 \$263787 \$263532 \$263788 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13963 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263788
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13964 \$263448 \$263530 \$263533 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13965 VSS|anode|cathode|vss \$263530 \$263786 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13966 \$263786 d|z$75 \$263531 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13967 VSS|anode|cathode|vss \$263531 \$263532 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13968 \$263532 \$263447 \$263448 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13969 VSS|anode|cathode|vss \$263534 \$263533 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13970 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$264078
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13971 \$264078 \$263448 \$263534 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13972 VSS|anode|cathode|vss \$263534 R[20]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13973 VSS|anode|cathode|vss cp|i|z$6 \$263535 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13974 VSS|anode|cathode|vss \$263535 \$263449 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13975 \$263536 \$263449 \$263771 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13976 \$263771 \$263537 \$263772 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13977 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263772
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13978 \$263450 \$263535 \$263538 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13979 VSS|anode|cathode|vss \$263535 \$263767 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13980 \$263767 d|z$76 \$263536 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13981 VSS|anode|cathode|vss \$263536 \$263537 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13982 \$263537 \$263449 \$263450 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13983 VSS|anode|cathode|vss \$263539 \$263538 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$13984 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$264103
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$13985 \$264103 \$263450 \$263539 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$13986 VSS|anode|cathode|vss \$263539 R[19]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$13987 VSS|anode|cathode|vss cp|i|z$6 \$263540 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13988 VSS|anode|cathode|vss \$263540 \$263451 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13989 \$263541 \$263451 \$263749 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$13990 \$263749 \$263542 \$263753 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$13991 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263753
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$13992 \$263452 \$263540 \$263543 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$13993 VSS|anode|cathode|vss \$263540 \$263746 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$13994 \$263746 d|z$77 \$263541 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$13995 VSS|anode|cathode|vss \$263541 \$263542 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$13996 \$263542 \$263451 \$263452 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$13997 \$261300 cp|i|z$6 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$13998 VSS|anode|cathode|vss \$261300 \$261301 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$13999 VSS|anode|cathode|vss \$263544 \$263543 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14000 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$264109
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14001 \$264109 \$263452 \$263544 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14002 VSS|anode|cathode|vss \$261300 \$263114 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14003 \$263114 d|z$69 \$261302 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14004 \$261302 \$261301 \$263115 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14005 \$263115 \$261851 \$263116 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14006 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$263116
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14007 \$261851 \$261302 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14008 \$261851 \$261301 \$261304 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14009 \$261304 \$261300 \$263110 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14010 VSS|anode|cathode|vss \$263544 i0|i1|q$12 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14011 \$263545 a2|i|s|zn \$263546 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14012 \$263547 \$263453 \$263545 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14013 VSS|anode|cathode|vss i0|i1|q$9 \$263547 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14014 VSS|anode|cathode|vss i0|i1|q$10 \$263546 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14015 VSS|anode|cathode|vss a2|i|s|zn \$263453 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14016 VSS|anode|cathode|vss \$263545 i0|z$2 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14017 VSS|anode|cathode|vss \$266428 \$266702 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14018 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$267379
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14019 \$267379 \$265341 \$266428 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14020 VSS|anode|cathode|vss \$266428 i0|i1|q$3 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14021 VSS|anode|cathode|vss \$266429 \$266704 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14022 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$267372
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14023 \$267372 \$265345 \$266429 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14024 VSS|anode|cathode|vss \$266429 i0|i1|q$2 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14025 VSS|anode|cathode|vss \$266430 \$266706 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14026 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$267371
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14027 \$267371 \$265349 \$266430 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14028 VSS|anode|cathode|vss \$266430 R[17]|i0|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14029 VSS|anode|cathode|vss \$266431 \$266707 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14030 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$267364
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14031 \$267364 \$265353 \$266431 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14032 VSS|anode|cathode|vss \$266431 i0|i1|q$13 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14033 VSS|anode|cathode|vss \$266432 \$266708 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14034 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$267363
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14035 \$267363 \$265357 \$266432 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14036 VSS|anode|cathode|vss \$266432 i0|i1|q$11 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14037 \$265485 a2|i|s|zn \$265358 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14038 \$265485 i0|i1|q$12 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14039 VSS|anode|cathode|vss i0|i1|q$10 \$265486 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14040 \$265486 \$265359 \$265358 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14041 VSS|anode|cathode|vss a2|i|s|zn \$265359 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14042 VSS|anode|cathode|vss \$265358 i0|z$3 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14043 z$31 cp|i|z$6 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14044 VSS|anode|cathode|vss a1|a2|q \$267362 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14045 \$267362 a1|b|d|z \$265488 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14046 d|z$82 \$265488 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14047 \$265338 cp|i|z$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14048 VSS|anode|cathode|vss \$265338 \$265339 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14049 VSS|anode|cathode|vss \$265338 \$267380 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14050 \$267380 d|z$83 \$265479 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14051 \$265479 \$265339 \$267381 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14052 \$267381 \$266387 \$267382 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14053 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$267382
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14054 \$266387 \$265479 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14055 \$266387 \$265339 \$265341 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14056 \$265341 \$265338 \$266702 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14057 \$265342 cp|i|z$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14058 VSS|anode|cathode|vss \$265342 \$265343 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14059 VSS|anode|cathode|vss \$265342 \$267376 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14060 \$267376 d|z$84 \$265480 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14061 \$265480 \$265343 \$267377 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14062 \$267377 \$266388 \$267378 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14063 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$267378
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14064 \$266388 \$265480 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14065 \$266388 \$265343 \$265345 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14066 \$265345 \$265342 \$266704 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14067 \$265346 cp|i|z$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14068 VSS|anode|cathode|vss \$265346 \$265347 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14069 VSS|anode|cathode|vss \$265346 \$267373 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14070 \$267373 d|z$85 \$265481 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14071 \$265481 \$265347 \$267374 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14072 \$267374 \$266389 \$267375 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14073 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$267375
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14074 \$266389 \$265481 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14075 \$266389 \$265347 \$265349 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14076 \$265349 \$265346 \$266706 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14077 \$265350 cp|i|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14078 VSS|anode|cathode|vss \$265350 \$265351 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14079 VSS|anode|cathode|vss \$265350 \$267368 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14080 \$267368 d|z$79 \$265482 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14081 \$265482 \$265351 \$267369 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14082 \$267369 \$266390 \$267370 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14083 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$267370
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14084 \$266390 \$265482 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14085 \$266390 \$265351 \$265353 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14086 \$265353 \$265350 \$266707 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14087 \$265354 cp|i|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14088 VSS|anode|cathode|vss \$265354 \$265355 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14089 VSS|anode|cathode|vss \$265354 \$267365 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14090 \$267365 d|z$80 \$265484 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14091 \$265484 \$265355 \$267366 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14092 \$267366 \$266391 \$267367 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14093 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$267367
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14094 \$266391 \$265484 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14095 \$266391 \$265355 \$265357 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14096 \$265357 \$265354 \$266708 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14097 \$267880 s|zn$5 \$267881 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14098 \$267882 \$267883 \$267880 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14099 VSS|anode|cathode|vss i0|i1|q$2 \$267882 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14100 VSS|anode|cathode|vss i0|i1|q$1 \$267881 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14101 VSS|anode|cathode|vss s|zn$5 \$267883 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14102 VSS|anode|cathode|vss \$267880 d|z$81 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14103 \$267884 s|zn$5 \$267885 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14104 \$267886 \$267887 \$267884 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14105 VSS|anode|cathode|vss i0|i1|q \$267886 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14106 VSS|anode|cathode|vss i0|i1|q$6 \$267885 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14107 VSS|anode|cathode|vss s|zn$5 \$267887 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14108 VSS|anode|cathode|vss \$267884 d|z$86 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14109 VSS|anode|cathode|vss cp|i|z$7 \$267889 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14110 VSS|anode|cathode|vss \$267889 \$267890 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14111 \$267891 \$267890 \$268104 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14112 \$268104 \$267892 \$268102 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14113 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$268102
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14114 \$267893 \$267889 \$267894 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14115 VSS|anode|cathode|vss \$267889 \$268166 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14116 \$268166 d|z$86 \$267891 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14117 VSS|anode|cathode|vss \$267891 \$267892 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14118 \$267892 \$267890 \$267893 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14119 VSS|anode|cathode|vss \$267895 \$267894 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14120 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$268165
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14121 \$268165 \$267893 \$267895 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14122 VSS|anode|cathode|vss \$267895 i0|i1|q$6 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14123 VSS|anode|cathode|vss cp|i|z$7 \$267896 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14124 VSS|anode|cathode|vss \$267896 \$267897 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14125 \$267898 \$267897 \$268114 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14126 \$268114 \$267899 \$268113 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14127 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$268113
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14128 \$267900 \$267896 \$267901 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14129 VSS|anode|cathode|vss \$267896 \$268164 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14130 \$268164 d|z$88 \$267898 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14131 VSS|anode|cathode|vss \$267898 \$267899 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14132 \$267899 \$267897 \$267900 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14133 VSS|anode|cathode|vss \$267902 \$267901 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14134 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$268163
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14135 \$268163 \$267900 \$267902 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14136 VSS|anode|cathode|vss \$267902 i0|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14137 z$32 cp|i|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14138 VSS|anode|cathode|vss a1|b|d|z \$267904 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14139 \$267904 a1|zn$22 s|zn$5 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14140 s|zn$5 a2|zn$32 \$267904 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14141 \$267905 a2|i|s|zn \$267906 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14142 \$267907 \$267908 \$267905 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14143 VSS|anode|cathode|vss i0|i1|q$13 \$267907 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14144 VSS|anode|cathode|vss a1|i1|q \$267906 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14145 VSS|anode|cathode|vss a2|i|s|zn \$267908 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14146 VSS|anode|cathode|vss \$267905 i0|z$6 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14147 \$267910 a2|i|s|zn \$267911 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14148 \$267912 \$267913 \$267910 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14149 VSS|anode|cathode|vss i0|i1|q$11 \$267912 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14150 VSS|anode|cathode|vss i0|i1|q$13 \$267911 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14151 VSS|anode|cathode|vss a2|i|s|zn \$267913 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14152 VSS|anode|cathode|vss \$267910 i0|z$4 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14153 VSS|anode|cathode|vss a2|q \$268162 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14154 \$268162 a1|b|d|z \$267914 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14155 VSS|anode|cathode|vss \$267914 DOUT_EN|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14156 VSS|anode|cathode|vss i|z$115 \$267916 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14157 VSS|anode|cathode|vss \$267916 cp|i|z$4 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14158 VSS|anode|cathode|vss a1|a2|q$2 \$268161 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14159 \$268161 a1|i0|q$1 a1|zn$21 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14160 \$267917 d|s|zn \$267919 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14161 \$267920 \$267921 \$267917 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14162 VSS|anode|cathode|vss a1|i0|q$1 \$267920 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14163 VSS|anode|cathode|vss DATA|core|i0|i1|p2c \$267919
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3756625p AD=0.244125p
+ PS=2.27u PD=1.53u
M$14164 VSS|anode|cathode|vss d|s|zn \$267921 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14165 VSS|anode|cathode|vss \$267917 d|z$87 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14166 VSS|anode|cathode|vss a1|a2|q$2 \$268160 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14167 \$268160 a1|i0|q$1 \$267923 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14168 VSS|anode|cathode|vss \$267923 a1|a2|a4|z VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14169 VSS|anode|cathode|vss cp|i|z$6 \$267924 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14170 VSS|anode|cathode|vss \$267924 \$267925 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14171 \$267926 \$267925 \$268109 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14172 \$268109 \$267927 \$268111 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14173 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$268111
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14174 \$267928 \$267924 \$267929 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14175 VSS|anode|cathode|vss \$267924 \$268159 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14176 \$268159 a1|b|d|z \$267926 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14177 VSS|anode|cathode|vss \$267926 \$267927 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14178 \$267927 \$267925 \$267928 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14179 VSS|anode|cathode|vss \$267930 \$267929 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14180 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$268158
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14181 \$268158 \$267928 \$267930 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14182 VSS|anode|cathode|vss \$267930 a1|a2|q$1 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14183 a1|b|d|z CEB|a1|core|i|p2c VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14184 VSS|anode|cathode|vss cp|i|z$6 \$267932 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14185 VSS|anode|cathode|vss \$267932 \$267933 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14186 \$267934 \$267933 \$268105 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14187 \$268105 \$267935 \$268106 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14188 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$268106
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14189 \$267936 \$267932 \$267937 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14190 VSS|anode|cathode|vss \$267932 \$268157 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14191 \$268157 d|z$82 \$267934 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14192 VSS|anode|cathode|vss \$267934 \$267935 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14193 \$267935 \$267933 \$267936 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14194 VSS|anode|cathode|vss \$267938 \$267937 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14195 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$268156
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14196 \$268156 \$267936 \$267938 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14197 VSS|anode|cathode|vss \$267938 a1|a2|b|q|s VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14198 \$270063 s|zn$5 \$269998 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14199 \$270063 i0|i1|q$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14200 VSS|anode|cathode|vss i0|i1|q$1 \$270064 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14201 \$270064 \$269910 \$269998 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14202 VSS|anode|cathode|vss s|zn$5 \$269910 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14203 VSS|anode|cathode|vss \$269998 d|z$83 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14204 \$270065 s|zn$5 \$269999 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14205 \$270065 i0|i1|q$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14206 VSS|anode|cathode|vss i0|i1|q$6 \$270066 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14207 \$270066 \$269911 \$269999 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14208 VSS|anode|cathode|vss s|zn$5 \$269911 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14209 VSS|anode|cathode|vss \$269999 d|z$84 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14210 z$33 cp|i|z$7 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14211 cp|i|z$7 \$270000 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$14212 VSS|anode|cathode|vss i|z$115 \$270000 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14213 \$270068 s|zn$5 \$270001 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14214 \$270068 i0|i1|q VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14215 VSS|anode|cathode|vss DATA|core|i0|i1|p2c \$270069
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p
+ AD=0.1890375p PS=2.27u PD=1.335u
M$14216 \$270069 \$269912 \$270001 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14217 VSS|anode|cathode|vss s|zn$5 \$269912 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14218 VSS|anode|cathode|vss \$270001 d|z$88 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14219 \$270070 s|zn$6 \$270002 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14220 \$270070 i0|i1|q$6 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p PS=1.53u PD=2.27u
M$14221 VSS|anode|cathode|vss R[17]|i0|q \$270071 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14222 \$270071 \$269913 \$270002 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14223 VSS|anode|cathode|vss s|zn$6 \$269913 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14224 VSS|anode|cathode|vss \$270002 d|z$85 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14225 VSS|anode|cathode|vss \$270780 \$271740 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14226 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$271797
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14227 \$271797 \$270006 \$270780 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14228 VSS|anode|cathode|vss \$270780 a1|i1|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14229 VSS|anode|cathode|vss \$270782 \$271741 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14230 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$271790
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14231 \$271790 \$270010 \$270782 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14232 VSS|anode|cathode|vss \$270782 DOUT_DAT|c2p|core|i|q
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p
+ PS=4.01u PD=2.53u
M$14233 VSS|anode|cathode|vss \$270784 \$271742 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14234 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$271789
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14235 \$271789 \$270014 \$270784 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14236 VSS|anode|cathode|vss \$270784 a1|i0|q$1 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14237 VSS|anode|cathode|vss \$270786 \$271743 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14238 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$271782
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14239 \$271782 \$270787 \$270786 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14240 VSS|anode|cathode|vss \$270786 a2|i|q$1 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14241 a2|z$13 a2|i|q$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14242 d|z$89 \$270079 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14243 \$271744 a3|zn$10 \$271780 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14244 \$271780 a2|z$13 \$271781 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14245 \$271781 a1|a2|q$1 a1|zn$22 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14246 \$271744 a4|zn$6 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14247 cp|i|z$6 \$270018 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$14248 VSS|anode|cathode|vss i|z$115 \$270018 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14249 VSS|anode|cathode|vss \$270789 \$271745 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14250 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$271775
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14251 \$271775 \$270022 \$270789 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14252 VSS|anode|cathode|vss \$270789 a1|a2|q VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14253 \$270003 cp|i|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14254 VSS|anode|cathode|vss \$270003 \$270004 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14255 VSS|anode|cathode|vss \$270003 \$271794 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14256 \$271794 d|z$90 \$270072 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14257 \$270072 \$270004 \$271795 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14258 \$271795 \$270779 \$271796 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14259 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$271796
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14260 \$270779 \$270072 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14261 \$270779 \$270004 \$270006 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14262 \$270006 \$270003 \$271740 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14263 \$270007 cp|i|z$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14264 VSS|anode|cathode|vss \$270007 \$270008 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14265 VSS|anode|cathode|vss \$270007 \$271791 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14266 \$271791 d|z$91 \$270074 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14267 \$270074 \$270008 \$271792 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14268 \$271792 \$270781 \$271793 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14269 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$271793
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14270 \$270781 \$270074 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14271 \$270781 \$270008 \$270010 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14272 \$270010 \$270007 \$271741 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14273 \$270011 cp|i|z$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14274 VSS|anode|cathode|vss \$270011 \$270012 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14275 VSS|anode|cathode|vss \$270011 \$271786 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14276 \$271786 d|z$87 \$270075 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14277 \$270075 \$270012 \$271787 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14278 \$271787 \$270783 \$271788 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14279 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$271788
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14280 \$270783 \$270075 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14281 \$270783 \$270012 \$270014 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14282 \$270014 \$270011 \$271742 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14283 \$270015 cp|i|z$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14284 VSS|anode|cathode|vss \$270015 \$270016 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14285 VSS|anode|cathode|vss \$270015 \$271783 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14286 \$271783 d|s|zn \$270076 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14287 \$270076 \$270016 \$271784 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14288 \$271784 \$270785 \$271785 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14289 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$271785
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14290 \$270785 \$270076 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14291 \$270785 \$270016 \$270787 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14292 \$270787 \$270015 \$271743 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14293 VSS|anode|cathode|vss a2|q$1 \$271779 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14294 \$271779 a1|b|d|z \$270079 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14295 \$270019 cp|i|z$6 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14296 VSS|anode|cathode|vss \$270019 \$270020 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14297 VSS|anode|cathode|vss \$270019 \$271776 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14298 \$271776 d|z$89 \$270081 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14299 \$270081 \$270020 \$271777 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14300 \$271777 \$270788 \$271778 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14301 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$271778
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14302 \$270788 \$270081 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14303 \$270788 \$270020 \$270022 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14304 \$270022 \$270019 \$271745 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14305 VSS|anode|cathode|vss cp|i|z$7 \$272012 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14306 VSS|anode|cathode|vss \$272012 \$272013 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14307 \$272014 \$272013 \$272573 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14308 \$272573 \$272015 \$272571 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14309 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$272571
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14310 \$272016 \$272012 \$272017 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14311 VSS|anode|cathode|vss \$272012 \$272561 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14312 \$272561 d|z$92 \$272014 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14313 VSS|anode|cathode|vss \$272014 \$272015 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14314 \$272015 \$272013 \$272016 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14315 VSS|anode|cathode|vss \$272018 \$272017 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14316 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$272574
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14317 \$272574 \$272016 \$272018 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14318 VSS|anode|cathode|vss \$272018 a1|a2|q$3 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14319 VSS|anode|cathode|vss a1|a2|q$3 a3|zn$9 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14320 a3|zn$9 a2|q$2 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14321 \$272021 a1|a2|b|q|s \$272022 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.19775p AD=0.244125p PS=1.83u PD=1.53u
M$14322 \$272023 \$272024 \$272021 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14323 VSS|anode|cathode|vss i0|z$6 \$272023 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14324 VSS|anode|cathode|vss i1|zn \$272022 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3756625p AD=0.244125p PS=2.27u PD=1.53u
M$14325 VSS|anode|cathode|vss a1|a2|b|q|s \$272024 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14326 VSS|anode|cathode|vss \$272021 d|z$90 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14327 VSS|anode|cathode|vss cp|i|z$4 \$272025 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14328 VSS|anode|cathode|vss \$272025 \$272026 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14329 \$272027 \$272026 \$272581 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14330 \$272581 \$272028 \$272585 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14331 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$272585
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14332 \$272029 \$272025 \$272030 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14333 VSS|anode|cathode|vss \$272025 \$272582 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14334 \$272582 a2|d|z \$272027 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14335 VSS|anode|cathode|vss \$272027 \$272028 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14336 \$272028 \$272026 \$272029 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14337 VSS|anode|cathode|vss \$272031 \$272030 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14338 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$272586
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14339 \$272586 \$272029 \$272031 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14340 VSS|anode|cathode|vss \$272031 a2|q VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14341 z$34 cp|i|z$5 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14342 VSS|anode|cathode|vss cp|i|z$5 \$272033 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14343 VSS|anode|cathode|vss \$272033 \$272034 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14344 \$272035 \$272034 \$272593 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14345 \$272593 \$272036 \$272592 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14346 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$272592
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14347 \$272037 \$272033 \$272038 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14348 VSS|anode|cathode|vss \$272033 \$272594 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14349 \$272594 d|z$93 \$272035 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14350 VSS|anode|cathode|vss \$272035 \$272036 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14351 \$272036 \$272034 \$272037 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14352 VSS|anode|cathode|vss \$272039 \$272038 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14353 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$272596
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14354 \$272596 \$272037 \$272039 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14355 VSS|anode|cathode|vss \$272039 a1|i0|q$2 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14356 VSS|anode|cathode|vss a2|zn$33 \$272597 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14357 \$272597 a1|i0|q$2 a2|i|s|zn VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14358 VSS|anode|cathode|vss cp|i|z$5 \$272042 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14359 VSS|anode|cathode|vss \$272042 \$272043 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14360 \$272044 \$272043 \$272601 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14361 \$272601 \$272045 \$272600 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14362 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$272600
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14363 \$272046 \$272042 \$272047 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14364 VSS|anode|cathode|vss \$272042 \$272599 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14365 \$272599 d|s|z \$272044 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14366 VSS|anode|cathode|vss \$272044 \$272045 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14367 \$272045 \$272043 \$272046 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14368 VSS|anode|cathode|vss \$272048 \$272047 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14369 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$272602
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14370 \$272602 \$272046 \$272048 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14371 VSS|anode|cathode|vss \$272048 a1|a2|q$4 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14372 VSS|anode|cathode|vss cp|i|z$6 \$272050 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14373 VSS|anode|cathode|vss \$272050 \$272051 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14374 \$272052 \$272051 \$272606 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14375 \$272606 \$272053 \$272605 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14376 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$272605
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14377 \$272054 \$272050 \$272055 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14378 VSS|anode|cathode|vss \$272050 \$272604 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14379 \$272604 d|z$94 \$272052 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14380 VSS|anode|cathode|vss \$272052 \$272053 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14381 \$272053 \$272051 \$272054 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14382 VSS|anode|cathode|vss \$272056 \$272055 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14383 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$272589
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14384 \$272589 \$272054 \$272056 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14385 VSS|anode|cathode|vss \$272056 a2|q$1 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14386 VSS|anode|cathode|vss a1|a2|q a4|zn$6 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14387 a4|zn$6 a1|a2|b|q|s VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14388 VSS|anode|cathode|vss \$275260 \$276108 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14389 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$276127
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14390 \$276127 \$274513 \$275260 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14391 VSS|anode|cathode|vss \$275260 a2|q$2 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14392 d|z$92 \$274521 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14393 d|z$98 \$274522 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14394 d|z$95 \$274523 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14395 a1|z$17 a2|i|q$2 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14396 d|z$91 \$274526 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14397 a2|d|z a2|i|s|zn VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.3955p PS=2.53u PD=2.53u
M$14398 d|z$96 \$274527 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14399 d|z$97 \$274529 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14400 cp|i|z$5 \$274531 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.355125p PS=2.53u PD=2.27u
M$14401 VSS|anode|cathode|vss i|z$115 \$274531 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14402 \$274532 d|s|z \$274514 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.244125p AD=0.19775p PS=1.53u PD=1.83u
M$14403 \$274532 DATA|core|i0|i1|p2c VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.244125p AD=0.3756625p
+ PS=1.53u PD=2.27u
M$14404 VSS|anode|cathode|vss a1|i0|q$2 \$274533 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.505u AS=0.3756625p AD=0.1890375p PS=2.27u PD=1.335u
M$14405 \$274533 \$274424 \$274514 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.1890375p AD=0.19775p PS=1.335u PD=1.83u
M$14406 VSS|anode|cathode|vss d|s|z \$274424 VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.35u AS=0.355125p AD=0.19775p PS=2.27u PD=1.83u
M$14407 VSS|anode|cathode|vss \$274514 d|z$93 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.355125p AD=0.3955p PS=2.27u PD=2.53u
M$14408 \$276109 a3|zn$11 \$276116 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14409 \$276116 a2|zn$34 \$276117 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14410 \$276117 a1|zn$23 a2|zn$33 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14411 \$276109 a4|zn$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14412 d|s|z \$274535 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14413 VSS|anode|cathode|vss a1|a2|q$4 a3|zn$10 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14414 a3|zn$10 a2|q$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14415 VSS|anode|cathode|vss CEB|a1|core|i|p2c d|s|zn VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14416 d|s|zn a1|a2|q$1 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14417 d|z$94 \$274537 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14418 VSS|anode|cathode|vss \$275263 \$276110 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14419 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$276111
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14420 \$276111 \$274518 \$275263 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14421 VSS|anode|cathode|vss \$275263 a2|q$3 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14422 \$274510 cp|i|z$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14423 VSS|anode|cathode|vss \$274510 \$274511 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14424 VSS|anode|cathode|vss \$274510 \$276128 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14425 \$276128 d|z$98 \$274519 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14426 \$274519 \$274511 \$276125 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14427 \$276125 \$274520 \$276126 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14428 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$276126
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14429 \$274520 \$274519 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14430 \$274520 \$274511 \$274513 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14431 \$274513 \$274510 \$276108 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14432 VSS|anode|cathode|vss a1|a2|b|q|s \$276122 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14433 \$276122 a1|b|d|z \$274521 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14434 VSS|anode|cathode|vss a1|a2|q$3 \$276123 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14435 \$276123 a1|b|d|z \$274522 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14436 VSS|anode|cathode|vss a1|a2|q$5 \$276124 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14437 \$276124 a1|b|d|z \$274523 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14438 VSS|anode|cathode|vss a2|d|z \$276121 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14439 \$276121 a1|i1|q \$274526 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14440 VSS|anode|cathode|vss a2|i|q$2 \$276119 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14441 \$276119 a1|b|d|z \$274527 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14442 VSS|anode|cathode|vss a1|a2|q$2 \$276120 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14443 \$276120 a1|b|d|z \$274529 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14444 VSS|anode|cathode|vss a2|i|q$1 \$276118 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14445 \$276118 a1|b|d|z \$274535 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14446 VSS|anode|cathode|vss a1|a2|q$4 \$276115 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14447 \$276115 a1|b|d|z \$274537 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14448 \$274515 cp|i|z$6 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14449 VSS|anode|cathode|vss \$274515 \$274516 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14450 VSS|anode|cathode|vss \$274515 \$276112 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14451 \$276112 d|z$99 \$274538 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14452 \$274538 \$274516 \$276113 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14453 \$276113 \$274539 \$276114 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14454 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$276114
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14455 \$274539 \$274538 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14456 \$274539 \$274516 \$274518 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14457 \$274518 \$274515 \$276110 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14458 VSS|anode|cathode|vss cp|i|z$7 \$276915 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14459 VSS|anode|cathode|vss \$276915 \$276166 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14460 \$276916 \$276166 \$276961 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14461 \$276961 \$276917 \$276959 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14462 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$276959
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14463 \$276167 \$276915 \$276918 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14464 VSS|anode|cathode|vss \$276915 \$276960 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14465 \$276960 d|z$101 \$276916 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14466 VSS|anode|cathode|vss \$276916 \$276917 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14467 \$276917 \$276166 \$276167 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14468 VSS|anode|cathode|vss \$276919 \$276918 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14469 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$277012
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14470 \$277012 \$276167 \$276919 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14471 VSS|anode|cathode|vss \$276919 a1|a2|q$6 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14472 VSS|anode|cathode|vss a2|q$6 \$277011 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14473 \$277011 a1|b|d|z \$276921 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14474 VSS|anode|cathode|vss \$276921 d|z$100 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14475 VSS|anode|cathode|vss a1|a2|q$6 a4|zn$8 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14476 a4|zn$8 a2|q$6 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14477 \$276168 a3|zn$9 \$277013 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14478 \$277013 a2|zn$35 \$277015 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.2905p PS=1.53u PD=1.53u
M$14479 \$277015 a1|z$17 a2|zn$32 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14480 VSS|anode|cathode|vss a4|zn$8 \$276168 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14481 VSS|anode|cathode|vss a1|a2|q$5 a2|zn$35 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14482 a2|zn$35 a2|q$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14483 VSS|anode|cathode|vss cp|i|z$4 \$276924 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14484 VSS|anode|cathode|vss \$276924 \$276169 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14485 \$276925 \$276169 \$276957 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14486 \$276957 \$276926 \$276958 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14487 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$276958
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14488 \$276170 \$276924 \$276927 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14489 VSS|anode|cathode|vss \$276924 \$276956 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14490 \$276956 d|z$96 \$276925 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14491 VSS|anode|cathode|vss \$276925 \$276926 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14492 \$276926 \$276169 \$276170 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14493 VSS|anode|cathode|vss \$276928 \$276927 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14494 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$277014
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14495 \$277014 \$276170 \$276928 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14496 VSS|anode|cathode|vss \$276928 a1|a2|q$2 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14497 VSS|anode|cathode|vss cp|i|z$5 \$276929 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14498 VSS|anode|cathode|vss \$276929 \$276171 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14499 \$276930 \$276171 \$276954 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14500 \$276954 \$276931 \$276955 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14501 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$276955
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14502 \$276172 \$276929 \$276932 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14503 VSS|anode|cathode|vss \$276929 \$276953 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14504 \$276953 d|z$102 \$276930 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14505 VSS|anode|cathode|vss \$276930 \$276931 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14506 \$276931 \$276171 \$276172 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14507 VSS|anode|cathode|vss \$276933 \$276932 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14508 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$277010
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14509 \$277010 \$276172 \$276933 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14510 VSS|anode|cathode|vss \$276933 a2|q$4 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14511 VSS|anode|cathode|vss cp|i|z$5 \$276935 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14512 VSS|anode|cathode|vss \$276935 \$276173 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14513 \$276936 \$276173 \$276951 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14514 \$276951 \$276937 \$276950 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14515 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$276950
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14516 \$276174 \$276935 \$276938 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14517 VSS|anode|cathode|vss \$276935 \$276952 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14518 \$276952 d|z$103 \$276936 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14519 VSS|anode|cathode|vss \$276936 \$276937 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14520 \$276937 \$276173 \$276174 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14521 VSS|anode|cathode|vss \$276939 \$276938 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14522 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$277007
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14523 \$277007 \$276174 \$276939 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14524 VSS|anode|cathode|vss \$276939 a1|a2|q$7 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14525 VSS|anode|cathode|vss cp|i|z$6 \$276941 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14526 VSS|anode|cathode|vss \$276941 \$276175 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14527 \$276942 \$276175 \$276948 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14528 \$276948 \$276943 \$276949 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14529 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$276949
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14530 \$276176 \$276941 \$276944 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14531 VSS|anode|cathode|vss \$276941 \$276947 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14532 \$276947 d|z$104 \$276942 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14533 VSS|anode|cathode|vss \$276942 \$276943 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14534 \$276943 \$276175 \$276176 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14535 VSS|anode|cathode|vss \$276945 \$276944 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14536 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$277006
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14537 \$277006 \$276176 \$276945 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14538 VSS|anode|cathode|vss \$276945 a2|q$5 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14539 d|z$105 \$279198 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14540 d|z$101 \$279200 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14541 VSS|anode|cathode|vss \$279556 \$280217 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14542 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$280585
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14543 \$280585 \$279145 \$279556 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14544 VSS|anode|cathode|vss \$279556 a1|a2|q$5 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14545 VSS|anode|cathode|vss \$279557 \$280218 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14546 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$280595
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14547 \$280595 \$279149 \$279557 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14548 VSS|anode|cathode|vss \$279557 a2|i|q$2 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14549 VSS|anode|cathode|vss \$279558 \$280219 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14550 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$280597
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14551 \$280597 \$279153 \$279558 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14552 VSS|anode|cathode|vss \$279558 a1|a2|q$8 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14553 VSS|anode|cathode|vss \$279559 \$280220 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14554 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$280615
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14555 \$280615 \$279157 \$279559 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14556 VSS|anode|cathode|vss \$279559 a2|q$8 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14557 VSS|anode|cathode|vss a1|a2|q$2 a4|zn$7 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14558 a4|zn$7 a2|q$8 VSS|anode|cathode|vss VSS|anode|cathode|vss sg13_lv_nmos
+ L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14559 VSS|anode|cathode|vss \$279560 \$280221 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14560 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$280625
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14561 \$280625 \$279161 \$279560 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14562 VSS|anode|cathode|vss \$279560 a1|a2|q$9 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14563 d|z$104 \$279208 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14564 d|z$99 \$279209 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.6175p PS=2.53u PD=4.01u
M$14565 VSS|anode|cathode|vss a1|a2|q$6 \$280563 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14566 \$280563 a1|b|d|z \$279198 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14567 VSS|anode|cathode|vss a2|q$2 \$280575 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14568 \$280575 a1|b|d|z \$279200 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14569 \$279142 cp|i|z$7 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14570 VSS|anode|cathode|vss \$279142 \$279143 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14571 VSS|anode|cathode|vss \$279142 \$280581 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14572 \$280581 d|z$100 \$279201 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14573 \$279201 \$279143 \$280579 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14574 \$280579 \$279255 \$280578 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14575 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$280578
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14576 \$279255 \$279201 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14577 \$279255 \$279143 \$279145 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14578 \$279145 \$279142 \$280217 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14579 \$279146 cp|i|z$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14580 VSS|anode|cathode|vss \$279146 \$279147 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14581 VSS|anode|cathode|vss \$279146 \$280592 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14582 \$280592 d|z$106 \$279202 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14583 \$279202 \$279147 \$280590 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14584 \$280590 \$279256 \$280589 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14585 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$280589
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14586 \$279256 \$279202 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14587 \$279256 \$279147 \$279149 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14588 \$279149 \$279146 \$280218 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14589 \$279150 cp|i|z$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14590 VSS|anode|cathode|vss \$279150 \$279151 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14591 VSS|anode|cathode|vss \$279150 \$280603 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14592 \$280603 d|z$97 \$279203 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14593 \$279203 \$279151 \$280601 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14594 \$280601 \$279257 \$280599 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14595 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$280599
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14596 \$279257 \$279203 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14597 \$279257 \$279151 \$279153 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14598 \$279153 \$279150 \$280219 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14599 \$279154 cp|i|z$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14600 VSS|anode|cathode|vss \$279154 \$279155 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14601 VSS|anode|cathode|vss \$279154 \$280604 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14602 \$280604 d|z$107 \$279205 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14603 \$279205 \$279155 \$280612 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14604 \$280612 \$279258 \$280610 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14605 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$280610
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14606 \$279258 \$279205 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14607 \$279258 \$279155 \$279157 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14608 \$279157 \$279154 \$280220 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14609 \$279158 cp|i|z$6 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.19775p AD=0.25625p PS=1.83u PD=1.92u
M$14610 VSS|anode|cathode|vss \$279158 \$279159 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14611 VSS|anode|cathode|vss \$279158 \$280620 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14612 \$280620 d|z$108 \$279207 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14613 \$279207 \$279159 \$280618 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14614 \$280618 \$279259 \$280617 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14615 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$280617
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14616 \$279259 \$279207 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.1954p AD=0.2649375p PS=1.32u PD=2u
M$14617 \$279259 \$279159 \$279161 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14618 \$279161 \$279158 \$280221 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14619 VSS|anode|cathode|vss a1|a2|q$9 \$280622 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14620 \$280622 a1|b|d|z \$279208 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14621 VSS|anode|cathode|vss a2|q$5 \$280635 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14622 \$280635 a1|b|d|z \$279209 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14623 VSS|anode|cathode|vss cp|i|z$7 \$280738 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14624 VSS|anode|cathode|vss \$280738 \$280723 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14625 \$280739 \$280723 \$281235 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14626 \$281235 \$280740 \$281242 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14627 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$281242
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14628 \$280724 \$280738 \$280741 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14629 VSS|anode|cathode|vss \$280738 \$281237 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14630 \$281237 d|z$105 \$280739 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14631 VSS|anode|cathode|vss \$280739 \$280740 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14632 \$280740 \$280723 \$280724 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14633 VSS|anode|cathode|vss \$280742 \$280741 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14634 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$281239
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14635 \$281239 \$280724 \$280742 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14636 VSS|anode|cathode|vss \$280742 a2|q$6 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14637 VSS|anode|cathode|vss cp|i|z$4 \$280743 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14638 VSS|anode|cathode|vss \$280743 \$280725 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.25625p AD=0.19775p PS=1.92u PD=1.83u
M$14639 \$280744 \$280725 \$281247 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1313375p AD=0.101675p PS=1.18u PD=1.075u
M$14640 \$281247 \$280745 \$281246 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.101675p AD=0.101675p PS=1.075u PD=1.075u
M$14641 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$281246
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.245u AS=0.2649375p
+ AD=0.101675p PS=2u PD=1.075u
M$14642 \$280726 \$280743 \$280746 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.245u AS=0.1708875p AD=0.154925p PS=1.32u PD=1.73u
M$14643 VSS|anode|cathode|vss \$280743 \$281243 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.35u AS=0.41975p AD=0.14525p PS=3.31u PD=1.18u
M$14644 \$281243 d|z$95 \$280744 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.35u AS=0.14525p AD=0.1313375p PS=1.18u PD=1.18u
M$14645 VSS|anode|cathode|vss \$280744 \$280745 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.43u AS=0.2649375p AD=0.1954p PS=2u PD=1.32u
M$14646 \$280745 \$280725 \$280726 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.49u AS=0.1954p AD=0.1708875p PS=1.32u PD=1.32u
M$14647 VSS|anode|cathode|vss \$280747 \$280746 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.245u AS=0.3412125p AD=0.154925p PS=2.27u PD=1.73u
M$14648 VSS|anode|cathode|vss RST|a1|b|cdn|core|i|p2c \$281251
+ VSS|anode|cathode|vss sg13_lv_nmos L=0.13u W=0.7u AS=0.3412125p AD=0.2905p
+ PS=2.27u PD=1.53u
M$14649 \$281251 \$280726 \$280747 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14650 VSS|anode|cathode|vss \$280747 a2|q$7 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14651 VSS|anode|cathode|vss a2|q$7 \$281248 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14652 \$281248 a1|b|d|z \$280748 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14653 VSS|anode|cathode|vss \$280748 d|z$106 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14654 VSS|anode|cathode|vss a1|a2|q$8 \$281253 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14655 \$281253 a1|b|d|z \$280749 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14656 VSS|anode|cathode|vss \$280749 d|z$102 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14657 VSS|anode|cathode|vss a2|q$4 \$281252 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14658 \$281252 a1|b|d|z \$280750 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14659 VSS|anode|cathode|vss \$280750 d|z$107 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14660 VSS|anode|cathode|vss a1|a2|q$8 a3|zn$11 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14661 a3|zn$11 a2|q$4 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14662 VSS|anode|cathode|vss a2|q$8 \$281257 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14663 \$281257 a1|b|d|z \$280751 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14664 VSS|anode|cathode|vss \$280751 d|z$103 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14665 VSS|anode|cathode|vss a1|a2|q$7 a2|zn$34 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14666 a2|zn$34 a2|q$3 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14667 VSS|anode|cathode|vss a1|a2|q$7 \$281264 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.635u AS=0.580775p AD=0.263525p PS=3.88u PD=1.465u
M$14668 \$281264 a1|b|d|z \$280752 VSS|anode|cathode|vss sg13_lv_nmos L=0.13u
+ W=0.635u AS=0.263525p AD=0.358775p PS=1.465u PD=2.4u
M$14669 VSS|anode|cathode|vss \$280752 d|z$108 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.6175p AD=0.3955p PS=4.01u PD=2.53u
M$14670 VSS|anode|cathode|vss a1|a2|q$9 a1|zn$23 VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.3955p AD=0.2905p PS=2.53u PD=1.53u
M$14671 a1|zn$23 a2|q$5 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=0.7u AS=0.2905p AD=0.3955p PS=1.53u PD=2.53u
M$14672 CEB|a1|core|i|p2c \$286830 VSS|anode|cathode|vss VSS|anode|cathode|vss
+ sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u PD=6.18u
M$14673 VSSIO|anode|cathode|guard|iovss \$40710 AVDD|anode|cathode|pad|vdd
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$14693 VSSIO|anode|cathode|guard|iovss gate|ngate|o
+ anode|cathode|pad|pad_adc_result_0_pad VSS|anode|cathode|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$14701 VSSIO|anode|cathode|guard|iovss gate|ngate|o$1
+ anode|cathode|pad|pad_adc_result_1_pad VSS|anode|cathode|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$14709 VSSIO|anode|cathode|guard|iovss gate|ngate|o$2
+ anode|cathode|pad|pad_adc_result_2_pad VSS|anode|cathode|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$14717 VSSIO|anode|cathode|guard|iovss gate|ngate|o$3
+ anode|cathode|pad|pad_adc_result_3_pad VSS|anode|cathode|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$14725 VSSIO|anode|cathode|guard|iovss gate|ngate|o$4
+ anode|cathode|pad|pad_adc_result_4_pad VSS|anode|cathode|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$14733 VSSIO|anode|cathode|guard|iovss gate|ngate|o$5
+ anode|cathode|pad|pad_adc_valid_pad VSS|anode|cathode|vss sg13_hv_nmos L=0.6u
+ W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$14741 VSSIO|anode|cathode|guard|iovss gate|ngate|o$6
+ anode|cathode|pad|pad_adc_sample_pad VSS|anode|cathode|vss sg13_hv_nmos
+ L=0.6u W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$14749 \$63424 RESULT[0]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14750 VSS|anode|cathode|vss \$63550 \$63425 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14751 VSS|anode|cathode|vss \$63425 gate|ngate|o VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14752 \$63426 RESULT[0]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14753 VSS|anode|cathode|vss \$63551 \$63427 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14754 VSS|anode|cathode|vss \$63427 gate|o|pgate VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14755 \$63428 RESULT[1]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14756 VSS|anode|cathode|vss \$63553 \$63429 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14757 VSS|anode|cathode|vss \$63429 gate|ngate|o$1 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14758 \$63430 RESULT[1]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14759 VSS|anode|cathode|vss \$63554 \$63431 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14760 VSS|anode|cathode|vss \$63431 gate|o|pgate$1 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14761 \$63432 RESULT[2]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14762 VSS|anode|cathode|vss \$63556 \$63433 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14763 VSS|anode|cathode|vss \$63433 gate|ngate|o$2 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14764 \$63434 RESULT[2]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14765 VSS|anode|cathode|vss \$63557 \$63435 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14766 VSS|anode|cathode|vss \$63435 gate|o|pgate$2 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14767 \$63436 RESULT[3]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14768 VSS|anode|cathode|vss \$63559 \$63437 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14769 VSS|anode|cathode|vss \$63437 gate|ngate|o$3 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14770 \$63438 RESULT[3]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14771 VSS|anode|cathode|vss \$63560 \$63439 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14772 VSS|anode|cathode|vss \$63439 gate|o|pgate$3 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14773 \$63440 RESULT[4]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14774 VSS|anode|cathode|vss \$63562 \$63441 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14775 VSS|anode|cathode|vss \$63441 gate|ngate|o$4 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14776 \$63442 RESULT[4]|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14777 VSS|anode|cathode|vss \$63563 \$63443 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14778 VSS|anode|cathode|vss \$63443 gate|o|pgate$4 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14779 \$63444 VALID|a3|c2p|core|i|z VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14780 VSS|anode|cathode|vss \$63565 \$63445 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14781 VSS|anode|cathode|vss \$63445 gate|ngate|o$5 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14782 \$63446 VALID|a3|c2p|core|i|z VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14783 VSS|anode|cathode|vss \$63566 \$63447 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14784 VSS|anode|cathode|vss \$63447 gate|o|pgate$5 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14785 \$63448 SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14786 VSS|anode|cathode|vss \$63568 \$63449 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14787 VSS|anode|cathode|vss \$63449 gate|ngate|o$6 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14788 \$63450 SAMPLE|a1|c2p|core|i|z VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$14789 VSS|anode|cathode|vss \$63569 \$63451 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$14790 VSS|anode|cathode|vss \$63451 gate|o|pgate$6 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$14791 VSS|anode|cathode|vss core \$64423 VSS|anode|cathode|vss sg13_hv_nmos
+ L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$14792 VSS|anode|cathode|vss core$1 \$64425 VSS|anode|cathode|vss sg13_hv_nmos
+ L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$14793 VSS|anode|cathode|vss core$2 \$90574 VSS|anode|cathode|vss sg13_hv_nmos
+ L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$14794 VSSIO|anode|cathode|guard|iovss \$104193
+ anode|cathode|pad|pad_adc_vrefp_pad VSS|anode|cathode|vss sg13_hv_nmos L=0.6u
+ W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$14814 VSSIO|anode|cathode|guard|iovss in|pin2 gate|out VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.5u W=108u AS=23.22p AD=20.52p PS=131.16u PD=112.56u
M$14820 VSSIO|anode|cathode|guard|iovss in|pin2 VSSIO|anode|cathode|guard|iovss
+ VSS|anode|cathode|vss sg13_hv_nmos L=9.5u W=126u AS=23.94p AD=26.64p
+ PS=131.32u PD=149.92u
M$14840 VSSIO|anode|cathode|guard|iovss gate|out VDD|pad|pin1|supply|vdd
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=756.8u AS=344.608p AD=349.36p
+ PS=931.04u PD=933.2u
M$15012 VSSIO|anode|cathode|guard|iovss \$123893
+ anode|cathode|pad|pad_adc_vrefn_pad VSS|anode|cathode|vss sg13_hv_nmos L=0.6u
+ W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$15032 VSSIO|anode|cathode|guard|iovss \$144910
+ anode|cathode|pad|pad_adc_vin_pad VSS|anode|cathode|vss sg13_hv_nmos L=0.6u
+ W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$15052 VSSIO|anode|cathode|guard|iovss in|pin2$1 gate|out$1
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.5u W=108u AS=23.22p AD=20.52p
+ PS=131.16u PD=112.56u
M$15058 VSSIO|anode|cathode|guard|iovss in|pin2$1
+ VSSIO|anode|cathode|guard|iovss VSS|anode|cathode|vss sg13_hv_nmos L=9.5u
+ W=126u AS=23.94p AD=26.64p PS=131.32u PD=149.92u
M$15078 VSSIO|anode|cathode|guard|iovss gate|out$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply VSS|anode|cathode|vss sg13_hv_nmos
+ L=0.6u W=756.8u AS=344.608p AD=349.36p PS=931.04u PD=933.2u
M$15250 VSSIO|anode|cathode|guard|iovss \$166059
+ anode|cathode|pad|pad_adc_vip_pad VSS|anode|cathode|vss sg13_hv_nmos L=0.6u
+ W=88u AS=40.7p AD=40.7p PS=110.9u PD=110.9u
M$15270 VSSIO|anode|cathode|guard|iovss \$192133 anode|cathode|pad
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15290 VSSIO|anode|cathode|guard|iovss gate|ngate|o$7
+ anode|cathode|pad|pad_miso_pad VSS|anode|cathode|vss sg13_hv_nmos L=0.6u
+ W=35.2u AS=16.676p AD=16.676p PS=47.18u PD=47.18u
M$15298 \$200627 DOUT_DAT|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15299 VSS|anode|cathode|vss \$200626 \$201363 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15300 \$202320 DOUT_DAT|c2p|core|i|q VSS|anode|cathode|vss
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p
+ PS=4.48u PD=2.28u
M$15301 VSS|anode|cathode|vss \$202259 \$202581 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u PD=4.48u
M$15302 VSS|anode|cathode|vss \$201363 gate|ngate|o$7 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$15303 VSS|anode|cathode|vss \$202581 gate|o|pgate$7 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u PD=4.48u
M$15304 VSSIO|anode|cathode|guard|iovss \$220268 anode|cathode|pad$1
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15324 VSS|anode|cathode|vss core$3 \$231093 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$15325 VSSIO|anode|cathode|guard|iovss \$249093 anode|cathode|pad$2
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15345 VSS|anode|cathode|vss core$4 \$258894 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$15346 VSSIO|anode|cathode|guard|iovss \$276913 anode|cathode|pad$3
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15366 VSS|anode|cathode|vss core$5 \$286830 VSS|anode|cathode|vss
+ sg13_hv_nmos L=0.45u W=2.65u AS=0.901p AD=0.901p PS=5.98u PD=5.98u
M$15367 VSSIO|anode|cathode|guard|iovss \$335158 anode|cathode|pad$4
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15387 VSSIO|anode|cathode|guard|iovss \$335159 anode|cathode|pad$5
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15407 VSSIO|anode|cathode|guard|iovss \$335160 anode|cathode|pad$6
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15427 VSSIO|anode|cathode|guard|iovss \$335161 anode|cathode|pad$7
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15447 VSSIO|anode|cathode|guard|iovss \$335162 anode|cathode|pad$8
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15467 VSSIO|anode|cathode|guard|iovss \$335163 anode|cathode|pad$9
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15487 VSSIO|anode|cathode|guard|iovss \$335164 anode|cathode|pad$10
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15507 VSSIO|anode|cathode|guard|iovss \$335165 anode|cathode|pad$11
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15527 VSSIO|anode|cathode|guard|iovss \$335166 anode|cathode|pad$12
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15547 VSSIO|anode|cathode|guard|iovss \$335167 anode|cathode|pad$13
+ VSS|anode|cathode|vss sg13_hv_nmos L=0.6u W=88u AS=40.7p AD=40.7p PS=110.9u
+ PD=110.9u
M$15567 RST|a1|b|cdn|core|i|p2c \$64423 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15568 CLK|core|i|p2c \$64425 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p PS=10.18u PD=10.18u
M$15569 \$63550 RESULT[0]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15570 \$63551 RESULT[0]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15571 \$63553 RESULT[1]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15572 \$63554 RESULT[1]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15573 \$63556 RESULT[2]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15574 \$63557 RESULT[2]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15575 \$63559 RESULT[3]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15576 \$63560 RESULT[3]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15577 \$63562 RESULT[4]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15578 \$63563 RESULT[4]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15579 \$63565 VALID|a3|c2p|core|i|z VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15580 \$63566 VALID|a3|c2p|core|i|z VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15581 \$63568 SAMPLE|a1|c2p|core|i|z VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15582 \$63569 SAMPLE|a1|c2p|core|i|z VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$15583 \$89697 \$90053 \$89697 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$15619 \$89698 \$90054 \$89698 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$15655 \$89699 \$90055 \$89699 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$15691 \$89700 \$90056 \$89700 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$15727 \$89701 \$90057 \$89701 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$15763 \$89702 \$90058 \$89702 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$15799 \$89703 \$90059 \$89703 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$15835 \$89704 \$90060 \$89704 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$15871 \$89705 \$90061 \$89705 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$15907 \$89706 \$90062 \$89706 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$15943 GO|a2|core|p2c \$90574 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p PS=10.18u PD=10.18u
M$16304 \$91546 a2|zn d|zn VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$16305 d|zn a1|z \$91546 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$16306 \$91546 b|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$16307 \$94944 \$95043 \$94944 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16319 \$90053 z$6 \$93030 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16320 \$93030 zn$1 \$93030 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16322 \$90053 zn$1 \$90053 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$16335 \$93031 z$6 \$90053 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16338 \$93031 zn$1 \$93031 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16351 \$93032 z$6 \$90053 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16354 \$93032 zn$1 \$93032 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16355 \$94945 \$95044 \$94945 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1382.4u AS=590.976p AD=590.976p PS=2482.56u PD=2482.56u
M$16367 \$90054 z$6 \$93033 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16368 \$93033 zn$1 \$93033 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16370 \$90054 zn$1 \$90054 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$16383 \$93034 z$6 \$90054 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16386 \$93034 zn$1 \$93034 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16399 \$93035 z$6 \$90054 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16402 \$93035 zn$1 \$93035 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16415 \$90055 z$6 \$93036 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16416 \$93036 zn$1 \$93036 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16418 \$90055 zn$1 \$90055 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$16431 \$93037 z$6 \$90055 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16434 \$93037 zn$1 \$93037 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16447 \$93038 z$6 \$90055 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16450 \$93038 zn$1 \$93038 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16463 \$90056 z$6 \$93039 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16464 \$93039 zn$1 \$93039 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16466 \$90056 zn$1 \$90056 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$16479 \$93040 z$6 \$90056 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16482 \$93040 zn$1 \$93040 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16495 \$93041 z$6 \$90056 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16498 \$93041 zn$1 \$93041 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16511 \$90057 z$6 \$93042 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16512 \$93042 zn$1 \$93042 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16514 \$90057 zn$1 \$90057 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$16527 \$93043 z$6 \$90057 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16530 \$93043 zn$1 \$93043 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16543 \$93044 z$6 \$90057 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16546 \$93044 zn$1 \$93044 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16559 \$90058 z$6 \$93045 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16560 \$93045 zn$1 \$93045 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16562 \$90058 zn$1 \$90058 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$16575 \$93046 z$6 \$90058 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16578 \$93046 zn$1 \$93046 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16591 \$93047 z$6 \$90058 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16594 \$93047 zn$1 \$93047 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16607 \$90059 z$6 \$93048 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16608 \$93048 zn$1 \$93048 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16610 \$90059 zn$1 \$90059 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$16623 \$93049 z$6 \$90059 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16626 \$93049 zn$1 \$93049 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16639 \$93050 z$6 \$90059 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16642 \$93050 zn$1 \$93050 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16655 \$90060 z$6 \$93051 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16656 \$93051 zn$1 \$93051 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16658 \$90060 zn$1 \$90060 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$16671 \$93052 z$6 \$90060 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16674 \$93052 zn$1 \$93052 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16687 \$93053 z$6 \$90060 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16690 \$93053 zn$1 \$93053 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16703 \$90061 z$6 \$93054 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16704 \$93054 zn$1 \$93054 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16706 \$90061 zn$1 \$90061 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$16719 \$93055 z$6 \$90061 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16722 \$93055 zn$1 \$93055 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16735 \$93056 z$6 \$90061 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16738 \$93056 zn$1 \$93056 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16739 \$94946 \$95045 \$94946 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$16751 \$90062 z$6 \$93057 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16752 \$93057 zn$1 \$93057 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16754 \$90062 zn$1 \$90062 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$16767 \$93058 z$6 \$90062 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16770 \$93058 zn$1 \$93058 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16783 \$93059 z$6 \$90062 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$16786 \$93059 zn$1 \$93059 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$16787 VDD|pad|pin1|supply|vdd a1|z$3 \$94578 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$16788 \$94578 a2|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$16789 VDD|pad|pin1|supply|vdd \$94578 d|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$16790 b|zn$1 a1|a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$16791 VDD|pad|pin1|supply|vdd GO|a2|core|p2c b|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$16792 b|zn$1 a2|a3|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$16793 a1|z$1 a1|b|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$16794 a1|z$2 a1|b|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$17155 \$100313 \$100687 \$100313 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$17167 \$95043 z$6 \$98295 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17168 \$98295 zn$1 \$98295 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17170 \$95043 zn$1 \$95043 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17183 \$98296 z$6 \$95043 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17186 \$98296 zn$1 \$98296 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17199 \$98297 z$6 \$95043 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17202 \$98297 zn$1 \$98297 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17215 \$95044 z$4 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=19.2u
+ AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$17216 a2 z$1 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u
+ AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$17218 \$95044 z$1 \$95044 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$17231 VIP|core|padres z$7 \$95044 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=19.2u AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$17232 \$95044 z$3 \$95044 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$17234 VIP|core|padres z$3 VIP|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$17247 VIN|core|padres z$2 \$95044 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=19.2u AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$17248 \$95044 zn \$95044 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$17250 VIN|core|padres zn VIN|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$17299 \$100314 \$100688 \$100314 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=691.2u AS=295.488p AD=295.488p PS=1241.28u PD=1241.28u
M$17587 \$100315 \$100689 \$100315 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$17599 \$95045 z$6 \$98300 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17600 \$98300 zn$1 \$98300 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17602 \$95045 zn$1 \$95045 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$17615 \$98301 z$6 \$95045 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17618 \$98301 zn$1 \$98301 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17631 \$98302 z$6 \$95045 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$17634 \$98302 zn$1 \$98302 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$17635 \$97578 \$97512 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$17636 VDD|pad|pin1|supply|vdd cp|z \$97512 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$17637 \$99205 \$99051 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$17638 VDD|pad|pin1|supply|vdd cp|z$1 \$99051 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$17639 \$97513 \$97512 \$97562 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$17640 \$97562 \$97579 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$17641 \$98709 \$97578 \$97563 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$17642 \$97563 \$97580 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$17643 \$98054 d|z$1 \$97513 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$17644 VDD|pad|pin1|supply|vdd \$97513 \$97579 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$17645 VDD|pad|pin1|supply|vdd \$97578 \$98054 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$17646 \$97579 \$97512 \$98709 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$17647 VDD|pad|pin1|supply|vdd \$98709 \$97580 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$17648 VDD|pad|pin1|supply|vdd \$99205 \$100205 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$17649 \$100205 d|zn$1 \$99052 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$17650 \$99052 \$99051 \$100208 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$17651 VDD|pad|pin1|supply|vdd \$99054 \$100208 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$17652 \$99054 \$99052 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$17653 \$99054 \$99051 \$99053 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$17654 \$99053 \$99205 \$100207 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$17655 VDD|pad|pin1|supply|vdd \$99206 \$100207 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$17656 VDD|pad|pin1|supply|vdd \$99053 \$99206 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$17657 \$96515 a2|zn$1 d|zn$1 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$17658 d|zn$1 a1|z$4 \$96515 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$17659 \$96515 b|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$17660 b|i|q$1 \$97580 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$17661 RESULT[3]|c2p|core|i|q \$99206 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$18022 \$105989 \$106438 \$105989 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$18034 \$100687 z$6 \$104202 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18035 \$104202 zn$1 \$104202 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18037 \$100687 zn$1 \$100687 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$18050 \$104203 z$6 \$100687 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18053 \$104203 zn$1 \$104203 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18066 \$104204 z$6 \$100687 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18069 \$104204 zn$1 \$104204 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18166 \$105990 \$106439 \$105990 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=345.6u AS=147.744p AD=147.744p PS=620.64u PD=620.64u
M$18178 \$100688 z$7 VREFH|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$18179 VREFH|core|padres z$3 VREFH|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$18181 \$100688 z$3 \$100688 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$18194 a2 z$9 \$100688 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u
+ AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$18195 \$100688 z \$100688 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$18197 a2 z a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$18210 a2$1 z$8 \$100688 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$18211 \$100688 z$5 \$100688 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$18213 a2$1 z$5 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$18454 \$105991 \$106440 \$105991 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$18466 \$100689 z$6 \$104207 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18467 \$104207 zn$1 \$104207 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18469 \$100689 zn$1 \$100689 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$18482 \$104208 z$6 \$100689 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18485 \$104208 zn$1 \$104208 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18498 \$104209 z$6 \$100689 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18501 \$104209 zn$1 \$104209 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18502 \$102486 \$102482 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$18503 VDD|pad|pin1|supply|vdd cp|z$1 \$102482 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$18504 \$106441 a2|z$2 b|zn VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$18505 b|zn a1|i|q \$106441 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$18506 \$106441 RST|a1|b|cdn|core|i|p2c VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p
+ PS=2.03u PD=3.53u
M$18507 VDD|pad|pin1|supply|vdd \$102486 \$103538 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$18508 \$103538 d|zn$2 \$102483 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$18509 \$102483 \$102482 \$103537 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$18510 VDD|pad|pin1|supply|vdd \$102487 \$103537 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$18511 \$102487 \$102483 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$18512 \$102487 \$102482 \$102484 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$18513 \$102484 \$102486 \$103536 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$18514 VDD|pad|pin1|supply|vdd \$102761 \$103536 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$18515 VDD|pad|pin1|supply|vdd \$102484 \$102761 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$18516 VDD|pad|pin1|supply|vdd a1|z$3 \$105690 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$18517 \$105690 a2|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$18518 VDD|pad|pin1|supply|vdd \$105690 d|z$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$18519 \$106442 a2|zn$2 d|zn$3 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$18520 d|zn$3 a1|z$5 \$106442 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$18521 \$106442 b|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$18522 RESULT[0]|c2p|core|i|q \$102761 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$18883 a1|z$5 RESULT[2]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$18884 b|zn$2 a1|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$18885 VDD|pad|pin1|supply|vdd a2|i|q b|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$18886 b|zn$2 a1|a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$18887 \$107306 \$106803 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$18888 VDD|pad|pin1|supply|vdd cp|z \$106803 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$18889 \$106804 \$106803 \$107234 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$18890 \$107234 \$107307 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$18891 \$107993 \$107306 \$107230 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$18892 \$107230 \$107783 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$18893 \$107392 d|z \$106804 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$18894 VDD|pad|pin1|supply|vdd \$106804 \$107307 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$18895 VDD|pad|pin1|supply|vdd \$107306 \$107392 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$18896 \$107307 \$106803 \$107993 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$18897 VDD|pad|pin1|supply|vdd \$107993 \$107783 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$18898 b|i|q \$107783 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$18899 a1|z$6 a1|b|i|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$18900 \$110982 \$111646 \$110982 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$18912 \$106438 z$6 \$109162 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18913 \$109162 zn$1 \$109162 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18915 \$106438 zn$1 \$106438 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$18928 \$109163 z$6 \$106438 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18931 \$109163 zn$1 \$109163 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$18944 \$109164 z$6 \$106438 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$18947 \$109164 zn$1 \$109164 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19044 \$110983 \$111647 \$110983 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=172.8u AS=73.872p AD=73.872p PS=310.32u PD=310.32u
M$19056 \$106439 z$7 VREFH|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19059 \$106439 z$3 \$106439 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19072 a2 z$12 \$106439 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19073 \$106439 z$11 \$106439 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19075 a2 z$11 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19088 a2$1 z$10 \$106439 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$19089 \$106439 z$13 \$106439 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19091 a2$1 z$13 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19092 \$110984 \$111648 \$110984 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19140 \$110985 \$111649 \$110985 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19332 \$110986 \$111650 \$110986 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19344 \$106440 z$6 \$109165 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19345 \$109165 zn$1 \$109165 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19347 \$106440 zn$1 \$106440 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$19360 \$109166 z$6 \$106440 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19363 \$109166 zn$1 \$109166 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19376 \$109167 z$6 \$106440 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19379 \$109167 zn$1 \$109167 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19380 \$110275 \$109669 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$19381 VDD|pad|pin1|supply|vdd cp|z \$109669 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$19382 \$109670 \$109669 \$110121 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$19383 \$110121 \$109671 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$19384 \$110890 \$110275 \$110130 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$19385 \$110130 \$110361 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$19386 \$110312 d|z$2 \$109670 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$19387 VDD|pad|pin1|supply|vdd \$109670 \$109671 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$19388 VDD|pad|pin1|supply|vdd \$110275 \$110312 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$19389 \$109671 \$109669 \$110890 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$19390 VDD|pad|pin1|supply|vdd \$110890 \$110361 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$19391 a1|z$8 RESULT[1]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$19392 VDD|pad|pin1|supply|vdd a2|d|zn \$109647 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$19393 \$109647 a1|z$9 d|zn$4 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$19394 d|zn$4 b|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$19395 VDD|pad|pin1|supply|vdd a2|zn$3 \$109641 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$19396 \$109641 a1|z$6 d|zn$5 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$19397 d|zn$5 b|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$19398 b|q \$110361 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$19399 VDD|pad|pin1|supply|vdd i|z$3 \$108731 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$19400 VDD|pad|pin1|supply|vdd \$108731 cp|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$19761 a1|a2|a3|z RST|a1|b|cdn|core|i|p2c VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$19762 VDD|pad|pin1|supply|vdd i|z$3 \$111651 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$19763 VDD|pad|pin1|supply|vdd \$111651 cp|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$19764 \$111966 \$111445 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$19765 VDD|pad|pin1|supply|vdd cp|z$1 \$111445 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$19766 VDD|pad|pin1|supply|vdd \$111966 \$112733 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$19767 \$112733 d|zn \$111446 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$19768 \$111446 \$111445 \$112732 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$19769 VDD|pad|pin1|supply|vdd \$111652 \$112732 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$19770 \$111652 \$111446 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$19771 \$111652 \$111445 \$111447 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$19772 \$111447 \$111966 \$112735 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$19773 VDD|pad|pin1|supply|vdd \$111967 \$112735 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$19774 VDD|pad|pin1|supply|vdd \$111447 \$111967 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$19775 RESULT[4]|c2p|core|i|q \$111967 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$19776 \$116315 \$116455 \$116315 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19788 \$111646 z$6 \$114499 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19789 \$114499 zn$1 \$114499 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19791 \$111646 zn$1 \$111646 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$19804 \$114500 z$6 \$111646 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19807 \$114500 zn$1 \$114500 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19820 \$114501 z$6 \$111646 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19823 \$114501 zn$1 \$114501 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19824 \$116316 \$116456 \$116316 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19872 \$116317 \$116457 \$116317 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19920 \$116318 \$116458 \$116318 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19932 \$111647 z$7 VREFH|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19935 \$111647 z$3 \$111647 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19948 a2 z$14 \$111647 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19949 \$111647 z$15 \$111647 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19951 a2 z$15 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19964 a2$1 z$16 \$111647 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$19965 \$111647 z$19 \$111647 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19967 a2$1 z$19 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19968 \$116319 \$116459 \$116319 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$19980 \$111648 z$7 VREFH|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19983 \$111648 z$3 \$111648 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19996 a2 z$17 \$111648 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$19997 \$111648 z$25 \$111648 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$19999 a2 z$25 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20012 a2$1 z$21 \$111648 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20013 \$111648 z$23 \$111648 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20015 a2$1 z$23 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20016 \$116320 \$116460 \$116320 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20028 \$111649 z$7 VREFH|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20031 \$111649 z$3 \$111649 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20044 a2 z$18 \$111649 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20045 \$111649 zn$2 \$111649 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20047 a2 zn$2 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20060 a2$1 z$18 \$111649 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20063 a2$1 zn$2 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20064 \$116321 \$116461 \$116321 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20112 \$116322 \$116462 \$116322 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20160 \$116323 \$116463 \$116323 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20208 \$116324 \$116464 \$116324 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$20220 \$111650 z$6 \$114502 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20221 \$114502 zn$1 \$114502 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20223 \$111650 zn$1 \$111650 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20236 \$114503 z$6 \$111650 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20239 \$114503 zn$1 \$114503 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20252 \$114504 z$6 \$111650 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20255 \$114504 zn$1 \$114504 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20256 \$114519 \$114505 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20257 VDD|pad|pin1|supply|vdd cp|z \$114505 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20258 VDD|pad|pin1|supply|vdd \$114519 \$115721 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$20259 \$115721 d|z$3 \$114506 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$20260 \$114506 \$114505 \$115716 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$20261 VDD|pad|pin1|supply|vdd \$114520 \$115716 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$20262 \$114520 \$114506 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$20263 \$114520 \$114505 \$114507 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$20264 \$114507 \$114519 \$115717 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$20265 VDD|pad|pin1|supply|vdd \$114892 \$115717 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$20266 VDD|pad|pin1|supply|vdd \$114507 \$114892 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$20267 VDD|pad|pin1|supply|vdd a1|z$7 \$113285 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20268 \$113285 a2|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$20269 VDD|pad|pin1|supply|vdd \$113285 SAMPLE|a1|c2p|core|i|z
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p
+ PS=2.03u PD=3.53u
M$20270 b|i|q$3 \$114892 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$20631 AVDD|anode|cathode|pad|vdd i|z$2 \$126395 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$20633 AVDD|anode|cathode|pad|vdd \$126395 i|z$10 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$20637 AVDD|anode|cathode|pad|vdd i|zn \$124561 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$20639 AVDD|anode|cathode|pad|vdd \$124561 i|z$5 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$20643 \$116455 z$6 \$119711 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20644 \$119711 zn$1 \$119711 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20645 AVDD|anode|cathode|pad|vdd \$126398 \$126182 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$20646 \$126397 i|z$10 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$20647 \$124562 i|z|zn$3 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$20648 AVDD|anode|cathode|pad|vdd \$123895 \$124563 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$20650 \$123895 \$124562 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20651 AVDD|anode|cathode|pad|vdd \$124563 i|z$1 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20652 \$126398 \$126397 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20653 AVDD|anode|cathode|pad|vdd \$126182 i|z$11 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20654 \$116455 zn$1 \$116455 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20655 AVDD|anode|cathode|pad|vdd \$126830 i|z$109 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$20657 AVDD|anode|cathode|pad|vdd i|z$15 \$126830 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20658 \$124565 i|z$6 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$20664 AVDD|anode|cathode|pad|vdd \$124565 i|z|zn AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$20680 \$119712 z$6 \$116455 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20681 AVDD|anode|cathode|pad|vdd i|zn$6 \$126400 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$20687 AVDD|anode|cathode|pad|vdd \$126400 z$7 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$20705 \$119712 zn$1 \$119712 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20706 \$119713 z$6 \$116455 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20709 \$119713 zn$1 \$119713 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20710 \$116456 z$6 \$119714 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20711 \$119714 zn$1 \$119714 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20713 \$116456 zn$1 \$116456 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20714 \$119715 z$6 \$116456 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20717 \$119715 zn$1 \$119715 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20718 \$119716 z$6 \$116456 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20721 \$119716 zn$1 \$119716 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20722 \$116457 z$6 \$119717 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20723 \$119717 zn$1 \$119717 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20725 \$116457 zn$1 \$116457 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20726 \$119718 z$6 \$116457 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20729 \$119718 zn$1 \$119718 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20730 \$119719 z$6 \$116457 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20733 \$119719 zn$1 \$119719 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20734 \$124568 i|z$7 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$20740 AVDD|anode|cathode|pad|vdd \$124568 z$21 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$20756 \$116458 z$6 \$119720 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20757 AVDD|anode|cathode|pad|vdd i|zn$2 \$126401 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$20763 AVDD|anode|cathode|pad|vdd \$126401 i|z|zn$1 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$20779 \$119720 zn$1 \$119720 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20781 \$116458 zn$1 \$116458 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20782 \$119721 z$6 \$116458 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20785 \$119721 zn$1 \$119721 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20786 \$119722 z$6 \$116458 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20789 \$119722 zn$1 \$119722 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20790 \$116459 z$6 \$119723 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20791 \$119723 zn$1 \$119723 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20793 \$116459 zn$1 \$116459 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20794 \$119724 z$6 \$116459 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20795 AVDD|anode|cathode|pad|vdd i|z$16 \$126403 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$20801 AVDD|anode|cathode|pad|vdd \$126403 z$15 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$20819 \$119724 zn$1 \$119724 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20820 \$119725 z$6 \$116459 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20823 \$119725 zn$1 \$119725 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20824 \$116460 z$6 \$119726 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20825 \$119726 zn$1 \$119726 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20827 \$116460 zn$1 \$116460 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20828 \$119727 z$6 \$116460 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20831 \$119727 zn$1 \$119727 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20832 \$119728 z$6 \$116460 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20835 \$119728 zn$1 \$119728 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20836 \$116461 z$6 \$119729 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20837 \$119729 zn$1 \$119729 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20839 \$116461 zn$1 \$116461 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20840 \$119730 z$6 \$116461 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20843 \$119730 zn$1 \$119730 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20844 \$119731 z$6 \$116461 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20847 AVDD|anode|cathode|pad|vdd \$126405 \$126183 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$20848 \$126404 i|zn$8 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$20849 \$119731 zn$1 \$119731 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20850 \$126405 \$126404 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20851 AVDD|anode|cathode|pad|vdd \$126183 i|z$12 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20852 i|zn$1 i|z|zn$1 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$20860 \$116462 z$6 \$119732 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20861 \$119732 zn$1 \$119732 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20863 \$116462 zn$1 \$116462 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20864 \$119733 z$6 \$116462 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20867 \$119733 zn$1 \$119733 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20868 \$119734 z$6 \$116462 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20871 \$119734 zn$1 \$119734 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20872 \$116463 z$6 \$119735 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20873 \$119735 zn$1 \$119735 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20874 AVDD|anode|cathode|pad|vdd \$126410 \$126184 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$20875 \$126408 i|z$13 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$20877 \$126410 \$126408 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20878 AVDD|anode|cathode|pad|vdd \$126184 i|z$14 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20879 \$116463 zn$1 \$116463 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20880 AVDD|anode|cathode|pad|vdd RESULT[1]|c2p|core|i|q \$126412
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p
+ AD=2.8813375p PS=12.07u PD=12.18u
M$20886 AVDD|anode|cathode|pad|vdd \$126412 i|z|zn$2 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$20902 \$119736 z$6 \$116463 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20905 \$119736 zn$1 \$119736 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20906 \$119737 z$6 \$116463 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20909 \$119737 zn$1 \$119737 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20910 AVDD|anode|cathode|pad|vdd \$126415 \$126185 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$20911 \$126414 i|z|zn$5 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$20912 \$116464 z$6 \$119738 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20913 AVDD|anode|cathode|pad|vdd \$124622 i|z$9 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$20915 AVDD|anode|cathode|pad|vdd i|z$8 \$124622 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20916 \$126415 \$126414 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20917 AVDD|anode|cathode|pad|vdd \$126185 i|z$81 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20918 \$119738 zn$1 \$119738 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20920 \$116464 zn$1 \$116464 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$20921 \$119739 z$6 \$116464 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20924 \$119739 zn$1 \$119739 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20925 \$119740 z$6 \$116464 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$20928 \$119740 zn$1 \$119740 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$20929 VDD|pad|pin1|supply|vdd a1|i|q \$120649 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$20930 VDD|pad|pin1|supply|vdd a2|i|q \$120650 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.4185p PS=2.03u PD=2.03u
M$20931 \$120650 \$120649 \$120651 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.4185p AD=0.249p PS=2.03u PD=1.43u
M$20932 \$120651 a1|i|q \$120652 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.249p AD=0.249p PS=1.43u PD=1.43u
M$20933 VDD|pad|pin1|supply|vdd \$120650 \$120652 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.249p PS=2.03u PD=1.43u
M$20934 VDD|pad|pin1|supply|vdd \$120651 a2|a3|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$20935 \$119240 i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.339p AD=0.4185p PS=2.33u PD=2.03u
M$20936 VDD|pad|pin1|supply|vdd \$119240 i|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$20937 a2|zn$4 a1|b|i|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20938 VDD|pad|pin1|supply|vdd a1|a2|a3|z a2|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$20939 a2|zn$4 a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20940 \$126417 \$126076 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20941 VDD|pad|pin1|supply|vdd cp|z$2 \$126076 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20942 \$124570 \$123896 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20943 VDD|pad|pin1|supply|vdd cp|z$2 \$123896 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20944 a2|z$2 a2|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$20945 \$126077 \$126076 \$126338 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$20946 \$126338 \$126186 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$20947 \$126943 \$126417 \$126340 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$20948 \$126340 \$126418 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$20949 \$126658 d|zn$8 \$126077 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$20950 VDD|pad|pin1|supply|vdd \$126077 \$126186 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$20951 VDD|pad|pin1|supply|vdd \$126417 \$126658 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$20952 \$126186 \$126076 \$126943 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$20953 VDD|pad|pin1|supply|vdd \$126943 \$126418 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$20954 a2|z$3 \$120653 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20955 VDD|pad|pin1|supply|vdd b|i|q$2 \$122130 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$20956 \$122130 a1|b|i|q$1 \$120653 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$20957 \$120653 a2|zn$5 \$122130 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20958 VDD|pad|pin1|supply|vdd \$124570 \$125935 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$20959 \$125935 d|zn$7 \$123897 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$20960 \$123897 \$123896 \$125936 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$20961 VDD|pad|pin1|supply|vdd \$123898 \$125936 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$20962 \$123898 \$123897 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$20963 \$123898 \$123896 \$123899 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$20964 \$123899 \$124570 \$125927 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$20965 VDD|pad|pin1|supply|vdd \$124571 \$125927 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$20966 VDD|pad|pin1|supply|vdd \$123899 \$124571 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$20967 VDD|pad|pin1|supply|vdd a2|zn$3 \$119588 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20968 \$119588 a1|z$10 d|zn$6 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$20969 d|zn$6 b|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20970 z$20 i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$20971 VDD|pad|pin1|supply|vdd a1|i|q \$120654 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$20972 \$120654 a2|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$20973 VDD|pad|pin1|supply|vdd \$120654 VALID|a3|c2p|core|i|z
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p
+ PS=2.03u PD=3.53u
M$20974 a1|b|i|q$3 \$126418 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$20975 RESULT[1]|c2p|core|i|q \$124571 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$20976 AVDD|anode|cathode|pad|vdd \$128040 i|z$75 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$20978 AVDD|anode|cathode|pad|vdd i|z \$128040 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$20979 i|z|zn$1 i|zn$1 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$20987 \$127585 i|z$67 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$20993 AVDD|anode|cathode|pad|vdd \$127585 z$3 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21009 \$127586 i|z$17 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21010 AVDD|anode|cathode|pad|vdd \$127588 \$127589 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21011 \$127588 \$127586 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21012 AVDD|anode|cathode|pad|vdd \$127589 i|z$18 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21013 AVDD|anode|cathode|pad|vdd \$128041 i|z$19 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21015 AVDD|anode|cathode|pad|vdd i|z$27 \$128041 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21016 AVDD|anode|cathode|pad|vdd \$128043 i|z$20 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21018 AVDD|anode|cathode|pad|vdd i|z$28 \$128043 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21019 \$127594 i|z$21 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21025 AVDD|anode|cathode|pad|vdd \$127594 z$12 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21041 \$127595 RESULT[4]|c2p|core|i|q AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p
+ AD=2.713175p PS=12.18u PD=12.07u
M$21047 AVDD|anode|cathode|pad|vdd \$127595 i|z|zn$4 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21063 \$127598 i|z$22 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21069 AVDD|anode|cathode|pad|vdd \$127598 a1|i|z|zn
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p
+ PS=32.48u PD=33.98u
M$21085 \$127600 i|z$23 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21086 AVDD|anode|cathode|pad|vdd \$127602 \$127603 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21087 \$127602 \$127600 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21088 AVDD|anode|cathode|pad|vdd \$127603 i|z$32 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21089 i|zn$3 i|z|zn$5 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21097 \$127605 RESULT[2]|c2p|core|i|q AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p
+ AD=2.713175p PS=12.18u PD=12.07u
M$21103 AVDD|anode|cathode|pad|vdd \$127605 i|z|zn$5 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21119 \$127608 i|z$24 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21125 AVDD|anode|cathode|pad|vdd \$127608 z$1 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21141 AVDD|anode|cathode|pad|vdd \$128046 i|z$106 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21143 AVDD|anode|cathode|pad|vdd i|z$29 \$128046 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21144 AVDD|anode|cathode|pad|vdd \$128047 i|z$25 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21146 AVDD|anode|cathode|pad|vdd i|z$12 \$128047 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21147 AVDD|anode|cathode|pad|vdd \$128048 i|z$13 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21149 AVDD|anode|cathode|pad|vdd i|z$30 \$128048 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21150 i|z|zn$6 i|zn$4 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21158 \$127611 i|zn$4 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21159 AVDD|anode|cathode|pad|vdd \$127612 \$127613 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21160 \$127612 \$127611 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21161 AVDD|anode|cathode|pad|vdd \$127613 i|z$8 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21162 i|z|zn$3 i|zn$5 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21170 VDD|pad|pin1|supply|vdd i|z$31 \$127614 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$21171 VDD|pad|pin1|supply|vdd \$127614 i|z$26 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$21172 VDD|pad|pin1|supply|vdd CLK|core|i|p2c \$127616 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$21173 VDD|pad|pin1|supply|vdd \$127616 i|z$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$21174 i|zn$5 i|z|zn$3 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21182 i|zn$6 i|z|zn AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21190 AVDD|anode|cathode|pad|vdd a2|z$5 \$129460 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21191 \$129460 a1|z$12 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=0.996p AD=0.996p PS=4.06u PD=4.06u
M$21194 AVDD|anode|cathode|pad|vdd \$129460 i|z$6 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$21198 AVDD|anode|cathode|pad|vdd \$129462 \$129463 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21199 \$129461 i|z$38 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21200 \$129462 \$129461 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21201 AVDD|anode|cathode|pad|vdd \$129463 i|z$28 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21202 AVDD|anode|cathode|pad|vdd \$130202 i|z$33 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21204 AVDD|anode|cathode|pad|vdd i|z$42 \$130202 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21205 AVDD|anode|cathode|pad|vdd i|z$43 \$129465 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21207 AVDD|anode|cathode|pad|vdd \$129465 a2|z$4 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$21211 AVDD|anode|cathode|pad|vdd \$129468 \$129469 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21212 \$129467 i|z|zn$8 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21213 \$129468 \$129467 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21214 AVDD|anode|cathode|pad|vdd \$129469 i|z$34 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21215 AVDD|anode|cathode|pad|vdd \$129472 \$129473 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21216 \$129471 i|z$39 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21217 \$129472 \$129471 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21218 AVDD|anode|cathode|pad|vdd \$129473 i|z$35 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21219 AVDD|anode|cathode|pad|vdd \$130205 i|z$36 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21221 AVDD|anode|cathode|pad|vdd i|z$44 \$130205 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21222 AVDD|anode|cathode|pad|vdd i|z$45 \$129476 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21228 AVDD|anode|cathode|pad|vdd \$129476 z$9 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21244 AVDD|anode|cathode|pad|vdd i|z$46 \$129477 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21250 AVDD|anode|cathode|pad|vdd \$129477 z AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21266 AVDD|anode|cathode|pad|vdd i|z|zn$1 \$129478 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=3.205u AS=1.569325p AD=1.389325p PS=7.59u PD=6.09u
M$21269 AVDD|anode|cathode|pad|vdd \$129478 i|z$24 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=3.984p AD=4.164p PS=16.24u PD=17.74u
M$21277 AVDD|anode|cathode|pad|vdd i|z$5 \$129479 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21283 AVDD|anode|cathode|pad|vdd \$129479 a1|z$11 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21299 AVDD|anode|cathode|pad|vdd i|z$47 \$129481 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21305 AVDD|anode|cathode|pad|vdd \$129481 z$13 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21321 AVDD|anode|cathode|pad|vdd \$129483 \$129484 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21322 \$129482 i|z$25 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21323 \$129483 \$129482 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21324 AVDD|anode|cathode|pad|vdd \$129484 i|z$30 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21325 i|z|zn$2 i|zn$8 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21333 AVDD|anode|cathode|pad|vdd i|z$48 \$129485 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21339 AVDD|anode|cathode|pad|vdd \$129485 z$14 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21355 AVDD|anode|cathode|pad|vdd \$129487 \$129488 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21356 \$129486 a2|i|z AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21357 \$129487 \$129486 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21358 AVDD|anode|cathode|pad|vdd \$129488 i|z$2 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21359 AVDD|anode|cathode|pad|vdd \$129490 \$129491 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21360 \$129489 i|z$113 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21361 \$129490 \$129489 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21362 AVDD|anode|cathode|pad|vdd \$129491 i|z$29 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21363 z$6 \$130446 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$21364 i|zn$4 i|z|zn$6 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21372 i|z|zn$5 i|zn$3 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21380 i|zn$7 i|zn$2 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21388 AVDD|anode|cathode|pad|vdd \$129494 \$129495 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21389 \$129493 i|z$59 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21390 \$129494 \$129493 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21391 AVDD|anode|cathode|pad|vdd \$129495 i|z$37 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21392 AVDD|anode|cathode|pad|vdd \$130212 i|z$7 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21394 AVDD|anode|cathode|pad|vdd i|z$14 \$130212 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21395 AVDD|anode|cathode|pad|vdd RESULT[3]|c2p|core|i|q \$129497
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p
+ AD=2.8813375p PS=12.07u PD=12.18u
M$21401 AVDD|anode|cathode|pad|vdd \$129497 i|z|zn$7 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21417 a2|zn a1|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21418 VDD|pad|pin1|supply|vdd a1|a2|a3|z a2|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$21419 a2|zn a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21420 \$129355 cp|i|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.339p AD=0.4185p PS=2.33u PD=2.03u
M$21421 VDD|pad|pin1|supply|vdd \$129355 cp|z$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$21422 \$131975 a2$1 a1|c|i|zn AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$21426 AVDD|anode|cathode|pad|vdd a1|z$11 \$131975 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$21430 AVDD|anode|cathode|pad|vdd a2|b|z a1|c|i|zn AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=21.6u AS=9.144p AD=9.144p PS=38.04u PD=38.04u
M$21434 AVDD|anode|cathode|pad|vdd a1|c|i|zn$1 a1|c|i|zn
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=21.6u AS=8.964p AD=9.684p
+ PS=36.54u PD=42.54u
M$21438 \$131976 a2$1 a1|c|i|zn AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$21442 AVDD|anode|cathode|pad|vdd a1|z$11 \$131976 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$21454 \$131977 a2$1 a1|c|i|zn AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$21458 AVDD|anode|cathode|pad|vdd a1|z$11 \$131977 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$21470 \$131978 a2$1 a1|c|i|zn AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$21474 AVDD|anode|cathode|pad|vdd a1|z$11 \$131978 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$21486 AVDD|anode|cathode|pad|vdd a2|b|z a1|c|i|zn$1
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=21.6u AS=9.144p AD=9.144p
+ PS=38.04u PD=38.04u
M$21487 a1|c|i|zn$1 a1|c|i|zn AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=21.6u AS=8.964p AD=9.684p
+ PS=36.54u PD=42.54u
M$21490 AVDD|anode|cathode|pad|vdd \$131123 z$22 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21492 AVDD|anode|cathode|pad|vdd i|z$55 \$131123 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21493 \$130777 i|z$33 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21494 AVDD|anode|cathode|pad|vdd \$130749 \$130778 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21495 \$130749 \$130777 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21496 AVDD|anode|cathode|pad|vdd \$130778 i|z$27 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21497 \$130779 i|z$40 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21503 AVDD|anode|cathode|pad|vdd \$130779 z$23 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21519 \$130781 i|zn$11 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21520 AVDD|anode|cathode|pad|vdd \$130750 \$130782 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21521 \$130750 \$130781 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21522 AVDD|anode|cathode|pad|vdd \$130782 i|z$56 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21523 i|zn$8 i|z|zn$2 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21531 \$130784 i|z$49 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21537 AVDD|anode|cathode|pad|vdd \$130784 z$17 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21553 \$130785 i|z$51 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21554 AVDD|anode|cathode|pad|vdd \$130751 \$130786 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21555 \$130751 \$130785 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21556 AVDD|anode|cathode|pad|vdd \$130786 i|z$62 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21557 \$130787 i|z$24 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21563 AVDD|anode|cathode|pad|vdd \$130787 z$1 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21579 \$130788 i|z$36 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21580 AVDD|anode|cathode|pad|vdd \$130752 \$130789 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21581 \$130752 \$130788 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21582 AVDD|anode|cathode|pad|vdd \$130789 i|z$52 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21583 \$130790 i|z$53 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21584 AVDD|anode|cathode|pad|vdd \$130754 \$130791 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21585 \$130754 \$130790 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21586 AVDD|anode|cathode|pad|vdd \$130791 i|z$57 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21587 \$131746 VALID|a3|c2p|core|i|z AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=3.984p
+ PS=17.74u PD=16.24u
M$21595 \$131746 a2|i|z \$131980 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=9.6u AS=3.984p AD=4.164p PS=16.24u PD=17.74u
M$21603 \$131980 SAMPLE|a1|c2p|core|i|z i|zn$9 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21611 a1|i|z|zn i|zn AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=7.2u AS=3.168p AD=3.168p PS=13.68u PD=13.68u
M$21617 z$18 \$130755 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$21618 i|zn$10 i|z|zn$7 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21626 \$130795 i|z|zn$2 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21627 AVDD|anode|cathode|pad|vdd \$130756 \$130796 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21628 \$130756 \$130795 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21629 AVDD|anode|cathode|pad|vdd \$130796 i|z$42 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21630 AVDD|anode|cathode|pad|vdd \$131124 i|z$58 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21632 AVDD|anode|cathode|pad|vdd i|z$35 \$131124 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21633 AVDD|anode|cathode|pad|vdd \$131125 i|z$59 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21635 AVDD|anode|cathode|pad|vdd i|z$1 \$131125 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21636 AVDD|anode|cathode|pad|vdd \$131126 i|z$48 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21638 AVDD|anode|cathode|pad|vdd i|z$57 \$131126 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21639 \$130799 i|z|zn$6 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21640 AVDD|anode|cathode|pad|vdd \$130757 \$130800 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21641 \$130757 \$130799 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21642 AVDD|anode|cathode|pad|vdd \$130800 i|z$114 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21643 \$130801 i|z$54 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21644 AVDD|anode|cathode|pad|vdd \$130759 \$130802 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21645 \$130759 \$130801 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21646 AVDD|anode|cathode|pad|vdd \$130802 i|z AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21647 \$131519 \$131519 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$21648 \$130803 i|z$41 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21649 AVDD|anode|cathode|pad|vdd \$130760 \$130804 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21650 \$130760 \$130803 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21651 AVDD|anode|cathode|pad|vdd \$130804 i|z$60 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21652 \$130806 i|zn$9 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=3.205u AS=1.569325p AD=1.389325p PS=7.59u PD=6.09u
M$21655 AVDD|anode|cathode|pad|vdd \$130806 i|z$22 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=3.984p AD=4.164p PS=16.24u PD=17.74u
M$21663 AVDD|anode|cathode|pad|vdd \$131127 i|z$54 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21665 AVDD|anode|cathode|pad|vdd i|z$37 \$131127 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21666 i|zn$2 SAMPLE|a1|c2p|core|i|z AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p
+ PS=17.74u PD=17.74u
M$21674 AVDD|anode|cathode|pad|vdd i|z$11 \$130807 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21676 AVDD|anode|cathode|pad|vdd \$130807 i|z$23 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$21680 \$130808 i|z$26 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$21686 AVDD|anode|cathode|pad|vdd \$130808 a2|i|z AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21702 VDD|pad|pin1|supply|vdd CLK|core|i|p2c \$130809 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$21703 VDD|pad|pin1|supply|vdd \$130809 i|z$61 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$21704 VDD|pad|pin1|supply|vdd i|z$61 \$130811 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$21705 VDD|pad|pin1|supply|vdd \$130811 i|z$31 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$21706 a2|z$1 \$131128 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21707 VDD|pad|pin1|supply|vdd b|q \$131981 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$21708 \$131981 a1|b|i|q$2 \$131128 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$21709 \$131128 a2|zn$5 \$131981 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21710 \$130812 \$130761 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21711 VDD|pad|pin1|supply|vdd cp|z$2 \$130761 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21712 RESULT[2]|c2p|core|i|q \$131129 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$21713 a2$1 z$7 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=3.6u
+ AS=2.034p AD=2.034p PS=13.98u PD=13.98u
M$21714 a2 z$3 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.8u
+ AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21716 a2$1 z$3 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.8u
+ AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$21725 \$132451 a2 a1|c|i|zn$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$21729 AVDD|anode|cathode|pad|vdd a1|z$11 \$132451 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$21741 \$132453 a2 a1|c|i|zn$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$21745 AVDD|anode|cathode|pad|vdd a1|z$11 \$132453 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$21757 \$132454 a2 a1|c|i|zn$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$21761 AVDD|anode|cathode|pad|vdd a1|z$11 \$132454 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$21773 \$132455 a2 a1|c|i|zn$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.172p AD=2.172p PS=9.62u PD=9.62u
M$21777 AVDD|anode|cathode|pad|vdd a1|z$11 \$132455 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=2.172p AD=1.992p PS=9.62u PD=8.12u
M$21793 \$132448 a1|c|i|zn AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.36u AS=0.2034p
+ AD=0.2129625p PS=1.85u PD=1.415u
M$21794 AVDD|anode|cathode|pad|vdd \$132448 i|z$65 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.585u AS=0.2129625p AD=0.330525p PS=1.415u PD=2.3u
M$21795 AVDD|anode|cathode|pad|vdd a1|c|i|zn$1 \$130774
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.36u AS=0.2129625p
+ AD=0.2034p PS=1.415u PD=1.85u
M$21796 AVDD|anode|cathode|pad|vdd \$130774 i|z$55 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.585u AS=0.2129625p AD=0.330525p PS=1.415u PD=2.3u
M$21797 AVDD|anode|cathode|pad|vdd \$133160 a2|a3|z AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21799 AVDD|anode|cathode|pad|vdd i|z$65 \$133160 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21800 AVDD|anode|cathode|pad|vdd a2|z$4 \$132456 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21801 \$132456 a1|i|z|zn AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u AS=0.996p AD=0.996p
+ PS=4.06u PD=4.06u
M$21804 AVDD|anode|cathode|pad|vdd \$132456 i|z$66 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$21808 AVDD|anode|cathode|pad|vdd i|z$74 \$132458 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21814 AVDD|anode|cathode|pad|vdd \$132458 z$11 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21830 z$24 \$133352 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$21831 i|z|zn$7 i|zn$10 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21839 AVDD|anode|cathode|pad|vdd i|z$75 \$132459 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21845 AVDD|anode|cathode|pad|vdd \$132459 z$25 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21861 AVDD|anode|cathode|pad|vdd i|z|zn \$132461 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=3.205u AS=1.569325p AD=1.389325p PS=7.59u PD=6.09u
M$21864 AVDD|anode|cathode|pad|vdd \$132461 i|z$67 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=3.984p AD=4.164p PS=16.24u PD=17.74u
M$21872 AVDD|anode|cathode|pad|vdd \$132464 \$132465 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21873 \$132463 i|z|zn$4 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21874 \$132464 \$132463 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21875 AVDD|anode|cathode|pad|vdd \$132465 i|z$63 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21876 AVDD|anode|cathode|pad|vdd i|z$76 \$132466 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21882 AVDD|anode|cathode|pad|vdd \$132466 z$10 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21898 AVDD|anode|cathode|pad|vdd i|z$58 \$132467 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21904 AVDD|anode|cathode|pad|vdd \$132467 z$19 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21920 AVDD|anode|cathode|pad|vdd \$133164 i|z$74 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21922 AVDD|anode|cathode|pad|vdd i|z$101 \$133164 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21923 AVDD|anode|cathode|pad|vdd \$132469 \$132470 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21924 \$132468 i|zn$10 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21925 \$132469 \$132468 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21926 AVDD|anode|cathode|pad|vdd \$132470 i|z$68 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21927 i|zn$11 i|z|zn$8 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$21935 z$2 \$133354 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$21936 AVDD|anode|cathode|pad|vdd b|i|q \$132473 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21942 AVDD|anode|cathode|pad|vdd \$132473 i|z|zn$8 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$21958 AVDD|anode|cathode|pad|vdd \$133168 i|z$69 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21960 AVDD|anode|cathode|pad|vdd i|z$77 \$133168 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21961 AVDD|anode|cathode|pad|vdd \$132476 \$132477 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21962 \$132475 i|z$72 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21963 \$132476 \$132475 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21964 AVDD|anode|cathode|pad|vdd \$132477 i|z$64 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21965 AVDD|anode|cathode|pad|vdd \$132479 \$132480 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21966 \$132478 i|z$69 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21967 \$132479 \$132478 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21968 AVDD|anode|cathode|pad|vdd \$132480 i|z$70 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21969 AVDD|anode|cathode|pad|vdd \$133170 i|z$46 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21971 AVDD|anode|cathode|pad|vdd i|z$79 \$133170 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21972 AVDD|anode|cathode|pad|vdd \$132483 \$132484 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21973 \$132482 i|z$103 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21974 \$132483 \$132482 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21975 AVDD|anode|cathode|pad|vdd \$132484 i|z$112 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21976 AVDD|anode|cathode|pad|vdd \$132486 \$132487 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$21977 \$132485 i|z$73 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$21978 \$132486 \$132485 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$21979 AVDD|anode|cathode|pad|vdd \$132487 i|z$71 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21980 AVDD|anode|cathode|pad|vdd \$133171 i|z$16 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$21982 AVDD|anode|cathode|pad|vdd i|z$80 \$133171 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$21983 AVDD|anode|cathode|pad|vdd b|i|q$1 \$132489 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$21989 AVDD|anode|cathode|pad|vdd \$132489 i|z|zn$9 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22005 \$132491 \$132446 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22006 VDD|pad|pin1|supply|vdd cp|z$1 \$132446 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22007 \$132447 \$132446 \$132714 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22008 \$132714 \$132492 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$22009 \$133356 \$132491 \$132715 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$22010 \$132715 \$132493 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$22011 \$132724 d|zn$4 \$132447 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$22012 VDD|pad|pin1|supply|vdd \$132447 \$132492 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$22013 VDD|pad|pin1|supply|vdd \$132491 \$132724 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$22014 \$132492 \$132446 \$133356 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$22015 VDD|pad|pin1|supply|vdd \$133356 \$132493 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$22016 a1|i|q$1 \$132493 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22017 VDD|pad|pin1|supply|vdd \$130812 \$132072 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$22018 \$132072 d|zn$3 \$130762 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$22019 \$130762 \$130761 \$132073 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22020 VDD|pad|pin1|supply|vdd \$130813 \$132073 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22021 \$130813 \$130762 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$22022 \$130813 \$130761 \$130763 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$22023 \$130763 \$130812 \$132068 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$22024 VDD|pad|pin1|supply|vdd \$131129 \$132068 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$22025 VDD|pad|pin1|supply|vdd \$130763 \$131129 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$22026 AVDD|anode|cathode|pad|vdd i|zn$1 \$135445 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22032 AVDD|anode|cathode|pad|vdd \$135445 z$4 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22048 z$26 \$133781 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22049 \$134212 \$134212 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22050 i|z|zn i|zn$6 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22058 \$133929 i|z$66 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22064 AVDD|anode|cathode|pad|vdd \$133929 a2|b|z AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22080 \$134213 \$134213 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22081 AVDD|anode|cathode|pad|vdd \$135447 \$135382 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22082 \$135446 i|z$9 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22083 \$133930 i|z$83 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22084 AVDD|anode|cathode|pad|vdd \$133783 \$133931 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22085 \$135447 \$135446 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22086 AVDD|anode|cathode|pad|vdd \$135382 i|z$97 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22087 \$133783 \$133930 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22088 AVDD|anode|cathode|pad|vdd \$133931 i|z$86 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22089 AVDD|anode|cathode|pad|vdd \$136356 i|z$50 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22091 AVDD|anode|cathode|pad|vdd i|z$62 \$136356 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22092 \$133933 i|zn$7 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=3.205u AS=1.569325p AD=1.389325p PS=7.59u PD=6.09u
M$22095 AVDD|anode|cathode|pad|vdd \$133933 a1|z$12 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=3.984p AD=4.164p PS=16.24u PD=17.74u
M$22103 AVDD|anode|cathode|pad|vdd \$133935 i|z$83 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22105 AVDD|anode|cathode|pad|vdd i|z$97 \$133935 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22106 AVDD|anode|cathode|pad|vdd \$133936 i|z$87 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22108 AVDD|anode|cathode|pad|vdd i|z$102 \$133936 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22109 \$133938 a1|i|z|zn AVDD|anode|cathode|pad|vdd
+ AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p
+ PS=3.53u PD=2.03u
M$22110 AVDD|anode|cathode|pad|vdd \$133784 \$133939 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22111 \$135448 \$135448 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22112 \$133784 \$133938 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22113 AVDD|anode|cathode|pad|vdd \$133939 i|z$43 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22114 \$133940 i|z$98 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22120 AVDD|anode|cathode|pad|vdd \$133940 z$8 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22136 AVDD|anode|cathode|pad|vdd i|zn$1 \$135449 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22142 AVDD|anode|cathode|pad|vdd \$135449 z$4 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22158 AVDD|anode|cathode|pad|vdd \$136357 i|z$21 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22160 AVDD|anode|cathode|pad|vdd i|z$86 \$136357 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22161 \$133941 i|z$84 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22162 AVDD|anode|cathode|pad|vdd \$133786 \$133942 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22163 AVDD|anode|cathode|pad|vdd \$135451 \$135383 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22164 \$135450 i|z|zn$9 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22165 \$133786 \$133941 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22166 AVDD|anode|cathode|pad|vdd \$133942 i|z$80 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22167 \$135451 \$135450 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22168 AVDD|anode|cathode|pad|vdd \$135383 i|z$96 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22169 \$133943 i|zn$3 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22170 AVDD|anode|cathode|pad|vdd \$133787 \$133944 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22171 \$133787 \$133943 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22172 AVDD|anode|cathode|pad|vdd \$133944 i|z$88 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22173 AVDD|anode|cathode|pad|vdd b|i|q$3 \$135452 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.6065125p AD=2.8813375p PS=12.07u PD=12.18u
M$22179 AVDD|anode|cathode|pad|vdd \$135452 i|z|zn$3 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22195 AVDD|anode|cathode|pad|vdd \$133946 i|z$82 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22197 AVDD|anode|cathode|pad|vdd i|z$89 \$133946 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22198 i|zn$12 i|z|zn$4 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22206 AVDD|anode|cathode|pad|vdd i|z$32 \$133949 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22208 AVDD|anode|cathode|pad|vdd \$133949 a2|z$5 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=4.8u AS=1.992p AD=2.172p PS=8.12u PD=9.62u
M$22212 AVDD|anode|cathode|pad|vdd \$135454 \$135384 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22213 \$135453 i|z$19 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22214 \$135454 \$135453 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22215 AVDD|anode|cathode|pad|vdd \$135384 i|z$105 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22216 AVDD|anode|cathode|pad|vdd \$135458 \$135385 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22217 \$135456 i|z$106 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22218 i|zn a1|i|z|zn AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=7.2u AS=3.168p AD=3.168p PS=13.68u PD=13.68u
M$22224 \$135458 \$135456 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22225 AVDD|anode|cathode|pad|vdd \$135385 i|z$101 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22226 AVDD|anode|cathode|pad|vdd \$133950 i|z$17 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22228 AVDD|anode|cathode|pad|vdd i|z$81 \$133950 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22229 \$133951 i|z$50 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22230 AVDD|anode|cathode|pad|vdd \$133788 \$133952 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22231 AVDD|anode|cathode|pad|vdd \$136358 i|z$103 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22233 AVDD|anode|cathode|pad|vdd i|z$56 \$136358 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22234 \$133788 \$133951 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22235 AVDD|anode|cathode|pad|vdd \$133952 i|z$79 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22236 z$27 \$136577 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22237 \$133953 i|z$87 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22243 AVDD|anode|cathode|pad|vdd \$133953 z$16 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22259 AVDD|anode|cathode|pad|vdd \$136359 i|z$38 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22261 AVDD|anode|cathode|pad|vdd i|z$88 \$136359 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22262 i|zn$13 i|z|zn$9 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22270 AVDD|anode|cathode|pad|vdd \$136360 i|z$107 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22272 AVDD|anode|cathode|pad|vdd i|z$94 \$136360 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22273 \$135460 \$135460 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22274 AVDD|anode|cathode|pad|vdd \$133954 i|z$39 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22276 AVDD|anode|cathode|pad|vdd i|z$18 \$133954 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22277 AVDD|anode|cathode|pad|vdd \$133955 i|z$41 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22279 AVDD|anode|cathode|pad|vdd i|z$34 \$133955 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22280 AVDD|anode|cathode|pad|vdd \$135463 \$135386 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22281 \$135461 i|z$108 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22282 \$135463 \$135461 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22283 AVDD|anode|cathode|pad|vdd \$135386 i|z$99 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22284 \$133956 i|z$78 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22290 AVDD|anode|cathode|pad|vdd \$133956 z$5 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22306 AVDD|anode|cathode|pad|vdd \$135466 \$135387 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22307 \$135464 i|z$109 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22308 \$135466 \$135464 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22309 AVDD|anode|cathode|pad|vdd \$135387 i|z$77 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22310 i|z|zn$4 i|zn$12 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22318 AVDD|anode|cathode|pad|vdd \$136361 i|z$110 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22320 AVDD|anode|cathode|pad|vdd i|z$104 \$136361 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22321 AVDD|anode|cathode|pad|vdd \$133957 i|z$45 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22323 AVDD|anode|cathode|pad|vdd i|z$90 \$133957 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22324 i|z|zn$8 i|zn$11 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22332 AVDD|anode|cathode|pad|vdd \$133959 i|z$91 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22334 AVDD|anode|cathode|pad|vdd i|z$92 \$133959 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22335 AVDD|anode|cathode|pad|vdd \$136362 i|z$73 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22337 AVDD|anode|cathode|pad|vdd i|z$68 \$136362 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22338 AVDD|anode|cathode|pad|vdd \$133962 i|z$98 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22340 AVDD|anode|cathode|pad|vdd i|z$99 \$133962 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22341 \$133964 b|i|q$2 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22347 AVDD|anode|cathode|pad|vdd \$133964 i|z|zn$6 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22363 AVDD|anode|cathode|pad|vdd \$136363 i|z$108 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22365 AVDD|anode|cathode|pad|vdd i|z$64 \$136363 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22366 AVDD|anode|cathode|pad|vdd \$135469 \$135388 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22367 \$135468 i|z$110 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22368 \$135469 \$135468 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22369 AVDD|anode|cathode|pad|vdd \$135388 i|z$92 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22370 AVDD|anode|cathode|pad|vdd \$135471 \$135389 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22371 \$135470 i|z$91 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22372 \$135471 \$135470 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22373 AVDD|anode|cathode|pad|vdd \$135389 i|z$90 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22374 AVDD|anode|cathode|pad|vdd \$136364 i|z$84 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22376 AVDD|anode|cathode|pad|vdd i|z$60 \$136364 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22377 \$133965 i|z|zn$7 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22378 AVDD|anode|cathode|pad|vdd \$133789 \$133966 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22379 \$133789 \$133965 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22380 AVDD|anode|cathode|pad|vdd \$133966 i|z$89 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22381 AVDD|anode|cathode|pad|vdd \$136365 i|z$40 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22383 AVDD|anode|cathode|pad|vdd i|z$105 \$136365 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22384 \$133967 i|z$85 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22385 AVDD|anode|cathode|pad|vdd \$133791 \$133968 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22386 AVDD|anode|cathode|pad|vdd \$136366 i|z$76 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22388 AVDD|anode|cathode|pad|vdd i|z$93 \$136366 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22389 \$133791 \$133967 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22390 AVDD|anode|cathode|pad|vdd \$133968 i|z$93 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22391 AVDD|anode|cathode|pad|vdd \$133970 i|z$49 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22393 AVDD|anode|cathode|pad|vdd i|z$70 \$133970 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22394 \$133971 i|z$82 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22395 AVDD|anode|cathode|pad|vdd \$133792 \$133972 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22396 \$133792 \$133971 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22397 AVDD|anode|cathode|pad|vdd \$133972 i|z$94 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22398 AVDD|anode|cathode|pad|vdd \$135473 \$135390 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22399 \$135472 i|z$20 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22400 AVDD|anode|cathode|pad|vdd \$133974 i|z$85 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22402 AVDD|anode|cathode|pad|vdd i|z$71 \$133974 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22403 \$135473 \$135472 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22404 AVDD|anode|cathode|pad|vdd \$135390 i|z$102 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22405 AVDD|anode|cathode|pad|vdd \$135475 \$135391 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22406 \$135474 i|z$111 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22407 i|z|zn$9 i|zn$13 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=4.164p AD=4.164p PS=17.74u PD=17.74u
M$22415 \$135475 \$135474 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22416 AVDD|anode|cathode|pad|vdd \$135391 i|z$44 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22417 AVDD|anode|cathode|pad|vdd \$136367 i|z$47 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22419 AVDD|anode|cathode|pad|vdd i|z$100 \$136367 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22420 \$133976 i|z$107 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22421 AVDD|anode|cathode|pad|vdd \$133793 \$133977 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22422 AVDD|anode|cathode|pad|vdd \$135477 \$135392 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22423 \$135476 i|zn$13 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22424 \$133793 \$133976 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22425 AVDD|anode|cathode|pad|vdd \$133977 i|z$100 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22426 \$135477 \$135476 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22427 AVDD|anode|cathode|pad|vdd \$135392 i|z$104 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22428 \$133978 i|zn$12 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22429 AVDD|anode|cathode|pad|vdd \$133794 \$133979 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22430 \$133794 \$133978 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22431 AVDD|anode|cathode|pad|vdd \$133979 i|z$95 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22432 AVDD|anode|cathode|pad|vdd \$133982 i|z$51 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22434 AVDD|anode|cathode|pad|vdd i|z$96 \$133982 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22435 AVDD|anode|cathode|pad|vdd \$136368 i|z$78 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22437 AVDD|anode|cathode|pad|vdd i|z$52 \$136368 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22438 AVDD|anode|cathode|pad|vdd \$133983 i|z$72 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22440 AVDD|anode|cathode|pad|vdd i|z$95 \$133983 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22441 \$135478 \$135241 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22442 VDD|pad|pin1|supply|vdd cp|z$2 \$135241 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22443 \$135242 \$135241 \$135431 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22444 \$135431 \$135393 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$22445 \$136579 \$135478 \$135429 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$22446 \$135429 \$135479 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$22447 \$136283 d|zn$6 \$135242 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$22448 VDD|pad|pin1|supply|vdd \$135242 \$135393 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$22449 VDD|pad|pin1|supply|vdd \$135478 \$136283 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$22450 \$135393 \$135241 \$136579 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$22451 VDD|pad|pin1|supply|vdd \$136579 \$135479 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$22452 VDD|pad|pin1|supply|vdd a2|a3|zn \$135183 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22453 \$135183 RST|a1|b|cdn|core|i|p2c b|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$22454 b|zn$4 a1|b|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22455 VDD|pad|pin1|supply|vdd i|z$4 \$133805 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$22456 VDD|pad|pin1|supply|vdd \$133805 cp|i|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$22457 a1|b|i|q$2 \$135479 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22458 \$135394 a2|zn$6 d|zn$2 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22459 d|zn$2 a1|z$13 \$135394 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$22460 \$135394 b|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22461 \$140500 \$140555 \$140500 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$22473 \$137560 \$137560 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22474 \$136908 i|zn$5 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.451625p PS=3.53u PD=2.03u
M$22475 AVDD|anode|cathode|pad|vdd \$136862 \$136909 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=0.85u AS=0.451625p AD=0.48025p PS=2.03u PD=2.83u
M$22476 \$136862 \$136908 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22477 AVDD|anode|cathode|pad|vdd \$136909 i|z$15 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22478 \$136910 i|zn$6 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22484 AVDD|anode|cathode|pad|vdd \$136910 z$7 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22524 \$140501 \$140556 \$140501 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$22560 \$140502 \$140557 \$140502 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$22596 \$136911 i|z$67 AVDD|anode|cathode|pad|vdd AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=6.395u AS=2.774675p AD=2.713175p PS=12.18u PD=12.07u
M$22602 AVDD|anode|cathode|pad|vdd \$136911 z$3 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=19.2u AS=7.968p AD=8.148p PS=32.48u PD=33.98u
M$22618 \$140503 \$140558 \$140503 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$22642 AVDD|anode|cathode|pad|vdd \$136912 i|z$113 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22644 AVDD|anode|cathode|pad|vdd i|z$114 \$136912 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22657 \$140504 \$140559 \$140504 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$22693 \$140505 \$140560 \$140505 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$22717 AVDD|anode|cathode|pad|vdd \$136915 i|z$53 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22719 AVDD|anode|cathode|pad|vdd i|z$112 \$136915 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22732 \$140506 \$140561 \$140506 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$22768 \$140507 \$140562 \$140507 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$22804 AVDD|anode|cathode|pad|vdd \$136916 i|z$111 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=2.4u AS=1.176p AD=0.996p PS=5.56u PD=4.06u
M$22806 AVDD|anode|cathode|pad|vdd i|z$63 \$136916 AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22807 \$140508 \$140563 \$140508 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$22843 \$140509 \$140564 \$140509 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$22879 \$136917 \$136863 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22880 VDD|pad|pin1|supply|vdd cp|i|z \$136863 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22881 VDD|pad|pin1|supply|vdd \$136917 \$138389 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$22882 \$138389 d|zn$9 \$136864 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$22883 \$136864 \$136863 \$138398 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22884 VDD|pad|pin1|supply|vdd \$136918 \$138398 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22885 \$136918 \$136864 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$22886 \$136918 \$136863 \$136865 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$22887 \$136865 \$136917 \$138397 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$22888 VDD|pad|pin1|supply|vdd \$136919 \$138397 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$22889 VDD|pad|pin1|supply|vdd \$136865 \$136919 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$22890 a1|b|i|q$1 \$136919 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$22891 VDD|pad|pin1|supply|vdd a1|z$3 \$140565 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22892 \$140565 a2|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$22893 VDD|pad|pin1|supply|vdd \$140565 d|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22894 \$136920 \$136866 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22895 VDD|pad|pin1|supply|vdd cp|z$3 \$136866 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22896 a2|zn$6 a1|b|i|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$22897 VDD|pad|pin1|supply|vdd a1|a2|a3|z a2|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$22898 a2|zn$6 a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$22899 VDD|pad|pin1|supply|vdd \$136920 \$138399 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$22900 \$138399 d|zn$10 \$136867 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$22901 \$136867 \$136866 \$138412 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22902 VDD|pad|pin1|supply|vdd \$136921 \$138412 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$22903 \$136921 \$136867 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$22904 \$136921 \$136866 \$136868 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$22905 \$136868 \$136920 \$138404 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$22906 VDD|pad|pin1|supply|vdd \$136922 \$138404 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$22907 VDD|pad|pin1|supply|vdd \$136868 \$136922 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$22908 a1|b|i|q \$136922 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$23269 \$142237 \$141920 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23270 VDD|pad|pin1|supply|vdd cp|z$3 \$141920 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23271 \$141921 \$141920 \$142598 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$23272 \$142598 \$142238 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$23273 \$143400 \$142237 \$142588 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$23274 \$142588 \$142239 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$23275 \$142596 d|zn$5 \$141921 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$23276 VDD|pad|pin1|supply|vdd \$141921 \$142238 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$23277 VDD|pad|pin1|supply|vdd \$142237 \$142596 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$23278 \$142238 \$141920 \$143400 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$23279 VDD|pad|pin1|supply|vdd \$143400 \$142239 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$23280 a2|i|q \$142239 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$23281 a2|z \$142241 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23282 VDD|pad|pin1|supply|vdd b|i|q \$142240 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$23283 \$142240 a1|b|i|q \$142241 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$23284 \$142241 a2|zn$5 \$142240 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23285 \$145966 \$146281 \$145966 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23297 \$140555 z$26 \$143729 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23298 \$143729 zn$3 \$143729 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23300 \$140555 zn$3 \$140555 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$23313 \$143730 z$26 \$140555 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23316 \$143730 zn$3 \$143730 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23329 \$143731 z$26 \$140555 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23332 \$143731 zn$3 \$143731 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23333 \$145967 \$146282 \$145967 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=1382.4u AS=590.976p AD=590.976p PS=2482.56u PD=2482.56u
M$23345 \$140556 z$26 \$143732 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23346 \$143732 zn$3 \$143732 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23348 \$140556 zn$3 \$140556 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$23361 \$143733 z$26 \$140556 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23364 \$143733 zn$3 \$143733 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23377 \$143734 z$26 \$140556 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23380 \$143734 zn$3 \$143734 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23381 \$145968 \$146283 \$145968 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=691.2u AS=295.488p AD=295.488p PS=1241.28u PD=1241.28u
M$23393 \$140557 z$26 \$143735 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23394 \$143735 zn$3 \$143735 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23396 \$140557 zn$3 \$140557 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$23409 \$143736 z$26 \$140557 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23412 \$143736 zn$3 \$143736 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23425 \$143737 z$26 \$140557 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23428 \$143737 zn$3 \$143737 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23429 \$145969 \$146284 \$145969 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=172.8u AS=73.872p AD=73.872p PS=310.32u PD=310.32u
M$23441 \$140558 z$26 \$143738 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23442 \$143738 zn$3 \$143738 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23444 \$140558 zn$3 \$140558 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$23457 \$143739 z$26 \$140558 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23460 \$143739 zn$3 \$143739 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23473 \$143740 z$26 \$140558 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23476 \$143740 zn$3 \$143740 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23477 \$145970 \$146285 \$145970 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23489 \$140559 z$26 \$143741 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23490 \$143741 zn$3 \$143741 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23492 \$140559 zn$3 \$140559 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$23505 \$143742 z$26 \$140559 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23508 \$143742 zn$3 \$143742 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23521 \$143743 z$26 \$140559 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23524 \$143743 zn$3 \$143743 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23525 \$145971 \$146286 \$145971 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23537 \$140560 z$26 \$143744 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23538 \$143744 zn$3 \$143744 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23540 \$140560 zn$3 \$140560 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$23553 \$143745 z$26 \$140560 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23556 \$143745 zn$3 \$143745 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23569 \$143746 z$26 \$140560 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23572 \$143746 zn$3 \$143746 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23585 \$140561 z$26 \$143747 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23586 \$143747 zn$3 \$143747 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23588 \$140561 zn$3 \$140561 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$23601 \$143748 z$26 \$140561 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23604 \$143748 zn$3 \$143748 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23617 \$143749 z$26 \$140561 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23620 \$143749 zn$3 \$143749 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23633 \$140562 z$26 \$143750 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23634 \$143750 zn$3 \$143750 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23636 \$140562 zn$3 \$140562 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$23649 \$143751 z$26 \$140562 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23652 \$143751 zn$3 \$143751 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23665 \$143752 z$26 \$140562 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23668 \$143752 zn$3 \$143752 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23681 \$140563 z$26 \$143753 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23682 \$143753 zn$3 \$143753 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23684 \$140563 zn$3 \$140563 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$23697 \$143754 z$26 \$140563 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23700 \$143754 zn$3 \$143754 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23713 \$143755 z$26 \$140563 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23716 \$143755 zn$3 \$143755 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23717 \$145972 \$146287 \$145972 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$23729 \$140564 z$26 \$143756 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23730 \$143756 zn$3 \$143756 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23732 \$140564 zn$3 \$140564 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$23745 \$143757 z$26 \$140564 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23748 \$143757 zn$3 \$143757 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23761 \$143758 z$26 \$140564 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$23764 \$143758 zn$3 \$143758 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$23765 \$145714 \$144911 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23766 VDD|pad|pin1|supply|vdd cp|z$3 \$144911 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23767 \$144913 \$144911 \$145557 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$23768 \$145557 \$144914 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.251625p PS=1.13u PD=1.58u
M$23769 \$146288 \$145714 \$145573 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$23770 \$145573 \$146170 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.1245p AD=0.37875p PS=1.13u PD=2.03u
M$23771 \$145963 d|z$4 \$144913 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$23772 VDD|pad|pin1|supply|vdd \$144913 \$144914 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.251625p AD=0.4002375p PS=1.58u PD=1.895u
M$23773 VDD|pad|pin1|supply|vdd \$145714 \$145963 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$23774 \$144914 \$144911 \$146288 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$23775 VDD|pad|pin1|supply|vdd \$146288 \$146170 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$23776 VDD|pad|pin1|supply|vdd a2|a3|zn \$144829 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$23777 \$144829 RST|a1|b|cdn|core|i|p2c b|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$23778 b|zn$5 a1|b|i|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$23779 b|i|q$2 \$146170 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$24140 \$151000 \$151285 \$151000 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$24152 \$146281 z$26 \$149147 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24153 \$149147 zn$3 \$149147 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24155 \$146281 zn$3 \$146281 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24168 \$149148 z$26 \$146281 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24171 \$149148 zn$3 \$149148 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24184 \$149149 z$26 \$146281 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24187 \$149149 zn$3 \$149149 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24200 \$146282 z$4 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=19.2u AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$24201 a2$1 z$1 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u
+ AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$24203 \$146282 z$1 \$146282 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$24216 VIN|core|padres z$7 \$146282 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=19.2u AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$24217 \$146282 z$3 \$146282 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$24219 VIN|core|padres z$3 VIN|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$24232 VIP|core|padres z$27 \$146282 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=19.2u AS=10.848p AD=10.848p PS=74.56u PD=74.56u
M$24233 \$146282 zn$5 \$146282 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$24235 VIP|core|padres zn$5 VIP|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$24248 \$146283 z$7 VREFL|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$24249 VREFL|core|padres z$3 VREFL|core|padres AVDD|anode|cathode|pad|vdd
+ sg13_lv_pmos L=0.13u W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$24251 \$146283 z$3 \$146283 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$24264 a2$1 z$9 \$146283 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=9.6u AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$24265 \$146283 z \$146283 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$24267 a2$1 z a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$24280 a2 z$8 \$146283 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=9.6u
+ AS=5.424p AD=5.424p PS=37.28u PD=37.28u
M$24281 \$146283 z$5 \$146283 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$24283 a2 z$5 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$24284 \$151001 \$151286 \$151001 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=345.6u AS=147.744p AD=147.744p PS=620.64u PD=620.64u
M$24296 \$146284 z$7 VREFL|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$24299 \$146284 z$3 \$146284 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24312 a2$1 z$14 \$146284 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$24313 \$146284 z$15 \$146284 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24315 a2$1 z$15 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24328 a2 z$16 \$146284 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$24329 \$146284 z$19 \$146284 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24331 a2 z$19 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24344 \$146285 z$7 VREFL|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24347 \$146285 z$3 \$146285 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24360 a2$1 z$17 \$146285 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24361 \$146285 z$25 \$146285 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24363 a2$1 z$25 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24376 a2 z$21 \$146285 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24377 \$146285 z$23 \$146285 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24379 a2 z$23 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24392 \$146286 z$7 VREFL|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24395 \$146286 z$3 \$146286 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24408 a2$1 z$24 \$146286 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24409 \$146286 zn$4 \$146286 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24411 a2$1 zn$4 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24424 a2 z$24 \$146286 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=1.2u
+ AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24427 a2 zn$4 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=0.6u
+ AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24572 \$151002 \$151287 \$151002 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$24584 \$146287 z$26 \$149150 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24585 \$149150 zn$3 \$149150 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24587 \$146287 zn$3 \$146287 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$24600 \$149151 z$26 \$146287 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24603 \$149151 zn$3 \$149151 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24616 \$149152 z$26 \$146287 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$24619 \$149152 zn$3 \$149152 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$24620 a1|z$3 \$146994 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$24621 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$147684
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p
+ PS=2.03u PD=2.03u
M$24622 \$147684 a1|i|q \$146994 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$24623 \$146994 a2|z$2 \$147684 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$24624 a2|z$6 \$150022 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$24625 VDD|pad|pin1|supply|vdd b|i|q$1 \$150823 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$24626 \$150823 a1|i|q$1 \$150022 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$24627 \$150022 a2|zn$5 \$150823 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$24628 VDD|pad|pin1|supply|vdd a2|zn$3 \$148996 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$24629 \$148996 a1|z$9 d|zn$9 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$24630 d|zn$9 b|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$24631 VDD|pad|pin1|supply|vdd a1|z$3 \$151288 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$24632 \$151288 a2|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$24633 VDD|pad|pin1|supply|vdd \$151288 d|z$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$24634 VDD|pad|pin1|supply|vdd a1|z$3 \$146995 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$24635 \$146995 a2|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$24636 VDD|pad|pin1|supply|vdd \$146995 d|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$24637 VDD|pad|pin1|supply|vdd cp|i|z \$146996 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.6u AS=0.4185p AD=0.339p PS=2.03u PD=2.33u
M$24638 VDD|pad|pin1|supply|vdd \$146996 cp|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.4185p AD=0.678p PS=2.03u PD=3.53u
M$24999 \$155911 \$156793 \$155911 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$25011 \$151285 z$26 \$154109 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25012 \$154109 zn$3 \$154109 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25014 \$151285 zn$3 \$151285 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$25027 \$154110 z$26 \$151285 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25030 \$154110 zn$3 \$154110 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25043 \$154111 z$26 \$151285 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25046 \$154111 zn$3 \$154111 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25155 \$151286 z$7 VREFL|core|padres AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$25158 \$151286 z$3 \$151286 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$25171 a2$1 z$12 \$151286 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=4.8u AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$25172 \$151286 z$11 \$151286 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$25174 a2$1 z$11 a2$1 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$25187 a2 z$10 \$151286 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=4.8u
+ AS=2.712p AD=2.712p PS=18.64u PD=18.64u
M$25188 \$151286 z$13 \$151286 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=2.4u AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$25190 a2 z$13 a2 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u W=2.4u
+ AS=1.356p AD=1.356p PS=9.32u PD=9.32u
M$25431 \$155912 \$156794 \$155912 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$25443 \$151287 z$26 \$154112 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25444 \$154112 zn$3 \$154112 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25446 \$151287 zn$3 \$151287 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$25459 \$154113 z$26 \$151287 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25462 \$154113 zn$3 \$154113 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25475 \$154114 z$26 \$151287 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25478 \$154114 zn$3 \$154114 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25479 a1|z$13 RESULT[0]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$25480 a2|z$7 \$155837 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$25481 VDD|pad|pin1|supply|vdd b|i|q$3 \$156836 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25482 \$156836 a1|b|i|q$3 \$155837 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25483 \$155837 a2|zn$5 \$156836 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$25484 VDD|pad|pin1|supply|vdd a2|a3|zn \$153820 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$25485 \$153820 RST|a1|b|cdn|core|i|p2c b|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25486 b|zn$6 a1|b|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$25487 VDD|pad|pin1|supply|vdd a2|zn$3 \$154645 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$25488 \$154645 a1|z$1 d|zn$10 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25489 d|zn$10 b|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$25490 a1|z RESULT[4]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$25491 VDD|pad|pin1|supply|vdd VALID|a3|c2p|core|i|z \$155838
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$25492 VDD|pad|pin1|supply|vdd \$155838 RD[8]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$25493 VDD|pad|pin1|supply|vdd SAMPLE|a1|c2p|core|i|z \$155840
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$25494 VDD|pad|pin1|supply|vdd \$155840 RD[9]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$25855 a2|zn$1 a1|b|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$25856 VDD|pad|pin1|supply|vdd a1|a2|a3|z a2|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$25857 a2|zn$1 a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$25858 \$161605 \$162307 \$161605 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$25870 \$156793 z$26 \$159940 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25871 \$159940 zn$3 \$159940 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25873 \$156793 zn$3 \$156793 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$25886 \$159941 z$26 \$156793 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25889 \$159941 zn$3 \$159941 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$25902 \$159942 z$26 \$156793 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$25905 \$159942 zn$3 \$159942 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26290 \$161606 \$162308 \$161606 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$26302 \$156794 z$26 \$159943 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26303 \$159943 zn$3 \$159943 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26305 \$156794 zn$3 \$156794 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$26318 \$159944 z$26 \$156794 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26321 \$159944 zn$3 \$159944 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26334 \$159945 z$26 \$156794 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26337 \$159945 zn$3 \$159945 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26338 \$159264 \$158745 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$26339 VDD|pad|pin1|supply|vdd cp|z$3 \$158745 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$26340 VDD|pad|pin1|supply|vdd \$159264 \$160281 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.885u AS=0.500025p AD=0.3493875p PS=2.9u PD=1.715u
M$26341 \$160281 a2|d|zn \$158746 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.75u AS=0.3493875p AD=0.251625p PS=1.715u PD=1.58u
M$26342 \$158746 \$158745 \$160283 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$26343 VDD|pad|pin1|supply|vdd \$158998 \$160283 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.251625p AD=0.1245p PS=1.58u PD=1.13u
M$26344 \$158998 \$158746 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.75u AS=0.4002375p AD=0.251625p PS=1.895u PD=1.58u
M$26345 \$158998 \$158745 \$158747 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.065u AS=0.4002375p AD=0.3406125p PS=1.895u PD=1.895u
M$26346 \$158747 \$159264 \$160278 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.3u AS=0.3406125p AD=0.1245p PS=1.895u PD=1.13u
M$26347 VDD|pad|pin1|supply|vdd \$159265 \$160278 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.3u AS=0.37875p AD=0.1245p PS=2.03u PD=1.13u
M$26348 VDD|pad|pin1|supply|vdd \$158747 \$159265 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.37875p AD=0.678p PS=2.03u PD=3.53u
M$26349 a2|zn$2 a1|b|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$26350 VDD|pad|pin1|supply|vdd a1|a2|a3|z a2|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$26351 a2|zn$2 a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$26352 a1|i|q \$159265 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$26713 \$163468 a2|zn$4 d|zn$7 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$26714 d|zn$7 a1|z$8 \$163468 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$26715 \$163468 b|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$26716 VDD|pad|pin1|supply|vdd a2|a3|zn \$163558 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$26717 \$163558 RST|a1|b|cdn|core|i|p2c a2|d|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$26718 \$167430 \$168095 \$167430 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$26730 \$162307 z$26 \$165672 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26731 \$165672 zn$3 \$165672 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26733 \$162307 zn$3 \$162307 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$26746 \$165673 z$26 \$162307 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26749 \$165673 zn$3 \$165673 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26762 \$165674 z$26 \$162307 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$26765 \$165674 zn$3 \$165674 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$26766 \$167431 \$168096 \$167431 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$26814 \$167432 \$168097 \$167432 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$26862 \$167433 \$168098 \$167433 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$26910 \$167434 \$168099 \$167434 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$26958 \$167435 \$168100 \$167435 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27006 \$167436 \$168101 \$167436 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27054 \$167437 \$168102 \$167437 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27102 \$167438 \$168103 \$167438 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27150 \$167439 \$168104 \$167439 AVDD|anode|cathode|pad|vdd sg13_lv_pmos
+ L=0.13u W=86.4u AS=36.936p AD=36.936p PS=155.16u PD=155.16u
M$27162 \$162308 z$26 \$165675 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27163 \$165675 zn$3 \$165675 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27165 \$162308 zn$3 \$162308 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27178 \$165676 z$26 \$162308 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27181 \$165676 zn$3 \$165676 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27194 \$165677 z$26 \$162308 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27197 \$165677 zn$3 \$165677 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27198 VDD|pad|pin1|supply|vdd a2|zn$3 \$164354 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$27199 \$164354 a1|z$2 d|zn$8 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$27200 d|zn$8 b|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$27201 VDD|pad|pin1|supply|vdd a2|a3|zn \$166704 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$27202 \$166704 RST|a1|b|cdn|core|i|p2c b|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$27203 b|zn$3 a1|b|i|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$27204 a2|zn$3 a1|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$27205 VDD|pad|pin1|supply|vdd a2|z$2 a2|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.498p PS=2.03u PD=2.03u
M$27206 a2|zn$3 a1|a2|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$27207 a1|z$7 a1|i|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$27568 \$168095 z$26 \$170779 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27569 \$170779 zn$3 \$170779 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27571 \$168095 zn$3 \$168095 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27572 \$170780 z$26 \$168095 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27575 \$170780 zn$3 \$170780 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27576 \$170781 z$26 \$168095 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27579 \$170781 zn$3 \$170781 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27580 \$168096 z$26 \$170782 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27581 \$170782 zn$3 \$170782 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27583 \$168096 zn$3 \$168096 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27584 \$170783 z$26 \$168096 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27587 \$170783 zn$3 \$170783 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27588 \$170784 z$26 \$168096 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27591 \$170784 zn$3 \$170784 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27592 \$168097 z$26 \$170785 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27593 \$170785 zn$3 \$170785 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27595 \$168097 zn$3 \$168097 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27596 \$170786 z$26 \$168097 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27599 \$170786 zn$3 \$170786 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27600 \$170787 z$26 \$168097 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27603 \$170787 zn$3 \$170787 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27604 \$168098 z$26 \$170788 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27605 \$170788 zn$3 \$170788 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27607 \$168098 zn$3 \$168098 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27608 \$170789 z$26 \$168098 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27611 \$170789 zn$3 \$170789 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27612 \$170790 z$26 \$168098 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27615 \$170790 zn$3 \$170790 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27616 \$168099 z$26 \$170791 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27617 \$170791 zn$3 \$170791 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27619 \$168099 zn$3 \$168099 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27620 \$170792 z$26 \$168099 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27623 \$170792 zn$3 \$170792 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27624 \$170793 z$26 \$168099 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27627 \$170793 zn$3 \$170793 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27628 \$168100 z$26 \$170794 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27629 \$170794 zn$3 \$170794 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27631 \$168100 zn$3 \$168100 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27632 \$170795 z$26 \$168100 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27635 \$170795 zn$3 \$170795 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27636 \$170796 z$26 \$168100 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27639 \$170796 zn$3 \$170796 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27640 \$168101 z$26 \$170797 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27641 \$170797 zn$3 \$170797 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27643 \$168101 zn$3 \$168101 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27644 \$170798 z$26 \$168101 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27647 \$170798 zn$3 \$170798 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27648 \$170799 z$26 \$168101 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27651 \$170799 zn$3 \$170799 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27652 \$168102 z$26 \$170800 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27653 \$170800 zn$3 \$170800 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27655 \$168102 zn$3 \$168102 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27656 \$170801 z$26 \$168102 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27659 \$170801 zn$3 \$170801 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27660 \$170802 z$26 \$168102 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27663 \$170802 zn$3 \$170802 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27664 \$168103 z$26 \$170803 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27665 \$170803 zn$3 \$170803 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27667 \$168103 zn$3 \$168103 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27668 \$170804 z$26 \$168103 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27671 \$170804 zn$3 \$170804 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27672 \$170805 z$26 \$168103 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27675 \$170805 zn$3 \$170805 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27676 \$168104 z$26 \$170806 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27677 \$170806 zn$3 \$170806 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27679 \$168104 zn$3 \$168104 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.8u AS=1.017p AD=1.017p PS=6.99u PD=6.99u
M$27680 \$170807 z$26 \$168104 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27683 \$170807 zn$3 \$170807 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27684 \$170808 z$26 \$168104 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=1.2u AS=0.678p AD=0.678p PS=4.66u PD=4.66u
M$27687 \$170808 zn$3 \$170808 AVDD|anode|cathode|pad|vdd sg13_lv_pmos L=0.13u
+ W=0.6u AS=0.339p AD=0.339p PS=2.33u PD=2.33u
M$27688 \$230018 \$229344 \$230017 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$27689 \$230018 R[48]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$27690 VDD|pad|pin1|supply|vdd i0|i1|q \$230019 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$27691 \$230019 s|zn \$230017 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$27692 a1|z$9 a1|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$27693 \$230022 \$229345 \$230021 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$27694 \$230022 R[56]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$27695 VDD|pad|pin1|supply|vdd i0|i1|q \$230023 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$27696 \$230023 s|zn$1 \$230021 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$27697 a1|z$10 a1|b|i|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p PS=3.53u PD=3.53u
M$27698 VDD|pad|pin1|supply|vdd \$213964 \$213964 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27699 VDD|pad|pin1|supply|vdd a2|a3|z \$170727 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.498p PS=3.53u PD=2.03u
M$27700 \$170727 RST|a1|b|cdn|core|i|p2c a2|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.2u AS=0.498p AD=0.678p PS=2.03u PD=3.53u
M$27701 a1|z$4 RESULT[3]|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.2u AS=0.678p AD=0.678p
+ PS=3.53u PD=3.53u
M$27702 \$230027 \$229346 \$230026 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$27703 \$230027 R[51]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$27704 VDD|pad|pin1|supply|vdd i0|i1|q$1 \$230028 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$27705 \$230028 s|zn \$230026 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$27706 VDD|pad|pin1|supply|vdd \$213965 \$213965 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27707 VDD|pad|pin1|supply|vdd R[13]|i|i0|q \$213461 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27708 VDD|pad|pin1|supply|vdd \$213461 RD[45]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27709 VDD|pad|pin1|supply|vdd R[15]|i|i0|q \$213462 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27710 VDD|pad|pin1|supply|vdd \$213462 RD[47]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27711 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a4|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27712 a4|zn$1 a2|z$9 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$27713 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a4|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27714 VDD|pad|pin1|supply|vdd i$2 \$213463 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27715 VDD|pad|pin1|supply|vdd \$213463 RD[3]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27716 a4|zn$1 RD[45]|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27717 VDD|pad|pin1|supply|vdd R[6]|i|i0|q \$213464 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27718 VDD|pad|pin1|supply|vdd \$213464 RD[38]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27719 VDD|pad|pin1|supply|vdd \$213970 \$213970 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27720 VDD|pad|pin1|supply|vdd \$215219 RD[30]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27721 VDD|pad|pin1|supply|vdd RD[38]|a2|z a1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27722 a1|zn$1 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$27723 VDD|pad|pin1|supply|vdd \$215220 RD[21]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27724 a1|zn$1 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27725 VDD|pad|pin1|supply|vdd R[12]|i|i0|q \$213466 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27726 VDD|pad|pin1|supply|vdd \$213466 RD[44]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27727 VDD|pad|pin1|supply|vdd RD[1]|a2|z a2|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27728 a2|zn$7 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$27729 VDD|pad|pin1|supply|vdd \$215221 RD[24]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27730 a2|zn$7 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27731 VDD|pad|pin1|supply|vdd \$215222 RD[23]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27732 VDD|pad|pin1|supply|vdd a3|zn a2|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27733 a2|zn$12 a2|zn$13 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$27734 VDD|pad|pin1|supply|vdd a1|zn$4 a2|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27735 VDD|pad|pin1|supply|vdd \$212052 \$212052 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27736 VDD|pad|pin1|supply|vdd R[14]|i|i0|q \$213468 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27737 VDD|pad|pin1|supply|vdd \$213468 RD[46]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27738 RD[1]|a2|z \$211248 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$27739 VDD|pad|pin1|supply|vdd i \$211248 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27740 a2|zn$12 a4|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27741 VDD|pad|pin1|supply|vdd \$213974 \$213974 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27742 VDD|pad|pin1|supply|vdd a2|zn$11 a1|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$27743 a1|zn$2 a1|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$27744 VDD|pad|pin1|supply|vdd R[2]|i|i0|q \$213469 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27745 VDD|pad|pin1|supply|vdd \$213469 RD[34]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27746 VDD|pad|pin1|supply|vdd \$212053 \$212053 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27747 VDD|pad|pin1|supply|vdd a2|zn$7 \$230032 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27748 \$230032 a1|zn$10 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$27749 RD[17]|a4|z \$215224 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27750 VDD|pad|pin1|supply|vdd R[8]|i|i0|q \$213470 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27751 VDD|pad|pin1|supply|vdd \$213470 RD[40]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27752 a1|z$14 \$230032 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27753 \$213978 \$213978 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27754 VDD|pad|pin1|supply|vdd RD[37]|a2|z a3|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27755 a3|zn a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$27756 RD[0]|a2|z \$211251 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$27757 VDD|pad|pin1|supply|vdd i$1 \$211251 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27758 \$213979 \$213979 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27759 a3|zn a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27760 VDD|pad|pin1|supply|vdd R[10]|i|i0|q \$213471 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27761 VDD|pad|pin1|supply|vdd \$213471 RD[42]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27762 RD[19]|a4|z \$211252 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27763 VDD|pad|pin1|supply|vdd RD[26]|a2|z a1|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27764 a1|zn$3 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$27765 RD[26]|a2|z \$211253 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27766 a1|zn$3 a2|a3|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27767 VDD|pad|pin1|supply|vdd R[5]|i|i0|q \$213472 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27768 VDD|pad|pin1|supply|vdd \$213472 RD[37]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27769 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27770 a2|zn$8 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$27771 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27772 VDD|pad|pin1|supply|vdd R[9]|i|i0|q \$213473 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27773 VDD|pad|pin1|supply|vdd \$213473 RD[41]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27774 a2|zn$8 RD[18]|a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27775 VDD|pad|pin1|supply|vdd R[3]|i|i0|q \$213474 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27776 VDD|pad|pin1|supply|vdd \$213474 RD[35]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27777 VDD|pad|pin1|supply|vdd a2|zn$20 a1|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$27778 a1|zn$8 a1|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$27779 VDD|pad|pin1|supply|vdd R[4]|i|i0|q \$213475 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27780 VDD|pad|pin1|supply|vdd \$213475 RD[36]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27781 VDD|pad|pin1|supply|vdd a2|zn$9 \$230037 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27782 \$230037 a1|zn$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$27783 VDD|pad|pin1|supply|vdd R[11]|i|i0|q \$213476 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27784 VDD|pad|pin1|supply|vdd \$213476 RD[43]|a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27785 a2|z$8 \$230037 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27786 \$213984 \$213984 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27787 VDD|pad|pin1|supply|vdd RD[34]|a2|z a1|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27788 a1|zn$6 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$27789 VDD|pad|pin1|supply|vdd \$213985 \$213985 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27790 VDD|pad|pin1|supply|vdd R[1]|i|i0|q \$213477 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27791 VDD|pad|pin1|supply|vdd \$213477 RD[33]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27792 a1|zn$6 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27793 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a4|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27794 a4|zn a2|z$9 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$27795 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a4|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27796 VDD|pad|pin1|supply|vdd \$213987 \$213987 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27797 VDD|pad|pin1|supply|vdd \$213988 \$213988 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27798 a4|zn RD[43]|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27799 \$213989 \$213989 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27800 VDD|pad|pin1|supply|vdd RD[28]|a2|z a2|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27801 a2|zn$10 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$27802 VDD|pad|pin1|supply|vdd i$3 \$213478 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27803 VDD|pad|pin1|supply|vdd \$213478 RD[2]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27804 a2|zn$10 a2|a3|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27805 VDD|pad|pin1|supply|vdd R[0]|i|i0|q \$213479 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27806 VDD|pad|pin1|supply|vdd \$213479 RD[32]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27807 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27808 a1|zn a2|z$9 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$27809 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a1|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27810 RD[28]|a2|z \$215232 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27811 VDD|pad|pin1|supply|vdd i$4 \$213480 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27812 VDD|pad|pin1|supply|vdd \$213480 RD[4]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27813 a1|zn RD[15]|a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27814 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27815 a2|zn$9 a2|z$9 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$27816 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27817 \$213993 \$213993 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27818 a2|zn$9 RD[9]|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$27819 VDD|pad|pin1|supply|vdd R[7]|i|i0|q \$213481 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$27820 VDD|pad|pin1|supply|vdd \$213481 RD[39]|a2|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$27821 \$230042 \$229361 \$230041 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$27822 \$230042 R[59]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$27823 VDD|pad|pin1|supply|vdd i0|i1|q$1 \$230043 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$27824 \$230043 s|zn$1 \$230041 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$27825 \$213995 \$213995 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27826 \$213996 \$213996 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27827 \$213997 \$213997 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$27828 \$200626 DOUT_DAT|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$27829 DATA|core|i0|i1|p2c \$231093 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$27830 \$202259 DOUT_DAT|c2p|core|i|q VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$27831 \$230012 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$27832 VDD|pad|pin1|supply|vdd \$230012 \$229341 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$27833 VDD|pad|pin1|supply|vdd \$229341 \$231312 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$27834 \$231312 d|z$8 \$230013 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$27835 \$230013 \$230012 \$231088 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$27836 \$231088 \$230014 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$27837 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$231088
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$27838 \$230014 \$230013 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$27839 \$230014 \$230012 \$229342 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$27840 \$229342 \$229341 \$231320 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$27841 VDD|pad|pin1|supply|vdd \$230016 \$231320 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$27842 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230016
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$27843 VDD|pad|pin1|supply|vdd \$229342 \$230016 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$27844 VDD|pad|pin1|supply|vdd \$230016 R[51]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$27845 VDD|pad|pin1|supply|vdd s|zn \$229344 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$27846 VDD|pad|pin1|supply|vdd \$230017 d|z$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$27847 VDD|pad|pin1|supply|vdd s|zn$1 \$229345 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$27848 VDD|pad|pin1|supply|vdd \$230021 d|z$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$27849 VDD|pad|pin1|supply|vdd s|zn \$229346 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$27850 VDD|pad|pin1|supply|vdd \$230026 d|z$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$27851 VDD|pad|pin1|supply|vdd s|zn$1 \$229361 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$27852 VDD|pad|pin1|supply|vdd \$230041 d|z$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$27853 \$230045 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$27854 VDD|pad|pin1|supply|vdd \$230045 \$229362 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$27855 VDD|pad|pin1|supply|vdd \$229362 \$231291 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$27856 \$231291 d|z$7 \$230046 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$27857 \$230046 \$230045 \$231092 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$27858 \$231092 \$230047 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$27859 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$231092
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$27860 \$230047 \$230046 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$27861 \$230047 \$230045 \$229363 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$27862 \$229363 \$229362 \$231283 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$27863 VDD|pad|pin1|supply|vdd \$230049 \$231283 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$27864 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$230049
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$27865 VDD|pad|pin1|supply|vdd \$229363 \$230049 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$27866 VDD|pad|pin1|supply|vdd \$230049 R[59]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$27867 \$231703 \$231480 \$231704 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$27868 \$231705 s|zn$2 \$231703 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$27869 VDD|pad|pin1|supply|vdd i0|i1|q$1 \$231705 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$27870 \$231704 R[35]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$27871 \$231480 s|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$27872 VDD|pad|pin1|supply|vdd \$231703 d|z$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$27873 VDD|pad|pin1|supply|vdd cp|z$4 \$231707 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$27874 VDD|pad|pin1|supply|vdd \$231707 \$231708 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$27875 VDD|pad|pin1|supply|vdd \$232243 \$231710 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$27876 \$231709 \$231707 \$231710 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$27877 VDD|pad|pin1|supply|vdd \$231708 \$232241 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$27878 \$232241 d|z$5 \$231709 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$27879 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$231710
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$27880 \$231711 \$231708 \$231745 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$27881 VDD|pad|pin1|supply|vdd \$232244 \$231745 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$27882 VDD|pad|pin1|supply|vdd \$231709 \$232243 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$27883 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232244
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$27884 VDD|pad|pin1|supply|vdd \$231711 \$232244 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$27885 \$232243 \$231707 \$231711 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$27886 VDD|pad|pin1|supply|vdd \$232244 R[48]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$27887 VDD|pad|pin1|supply|vdd cp|z$4 \$231712 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$27888 VDD|pad|pin1|supply|vdd \$231712 \$231713 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$27889 VDD|pad|pin1|supply|vdd \$232245 \$231715 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$27890 \$231714 \$231712 \$231715 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$27891 VDD|pad|pin1|supply|vdd \$231713 \$232242 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$27892 \$232242 d|z$6 \$231714 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$27893 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$231715
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$27894 \$231716 \$231713 \$231744 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$27895 VDD|pad|pin1|supply|vdd \$232246 \$231744 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$27896 VDD|pad|pin1|supply|vdd \$231714 \$232245 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$27897 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232246
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$27898 VDD|pad|pin1|supply|vdd \$231716 \$232246 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$27899 \$232245 \$231712 \$231716 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$27900 VDD|pad|pin1|supply|vdd \$232246 R[56]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$27901 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a4|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27902 VDD|pad|pin1|supply|vdd a2|z$9 a4|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27903 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a4|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27904 VDD|pad|pin1|supply|vdd RD[42]|a4|z a4|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27905 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a3|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27906 VDD|pad|pin1|supply|vdd a2|z$9 a3|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27907 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a3|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27908 VDD|pad|pin1|supply|vdd RD[41]|a4|z a3|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27909 VDD|pad|pin1|supply|vdd a3|zn$3 i1|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27910 VDD|pad|pin1|supply|vdd a2|z$10 i1|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27911 VDD|pad|pin1|supply|vdd a1|zn$9 i1|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27912 VDD|pad|pin1|supply|vdd a4|z i1|zn VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27913 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27914 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a2|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27915 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27916 VDD|pad|pin1|supply|vdd RD[21]|a4|z a2|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27917 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27918 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a1|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27919 VDD|pad|pin1|supply|vdd a1|z$15 a1|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27920 VDD|pad|pin1|supply|vdd RD[17]|a4|z a1|zn$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27921 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27922 VDD|pad|pin1|supply|vdd a2|z$9 a1|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27923 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a1|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27924 VDD|pad|pin1|supply|vdd RD[13]|a4|zn a1|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27925 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27926 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a2|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27927 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27928 VDD|pad|pin1|supply|vdd RD[19]|a4|z a2|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27929 VDD|pad|pin1|supply|vdd a3|zn$5 a2|zn$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27930 VDD|pad|pin1|supply|vdd a2|zn$14 a2|zn$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27931 VDD|pad|pin1|supply|vdd a1|zn$14 a2|zn$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27932 VDD|pad|pin1|supply|vdd a4|zn a2|zn$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27933 VDD|pad|pin1|supply|vdd a3|zn$7 a2|zn$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27934 VDD|pad|pin1|supply|vdd a2|zn$8 a2|zn$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27935 VDD|pad|pin1|supply|vdd a1|zn$3 a2|zn$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27936 VDD|pad|pin1|supply|vdd a4|zn$2 a2|zn$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27937 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a4|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27938 VDD|pad|pin1|supply|vdd a2|z$9 a4|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27939 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a4|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27940 VDD|pad|pin1|supply|vdd RD[44]|a4|z a4|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27941 VDD|pad|pin1|supply|vdd a3|zn$2 i1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27942 VDD|pad|pin1|supply|vdd a2|z$8 i1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27943 VDD|pad|pin1|supply|vdd a1|z$14 i1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27944 VDD|pad|pin1|supply|vdd a4|zn$4 i1|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27945 VDD|pad|pin1|supply|vdd RD[25]|a2|zn a4|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27946 VDD|pad|pin1|supply|vdd a1|a3|z a4|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27947 VDD|pad|pin1|supply|vdd a2|a3|z$1 a4|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27948 VDD|pad|pin1|supply|vdd a3|zn$1 a2|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27949 VDD|pad|pin1|supply|vdd a2|zn$10 a2|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27950 VDD|pad|pin1|supply|vdd a1|zn$13 a2|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27951 VDD|pad|pin1|supply|vdd a4|zn$3 a2|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27952 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27953 VDD|pad|pin1|supply|vdd a2|z$9 a1|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27954 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a1|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27955 VDD|pad|pin1|supply|vdd RD[11]|a4|zn a1|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27956 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27957 VDD|pad|pin1|supply|vdd a2|z$9 a1|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$27958 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a1|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$27959 VDD|pad|pin1|supply|vdd RD[8]|a4|z a1|zn$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27960 VDD|pad|pin1|supply|vdd RD[4]|a2|z a1|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27961 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$27962 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a1|zn$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$27963 \$231732 \$231484 \$231733 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$27964 \$231734 s|zn$1 \$231732 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$27965 VDD|pad|pin1|supply|vdd i0|i1|q$2 \$231734 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$27966 \$231733 R[58]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$27967 \$231484 s|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$27968 VDD|pad|pin1|supply|vdd \$231732 d|z$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$27969 VDD|pad|pin1|supply|vdd cp|i|z$1 \$231736 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$27970 VDD|pad|pin1|supply|vdd \$231736 \$231737 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$27971 VDD|pad|pin1|supply|vdd \$232249 \$231739 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$27972 \$231738 \$231736 \$231739 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$27973 VDD|pad|pin1|supply|vdd \$231737 \$232165 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$27974 \$232165 d|z$11 \$231738 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$27975 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$231739
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$27976 \$231740 \$231737 \$231743 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$27977 VDD|pad|pin1|supply|vdd \$232250 \$231743 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$27978 VDD|pad|pin1|supply|vdd \$231738 \$232249 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$27979 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$232250
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$27980 VDD|pad|pin1|supply|vdd \$231740 \$232250 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$27981 \$232249 \$231736 \$231740 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$27982 VDD|pad|pin1|supply|vdd \$232250 R[50]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$27983 \$233645 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$27984 VDD|pad|pin1|supply|vdd \$233645 \$233646 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$27985 VDD|pad|pin1|supply|vdd \$233646 \$235389 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$27986 \$235389 d|z$16 \$233647 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$27987 \$233647 \$233645 \$235337 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$27988 \$235337 \$233648 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$27989 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$235337
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$27990 \$233648 \$233647 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$27991 \$233648 \$233645 \$233649 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$27992 \$233649 \$233646 \$235390 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$27993 VDD|pad|pin1|supply|vdd \$233651 \$235390 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$27994 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$233651
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$27995 VDD|pad|pin1|supply|vdd \$233649 \$233651 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$27996 VDD|pad|pin1|supply|vdd \$233651 R[53]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$27997 \$233653 \$233655 \$233652 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$27998 \$233653 R[60]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$27999 VDD|pad|pin1|supply|vdd i0|i1|q$3 \$233654 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28000 \$233654 s|zn$1 \$233652 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28001 VDD|pad|pin1|supply|vdd s|zn$1 \$233655 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28002 VDD|pad|pin1|supply|vdd \$233652 d|z$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28003 \$233658 \$233660 \$233657 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28004 \$233658 R[55]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28005 VDD|pad|pin1|supply|vdd i0|i1|q$4 \$233659 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28006 \$233659 s|zn \$233657 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28007 VDD|pad|pin1|supply|vdd s|zn \$233660 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28008 VDD|pad|pin1|supply|vdd \$233657 d|z$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28009 \$233663 \$233665 \$233662 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28010 \$233663 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28011 VDD|pad|pin1|supply|vdd R[2]|i|i0|q \$233664 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28012 \$233664 s|z \$233662 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28013 VDD|pad|pin1|supply|vdd s|z \$233665 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28014 VDD|pad|pin1|supply|vdd \$233662 d|z$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28015 \$233668 \$233670 \$233667 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28016 \$233668 R[53]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28017 VDD|pad|pin1|supply|vdd i0|i1|q$5 \$233669 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28018 \$233669 s|zn \$233667 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28019 VDD|pad|pin1|supply|vdd s|zn \$233670 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28020 VDD|pad|pin1|supply|vdd \$233667 d|z$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28021 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a2|zn$18 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28022 a2|zn$18 a2|z$9 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$28023 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$18 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28024 a2|zn$18 RD[47]|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28025 VDD|pad|pin1|supply|vdd RD[30]|a2|z a3|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28026 a3|zn$4 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28027 a3|zn$4 a2|a3|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28028 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28029 a1|zn$15 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$28030 VDD|pad|pin1|supply|vdd a1|z$15 a1|zn$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28031 a1|zn$15 RD[23]|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28032 VDD|pad|pin1|supply|vdd RD[6]|a2|zn a1|zn$16 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28033 a1|zn$16 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28034 a1|zn$16 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28035 \$233679 a1|zn$2 \$235396 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$28036 \$235396 a2|zn$12 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$28037 VDD|pad|pin1|supply|vdd \$233679 i1|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28038 VDD|pad|pin1|supply|vdd RD[35]|a2|z a3|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28039 a3|zn$5 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28040 a3|zn$5 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28041 VDD|pad|pin1|supply|vdd RD[0]|a2|z a2|zn$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28042 a2|zn$19 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28043 a2|zn$19 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28044 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28045 a2|zn$20 a2|z$9 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$28046 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28047 a2|zn$20 RD[10]|a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28048 VDD|pad|pin1|supply|vdd RD[33]|a2|z a1|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28049 a1|zn$7 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28050 a1|zn$7 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28051 \$233688 a1|zn$8 \$235386 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$28052 \$235386 a2|zn$16 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$28053 VDD|pad|pin1|supply|vdd \$233688 i1|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28054 VDD|pad|pin1|supply|vdd RD[29]|a2|zn a2|zn$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28055 a2|zn$11 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28056 a2|zn$11 a2|a3|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28057 VDD|pad|pin1|supply|vdd a1|a3|z a3|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28058 a3|zn$6 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$28059 VDD|pad|pin1|supply|vdd a1|z$15 a3|zn$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28060 a3|zn$6 RD[16]|a4|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28061 VDD|pad|pin1|supply|vdd RD[2]|a2|z a3|zn$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28062 a3|zn$7 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28063 a3|zn$7 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28064 VDD|pad|pin1|supply|vdd a3|zn$6 a1|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28065 a1|zn$17 a2|zn$19 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$28066 VDD|pad|pin1|supply|vdd a1|zn$12 a1|zn$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28067 a1|zn$17 a4|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28068 VDD|pad|pin1|supply|vdd a2|zn$24 a1|zn$18 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$28069 a1|zn$18 a1|zn$19 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28070 \$233696 \$233698 \$233695 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28071 \$233696 R[50]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28072 VDD|pad|pin1|supply|vdd i0|i1|q$2 \$233697 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28073 \$233697 s|zn \$233695 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28074 VDD|pad|pin1|supply|vdd s|zn \$233698 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28075 VDD|pad|pin1|supply|vdd \$233695 d|z$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28076 \$233700 \$233702 \$233699 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28077 \$233700 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28078 VDD|pad|pin1|supply|vdd R[7]|i|i0|q \$233701 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28079 \$233701 s|z \$233699 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28080 VDD|pad|pin1|supply|vdd s|z \$233702 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28081 VDD|pad|pin1|supply|vdd \$233699 d|z$15 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28082 \$233704 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28083 VDD|pad|pin1|supply|vdd \$233704 \$233705 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28084 VDD|pad|pin1|supply|vdd \$233705 \$235376 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28085 \$235376 d|z$10 \$233706 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28086 \$233706 \$233704 \$235339 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28087 \$235339 \$233707 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28088 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$235339
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28089 \$233707 \$233706 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28090 \$233707 \$233704 \$233708 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28091 \$233708 \$233705 \$235375 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28092 VDD|pad|pin1|supply|vdd \$233710 \$235375 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28093 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$233710
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28094 VDD|pad|pin1|supply|vdd \$233708 \$233710 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28095 VDD|pad|pin1|supply|vdd \$233710 R[58]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28096 \$235807 \$235806 \$235865 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28097 \$235866 s|zn$2 \$235807 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28098 VDD|pad|pin1|supply|vdd i0|i1|q$5 \$235866 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28099 \$235865 R[37]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28100 \$235806 s|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28101 VDD|pad|pin1|supply|vdd \$235807 d|z$17 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28102 VDD|pad|pin1|supply|vdd cp|z$4 \$235808 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28103 VDD|pad|pin1|supply|vdd \$235808 \$235809 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28104 VDD|pad|pin1|supply|vdd \$236600 \$235810 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28105 \$235868 \$235808 \$235810 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28106 VDD|pad|pin1|supply|vdd \$235809 \$236507 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28107 \$236507 d|z$13 \$235868 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28108 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$235810
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28109 \$235811 \$235809 \$236504 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28110 VDD|pad|pin1|supply|vdd \$236644 \$236504 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28111 VDD|pad|pin1|supply|vdd \$235868 \$236600 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28112 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$236644
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28113 VDD|pad|pin1|supply|vdd \$235811 \$236644 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28114 \$236600 \$235808 \$235811 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28115 VDD|pad|pin1|supply|vdd \$236644 R[55]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28116 VDD|pad|pin1|supply|vdd cp|z$4 \$235812 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28117 VDD|pad|pin1|supply|vdd \$235812 \$235813 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28118 VDD|pad|pin1|supply|vdd \$236601 \$235814 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28119 \$235869 \$235812 \$235814 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28120 VDD|pad|pin1|supply|vdd \$235813 \$236508 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28121 \$236508 d|z$14 \$235869 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28122 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$235814
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28123 \$235815 \$235813 \$236511 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28124 VDD|pad|pin1|supply|vdd \$236645 \$236511 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28125 VDD|pad|pin1|supply|vdd \$235869 \$236601 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28126 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$236645
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28127 VDD|pad|pin1|supply|vdd \$235815 \$236645 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28128 \$236601 \$235812 \$235815 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28129 VDD|pad|pin1|supply|vdd \$236645 R[2]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28130 \$235818 \$235816 \$235870 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28131 \$235871 s|z \$235818 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28132 VDD|pad|pin1|supply|vdd R[6]|i|i0|q \$235871 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28133 \$235870 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28134 \$235816 s|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28135 VDD|pad|pin1|supply|vdd \$235818 d|z$18 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28136 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a2|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28137 VDD|pad|pin1|supply|vdd a2|z$9 a2|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$28138 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28139 VDD|pad|pin1|supply|vdd RD[46]|a4|z a2|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28140 VDD|pad|pin1|supply|vdd a2|zn$22 \$235874 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28141 VDD|pad|pin1|supply|vdd a1|zn$1 \$235874 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28142 VDD|pad|pin1|supply|vdd \$235874 a4|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28143 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28144 VDD|pad|pin1|supply|vdd a2|z$9 a2|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$28145 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28146 VDD|pad|pin1|supply|vdd RD[14]|a4|zn a2|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28147 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28148 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a2|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$28149 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28150 VDD|pad|pin1|supply|vdd RD[22]|a4|zn a2|zn$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28151 VDD|pad|pin1|supply|vdd cp|i|z$2 \$235819 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28152 VDD|pad|pin1|supply|vdd \$235819 \$235820 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28153 VDD|pad|pin1|supply|vdd \$236603 \$235821 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28154 \$235878 \$235819 \$235821 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28155 VDD|pad|pin1|supply|vdd \$235820 \$236524 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28156 \$236524 d|z$20 \$235878 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28157 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$235821
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28158 \$235822 \$235820 \$236527 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28159 VDD|pad|pin1|supply|vdd \$236646 \$236527 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28160 VDD|pad|pin1|supply|vdd \$235878 \$236603 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28161 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$236646
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28162 VDD|pad|pin1|supply|vdd \$235822 \$236646 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28163 \$236603 \$235819 \$235822 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28164 VDD|pad|pin1|supply|vdd \$236646 R[5]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28165 VDD|pad|pin1|supply|vdd RD[3]|a2|z a1|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28166 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28167 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a1|zn$14 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28168 \$235879 a1|zn$18 \$236532 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$28169 VDD|pad|pin1|supply|vdd a2|zn$17 \$236532 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$28170 VDD|pad|pin1|supply|vdd \$235879 i1|z$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28171 VDD|pad|pin1|supply|vdd a1|a3|z a1|zn$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28172 VDD|pad|pin1|supply|vdd a2|z$9 a1|zn$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$28173 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a1|zn$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28174 VDD|pad|pin1|supply|vdd RD[12]|a4|zn a1|zn$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28175 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$24 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28176 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a2|zn$24 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$28177 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$24 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28178 VDD|pad|pin1|supply|vdd RD[20]|a4|zn a2|zn$24 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28179 VDD|pad|pin1|supply|vdd RD[39]|a2|z a1|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28180 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a1|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28181 VDD|pad|pin1|supply|vdd a2|a3|zn$1 a1|zn$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28182 VDD|pad|pin1|supply|vdd RD[24]|a2|z a4|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28183 VDD|pad|pin1|supply|vdd a1|a3|z a4|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28184 VDD|pad|pin1|supply|vdd a2|a3|z$1 a4|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28185 VDD|pad|pin1|supply|vdd RD[27]|a2|zn a2|zn$25 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28186 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$25 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28187 VDD|pad|pin1|supply|vdd a2|a3|z$1 a2|zn$25 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28188 \$235885 a1|zn$20 \$236544 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$28189 VDD|pad|pin1|supply|vdd a2|zn$15 \$236544 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$28190 VDD|pad|pin1|supply|vdd \$235885 i1|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28191 \$235824 \$235823 \$235887 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28192 \$235888 s|zn$1 \$235824 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28193 VDD|pad|pin1|supply|vdd i0|i1|q$4 \$235888 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28194 \$235887 R[63]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28195 \$235823 s|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28196 VDD|pad|pin1|supply|vdd \$235824 d|z$19 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28197 VDD|pad|pin1|supply|vdd cp|i|z$1 \$235825 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28198 VDD|pad|pin1|supply|vdd \$235825 \$235826 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28199 VDD|pad|pin1|supply|vdd \$236605 \$235827 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28200 \$235890 \$235825 \$235827 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28201 VDD|pad|pin1|supply|vdd \$235826 \$236548 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28202 \$236548 d|z$15 \$235890 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28203 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$235827
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28204 \$235828 \$235826 \$236547 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28205 VDD|pad|pin1|supply|vdd \$236647 \$236547 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28206 VDD|pad|pin1|supply|vdd \$235890 \$236605 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28207 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$236647
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28208 VDD|pad|pin1|supply|vdd \$235828 \$236647 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28209 \$236605 \$235825 \$235828 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28210 VDD|pad|pin1|supply|vdd \$236647 R[7]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28211 \$237816 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28212 VDD|pad|pin1|supply|vdd \$237816 \$237799 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28213 VDD|pad|pin1|supply|vdd \$237799 \$239736 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28214 \$239736 d|z$12 \$237817 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28215 \$237817 \$237816 \$239582 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28216 \$239582 \$237818 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28217 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$239582
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28218 \$237818 \$237817 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28219 \$237818 \$237816 \$237800 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28220 \$237800 \$237799 \$239733 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28221 VDD|pad|pin1|supply|vdd \$237820 \$239733 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28222 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$237820
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28223 VDD|pad|pin1|supply|vdd \$237800 \$237820 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28224 VDD|pad|pin1|supply|vdd \$237820 R[60]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28225 \$237822 \$237801 \$237821 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28226 \$237822 R[57]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28227 VDD|pad|pin1|supply|vdd i0|i1|q$6 \$237823 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28228 \$237823 s|zn$1 \$237821 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28229 VDD|pad|pin1|supply|vdd s|zn$1 \$237801 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28230 VDD|pad|pin1|supply|vdd \$237821 d|z$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28231 \$237826 \$237802 \$237825 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28232 \$237826 R[62]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28233 VDD|pad|pin1|supply|vdd i0|i1|q$7 \$237827 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28234 \$237827 s|zn$1 \$237825 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28235 VDD|pad|pin1|supply|vdd s|zn$1 \$237802 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28236 VDD|pad|pin1|supply|vdd \$237825 d|z$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28237 \$237829 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28238 VDD|pad|pin1|supply|vdd \$237829 \$237803 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28239 VDD|pad|pin1|supply|vdd \$237803 \$239731 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28240 \$239731 d|z$18 \$237830 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28241 \$237830 \$237829 \$239583 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28242 \$239583 \$237831 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28243 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$239583
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28244 \$237831 \$237830 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28245 \$237831 \$237829 \$237804 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28246 \$237804 \$237803 \$239729 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28247 VDD|pad|pin1|supply|vdd \$237833 \$239729 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28248 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$237833
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28249 VDD|pad|pin1|supply|vdd \$237804 \$237833 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28250 VDD|pad|pin1|supply|vdd \$237833 R[6]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28251 VDD|pad|pin1|supply|vdd a3|zn$4 i1|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28252 i1|zn$2 a2|zn$21 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$28253 VDD|pad|pin1|supply|vdd a1|z$16 i1|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28254 i1|zn$2 a4|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28255 VDD|pad|pin1|supply|vdd a2|zn$23 \$237834 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28256 \$237834 a1|zn$16 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28257 a1|z$16 \$237834 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28258 \$237836 \$237806 \$237835 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28259 \$237836 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28260 VDD|pad|pin1|supply|vdd R[5]|i|i0|q \$237837 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28261 \$237837 s|z \$237835 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28262 VDD|pad|pin1|supply|vdd s|z \$237806 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28263 VDD|pad|pin1|supply|vdd \$237835 d|z$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28264 \$237838 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28265 VDD|pad|pin1|supply|vdd \$237838 \$237807 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28266 VDD|pad|pin1|supply|vdd \$237807 \$239723 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28267 \$239723 d|z$25 \$237839 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28268 \$237839 \$237838 \$239584 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28269 \$239584 \$237840 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28270 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$239584
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28271 \$237840 \$237839 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28272 \$237840 \$237838 \$237808 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28273 \$237808 \$237807 \$239722 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28274 VDD|pad|pin1|supply|vdd \$237842 \$239722 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28275 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$237842
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28276 VDD|pad|pin1|supply|vdd \$237808 \$237842 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28277 VDD|pad|pin1|supply|vdd \$237842 R[0]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28278 \$237844 \$237809 \$237843 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28279 \$237844 R[61]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28280 VDD|pad|pin1|supply|vdd i0|i1|q$5 \$237845 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28281 \$237845 s|zn$1 \$237843 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28282 VDD|pad|pin1|supply|vdd s|zn$1 \$237809 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28283 VDD|pad|pin1|supply|vdd \$237843 d|z$23 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28284 \$237848 \$237810 \$237847 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28285 \$237848 R[54]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28286 VDD|pad|pin1|supply|vdd i0|i1|q$7 \$237849 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28287 \$237849 s|zn \$237847 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28288 VDD|pad|pin1|supply|vdd s|zn \$237810 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28289 VDD|pad|pin1|supply|vdd \$237847 d|z$24 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28290 VDD|pad|pin1|supply|vdd a1|a2|a4|z s|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28291 s|zn$1 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28292 s|zn$1 a2|a3|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28293 \$237851 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28294 VDD|pad|pin1|supply|vdd \$237851 \$237812 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28295 VDD|pad|pin1|supply|vdd \$237812 \$239718 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28296 \$239718 d|z$26 \$237852 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28297 \$237852 \$237851 \$239585 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28298 \$239585 \$237853 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28299 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$239585
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28300 \$237853 \$237852 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28301 \$237853 \$237851 \$237813 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28302 \$237813 \$237812 \$239719 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28303 VDD|pad|pin1|supply|vdd \$237855 \$239719 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28304 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$237855
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28305 VDD|pad|pin1|supply|vdd \$237813 \$237855 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28306 VDD|pad|pin1|supply|vdd \$237855 R[4]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28307 \$237856 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28308 VDD|pad|pin1|supply|vdd \$237856 \$237814 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28309 VDD|pad|pin1|supply|vdd \$237814 \$239715 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28310 \$239715 d|z$19 \$237857 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28311 \$237857 \$237856 \$239586 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28312 \$239586 \$237858 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28313 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$239586
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28314 \$237858 \$237857 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28315 \$237858 \$237856 \$237815 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28316 \$237815 \$237814 \$239717 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28317 VDD|pad|pin1|supply|vdd \$237860 \$239717 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28318 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$237860
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28319 VDD|pad|pin1|supply|vdd \$237815 \$237860 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28320 VDD|pad|pin1|supply|vdd \$237860 R[63]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28321 VDD|pad|pin1|supply|vdd cp|z$4 \$240235 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28322 VDD|pad|pin1|supply|vdd \$240235 \$240236 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28323 VDD|pad|pin1|supply|vdd \$240571 \$240237 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28324 \$240301 \$240235 \$240237 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28325 VDD|pad|pin1|supply|vdd \$240236 \$240555 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28326 \$240555 d|z$21 \$240301 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28327 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240237
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28328 \$240238 \$240236 \$240552 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28329 VDD|pad|pin1|supply|vdd \$240877 \$240552 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28330 VDD|pad|pin1|supply|vdd \$240301 \$240571 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28331 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240877
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28332 VDD|pad|pin1|supply|vdd \$240238 \$240877 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28333 \$240571 \$240235 \$240238 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28334 VDD|pad|pin1|supply|vdd \$240877 R[57]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28335 VDD|pad|pin1|supply|vdd cp|i|z$2 \$240239 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28336 VDD|pad|pin1|supply|vdd \$240239 \$240240 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28337 VDD|pad|pin1|supply|vdd \$240572 \$240241 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28338 \$240302 \$240239 \$240241 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28339 VDD|pad|pin1|supply|vdd \$240240 \$240565 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28340 \$240565 d|z$22 \$240302 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28341 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240241
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28342 \$240242 \$240240 \$240560 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28343 VDD|pad|pin1|supply|vdd \$240878 \$240560 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28344 VDD|pad|pin1|supply|vdd \$240302 \$240572 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28345 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240878
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28346 VDD|pad|pin1|supply|vdd \$240242 \$240878 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28347 \$240572 \$240239 \$240242 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28348 VDD|pad|pin1|supply|vdd \$240878 R[62]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28349 \$240243 \$240244 \$240303 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28350 \$240304 s|zn \$240243 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28351 VDD|pad|pin1|supply|vdd i0|i1|q$3 \$240304 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28352 \$240303 R[52]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28353 \$240244 s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28354 VDD|pad|pin1|supply|vdd \$240243 d|z$27 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28355 VDD|pad|pin1|supply|vdd cp|i|z$2 \$240245 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28356 VDD|pad|pin1|supply|vdd \$240245 \$240246 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28357 VDD|pad|pin1|supply|vdd \$240573 \$240247 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28358 \$240306 \$240245 \$240247 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28359 VDD|pad|pin1|supply|vdd \$240246 \$240566 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28360 \$240566 d|z$27 \$240306 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28361 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240247
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28362 \$240248 \$240246 \$240561 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28363 VDD|pad|pin1|supply|vdd \$240880 \$240561 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28364 VDD|pad|pin1|supply|vdd \$240306 \$240573 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28365 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240880
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28366 VDD|pad|pin1|supply|vdd \$240248 \$240880 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28367 \$240573 \$240245 \$240248 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28368 VDD|pad|pin1|supply|vdd \$240880 R[52]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28369 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q \$240308 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28370 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q \$240308 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28371 VDD|pad|pin1|supply|vdd \$240308 a2|a3|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28372 VDD|pad|pin1|supply|vdd a2|zn$26 \$240309 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28373 VDD|pad|pin1|supply|vdd a1|zn$15 \$240309 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28374 VDD|pad|pin1|supply|vdd \$240309 a2|z$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28375 VDD|pad|pin1|supply|vdd a2|zn$18 \$240310 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28376 VDD|pad|pin1|supply|vdd a1|zn \$240310 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28377 VDD|pad|pin1|supply|vdd \$240310 a4|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28378 \$240249 \$240250 \$240311 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28379 \$240312 s|z \$240249 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28380 VDD|pad|pin1|supply|vdd R[0]|i|i0|q \$240312 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28381 \$240311 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28382 \$240250 s|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28383 VDD|pad|pin1|supply|vdd \$240249 d|z$25 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28384 VDD|pad|pin1|supply|vdd cp|i|z$3 \$240251 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28385 VDD|pad|pin1|supply|vdd \$240251 \$240252 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28386 VDD|pad|pin1|supply|vdd \$240574 \$240253 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28387 \$240313 \$240251 \$240253 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28388 VDD|pad|pin1|supply|vdd \$240252 \$240545 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28389 \$240545 d|z$23 \$240313 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28390 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240253
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28391 \$240254 \$240252 \$240541 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28392 VDD|pad|pin1|supply|vdd \$240881 \$240541 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28393 VDD|pad|pin1|supply|vdd \$240313 \$240574 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28394 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240881
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28395 VDD|pad|pin1|supply|vdd \$240254 \$240881 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28396 \$240574 \$240251 \$240254 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28397 VDD|pad|pin1|supply|vdd \$240881 R[61]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28398 VDD|pad|pin1|supply|vdd cp|i|z$1 \$240255 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28399 VDD|pad|pin1|supply|vdd \$240255 \$240256 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28400 VDD|pad|pin1|supply|vdd \$240575 \$240257 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28401 \$240314 \$240255 \$240257 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28402 VDD|pad|pin1|supply|vdd \$240256 \$240534 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28403 \$240534 d|z$24 \$240314 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28404 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240257
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28405 \$240258 \$240256 \$240521 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28406 VDD|pad|pin1|supply|vdd \$240882 \$240521 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28407 VDD|pad|pin1|supply|vdd \$240314 \$240575 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28408 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240882
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28409 VDD|pad|pin1|supply|vdd \$240258 \$240882 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28410 \$240575 \$240255 \$240258 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28411 VDD|pad|pin1|supply|vdd \$240882 R[54]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28412 VDD|pad|pin1|supply|vdd a2|zn$25 a1|zn$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$28413 VDD|pad|pin1|supply|vdd a1|zn$11 a1|zn$20 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28414 \$240259 \$240260 \$240315 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28415 \$240316 s|zn \$240259 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28416 VDD|pad|pin1|supply|vdd i0|i1|q$6 \$240316 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28417 \$240315 R[49]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28418 \$240260 s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28419 VDD|pad|pin1|supply|vdd \$240259 d|z$28 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28420 VDD|pad|pin1|supply|vdd cp|i|z$1 \$240261 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28421 VDD|pad|pin1|supply|vdd \$240261 \$240262 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28422 VDD|pad|pin1|supply|vdd \$240576 \$240263 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28423 \$240318 \$240261 \$240263 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28424 VDD|pad|pin1|supply|vdd \$240262 \$240515 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28425 \$240515 d|z$28 \$240318 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28426 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240263
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28427 \$240264 \$240262 \$240503 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28428 VDD|pad|pin1|supply|vdd \$240883 \$240503 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28429 VDD|pad|pin1|supply|vdd \$240318 \$240576 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28430 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$240883
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28431 VDD|pad|pin1|supply|vdd \$240264 \$240883 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28432 \$240576 \$240261 \$240264 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28433 VDD|pad|pin1|supply|vdd \$240883 R[49]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28434 \$242202 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28435 VDD|pad|pin1|supply|vdd \$242202 \$242148 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28436 VDD|pad|pin1|supply|vdd \$242148 \$244436 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28437 \$244436 d|z$9 \$242203 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28438 \$242203 \$242202 \$243744 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28439 \$243744 \$242204 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28440 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$243744
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28441 \$242204 \$242203 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28442 \$242204 \$242202 \$242149 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28443 \$242149 \$242148 \$244450 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28444 VDD|pad|pin1|supply|vdd \$242206 \$244450 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28445 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$242206
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28446 VDD|pad|pin1|supply|vdd \$242149 \$242206 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28447 VDD|pad|pin1|supply|vdd \$242206 R[35]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28448 \$242207 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28449 VDD|pad|pin1|supply|vdd \$242207 \$242150 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28450 VDD|pad|pin1|supply|vdd \$242150 \$244469 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28451 \$244469 d|z$29 \$242209 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28452 \$242209 \$242207 \$243745 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28453 \$243745 \$242210 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28454 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$243745
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28455 \$242210 \$242209 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28456 \$242210 \$242207 \$242151 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28457 \$242151 \$242150 \$244492 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28458 VDD|pad|pin1|supply|vdd \$242212 \$244492 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28459 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$242212
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28460 VDD|pad|pin1|supply|vdd \$242151 \$242212 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28461 VDD|pad|pin1|supply|vdd \$242212 R[34]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28462 \$242215 \$242152 \$242214 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28463 \$242215 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28464 VDD|pad|pin1|supply|vdd R[30]|i0|q \$242216 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28465 \$242216 s|z$1 \$242214 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28466 VDD|pad|pin1|supply|vdd s|z$1 \$242152 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28467 VDD|pad|pin1|supply|vdd \$242214 d|z$30 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28468 \$242219 \$243746 \$242218 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28469 \$242219 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28470 VDD|pad|pin1|supply|vdd R[27]|i0|q \$242220 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28471 \$242220 s|z$1 \$242218 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28472 VDD|pad|pin1|supply|vdd s|z$1 \$243746 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28473 VDD|pad|pin1|supply|vdd \$242218 d|z$31 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28474 z$28 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$28475 VDD|pad|pin1|supply|vdd RD[36]|a2|z a3|zn$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28476 a3|zn$1 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28477 a3|zn$1 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28478 \$242224 \$242156 \$242223 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28479 \$242224 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28480 VDD|pad|pin1|supply|vdd R[28]|i0|q \$242226 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28481 \$242226 s|z$1 \$242223 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28482 VDD|pad|pin1|supply|vdd s|z$1 \$242156 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28483 VDD|pad|pin1|supply|vdd \$242223 d|z$32 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28484 cp|i|z$2 \$242228 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$28485 VDD|pad|pin1|supply|vdd i|z$115 \$242228 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$28486 \$242230 \$242157 \$242229 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28487 \$242230 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28488 VDD|pad|pin1|supply|vdd R[31]|i0|q \$242232 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28489 \$242232 s|z$1 \$242229 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28490 VDD|pad|pin1|supply|vdd s|z$1 \$242157 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28491 VDD|pad|pin1|supply|vdd \$242229 d|z$33 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28492 \$242234 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28493 VDD|pad|pin1|supply|vdd \$242234 \$242158 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28494 VDD|pad|pin1|supply|vdd \$242158 \$244527 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28495 \$244527 d|z$34 \$242236 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28496 \$242236 \$242234 \$243747 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28497 \$243747 \$242237 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28498 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$243747
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28499 \$242237 \$242236 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28500 \$242237 \$242234 \$242159 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28501 \$242159 \$242158 \$244515 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28502 VDD|pad|pin1|supply|vdd \$242239 \$244515 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28503 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$242239
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28504 VDD|pad|pin1|supply|vdd \$242159 \$242239 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28505 VDD|pad|pin1|supply|vdd \$242239 R[39]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28506 \$242241 \$242160 \$242240 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28507 \$242241 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28508 VDD|pad|pin1|supply|vdd R[25]|i0|q \$242243 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28509 \$242243 s|z$1 \$242240 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28510 VDD|pad|pin1|supply|vdd s|z$1 \$242160 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28511 VDD|pad|pin1|supply|vdd \$242240 d|z$35 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28512 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q s|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28513 s|zn a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$28514 VDD|pad|pin1|supply|vdd a1|z$15 s|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$28515 s|zn a1|a2|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28516 VDD|pad|pin1|supply|vdd a1|a2|a4|z s|zn$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28517 s|zn$2 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28518 s|zn$2 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28519 \$242246 \$242163 \$242245 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28520 \$242246 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28521 VDD|pad|pin1|supply|vdd R[4]|i|i0|q \$242247 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28522 \$242247 s|z \$242245 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28523 VDD|pad|pin1|supply|vdd s|z \$242163 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28524 VDD|pad|pin1|supply|vdd \$242245 d|z$26 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28525 VDD|pad|pin1|supply|vdd RD[32]|a2|z a2|zn$27 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28526 a2|zn$27 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28527 a2|zn$27 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28528 \$242250 \$243748 \$242249 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28529 \$242250 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28530 VDD|pad|pin1|supply|vdd R[1]|i|i0|q \$242251 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28531 \$242251 s|z \$242249 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28532 VDD|pad|pin1|supply|vdd s|z \$243748 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28533 VDD|pad|pin1|supply|vdd \$242249 d|z$36 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28534 \$242253 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28535 VDD|pad|pin1|supply|vdd \$242253 \$242165 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28536 VDD|pad|pin1|supply|vdd \$242165 \$244481 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28537 \$244481 d|z$37 \$242255 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28538 \$242255 \$242253 \$243749 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28539 \$243749 \$242256 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28540 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$243749
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28541 \$242256 \$242255 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28542 \$242256 \$242253 \$242166 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28543 \$242166 \$242165 \$244475 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28544 VDD|pad|pin1|supply|vdd \$242258 \$244475 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28545 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$242258
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28546 VDD|pad|pin1|supply|vdd \$242166 \$242258 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28547 VDD|pad|pin1|supply|vdd \$242258 R[3]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28548 \$244529 \$244530 \$244563 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28549 \$244564 s|zn$2 \$244529 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28550 VDD|pad|pin1|supply|vdd i0|i1|q$7 \$244564 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28551 \$244563 R[38]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28552 \$244530 s|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28553 VDD|pad|pin1|supply|vdd \$244529 d|z$38 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28554 \$244531 \$244532 \$244566 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28555 \$244567 s|zn$3 \$244531 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28556 VDD|pad|pin1|supply|vdd R[45]|i0|q \$244567 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28557 \$244566 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28558 \$244532 s|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28559 VDD|pad|pin1|supply|vdd \$244531 d|z$39 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28560 VDD|pad|pin1|supply|vdd i|z$115 \$244534 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$28561 VDD|pad|pin1|supply|vdd \$244534 cp|z$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$28562 VDD|pad|pin1|supply|vdd cp|i|z$2 \$244535 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28563 VDD|pad|pin1|supply|vdd \$244535 \$244536 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28564 VDD|pad|pin1|supply|vdd \$244833 \$244537 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28565 \$244569 \$244535 \$244537 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28566 VDD|pad|pin1|supply|vdd \$244536 \$244831 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28567 \$244831 d|z$30 \$244569 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28568 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$244537
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28569 \$244538 \$244536 \$244830 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28570 VDD|pad|pin1|supply|vdd \$245494 \$244830 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28571 VDD|pad|pin1|supply|vdd \$244569 \$244833 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28572 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$245494
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28573 VDD|pad|pin1|supply|vdd \$244538 \$245494 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28574 \$244833 \$244535 \$244538 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28575 VDD|pad|pin1|supply|vdd \$245494 R[30]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28576 VDD|pad|pin1|supply|vdd cp|i|z$2 \$244539 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28577 VDD|pad|pin1|supply|vdd \$244539 \$244540 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28578 VDD|pad|pin1|supply|vdd \$244834 \$244541 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28579 \$244570 \$244539 \$244541 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28580 VDD|pad|pin1|supply|vdd \$244540 \$244829 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28581 \$244829 d|z$31 \$244570 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28582 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$244541
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28583 \$244542 \$244540 \$244828 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28584 VDD|pad|pin1|supply|vdd \$245495 \$244828 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28585 VDD|pad|pin1|supply|vdd \$244570 \$244834 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28586 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$245495
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28587 VDD|pad|pin1|supply|vdd \$244542 \$245495 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28588 \$244834 \$244539 \$244542 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28589 VDD|pad|pin1|supply|vdd \$245495 R[27]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28590 VDD|pad|pin1|supply|vdd RD[31]|a2|zn a3|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28591 VDD|pad|pin1|supply|vdd a1|a3|z a3|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28592 VDD|pad|pin1|supply|vdd a2|a3|z$1 a3|zn$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28593 VDD|pad|pin1|supply|vdd cp|i|z$2 \$244543 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28594 VDD|pad|pin1|supply|vdd \$244543 \$244544 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28595 VDD|pad|pin1|supply|vdd \$244835 \$244545 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28596 \$244571 \$244543 \$244545 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28597 VDD|pad|pin1|supply|vdd \$244544 \$244827 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28598 \$244827 d|z$33 \$244571 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28599 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$244545
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28600 \$244546 \$244544 \$244825 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28601 VDD|pad|pin1|supply|vdd \$245496 \$244825 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28602 VDD|pad|pin1|supply|vdd \$244571 \$244835 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28603 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$245496
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28604 VDD|pad|pin1|supply|vdd \$244546 \$245496 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28605 \$244835 \$244543 \$244546 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28606 VDD|pad|pin1|supply|vdd \$245496 R[31]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28607 VDD|pad|pin1|supply|vdd cp|i|z$3 \$244547 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28608 VDD|pad|pin1|supply|vdd \$244547 \$244548 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28609 VDD|pad|pin1|supply|vdd \$244836 \$244549 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28610 \$244572 \$244547 \$244549 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28611 VDD|pad|pin1|supply|vdd \$244548 \$244824 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28612 \$244824 d|z$40 \$244572 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28613 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$244549
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28614 \$244550 \$244548 \$244822 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28615 VDD|pad|pin1|supply|vdd \$245497 \$244822 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28616 VDD|pad|pin1|supply|vdd \$244572 \$244836 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28617 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$245497
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28618 VDD|pad|pin1|supply|vdd \$244550 \$245497 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28619 \$244836 \$244547 \$244550 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28620 VDD|pad|pin1|supply|vdd \$245497 R[32]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28621 VDD|pad|pin1|supply|vdd cp|i|z$3 \$244551 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28622 VDD|pad|pin1|supply|vdd \$244551 \$244552 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28623 VDD|pad|pin1|supply|vdd \$244837 \$244553 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28624 \$244574 \$244551 \$244553 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28625 VDD|pad|pin1|supply|vdd \$244552 \$244820 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28626 \$244820 d|z$35 \$244574 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28627 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$244553
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28628 \$244554 \$244552 \$244816 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28629 VDD|pad|pin1|supply|vdd \$245498 \$244816 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28630 VDD|pad|pin1|supply|vdd \$244574 \$244837 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28631 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$245498
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28632 VDD|pad|pin1|supply|vdd \$244554 \$245498 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28633 \$244837 \$244551 \$244554 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28634 VDD|pad|pin1|supply|vdd \$245498 R[25]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28635 VDD|pad|pin1|supply|vdd a2|a3|zn$1 \$244575 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28636 VDD|pad|pin1|supply|vdd a1|a3|z \$244575 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28637 VDD|pad|pin1|supply|vdd \$244575 a2|z$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28638 VDD|pad|pin1|supply|vdd cp|i|z$1 \$244555 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28639 VDD|pad|pin1|supply|vdd \$244555 \$244556 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28640 VDD|pad|pin1|supply|vdd \$244838 \$244557 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28641 \$244577 \$244555 \$244557 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28642 VDD|pad|pin1|supply|vdd \$244556 \$244815 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28643 \$244815 d|z$41 \$244577 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28644 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$244557
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28645 \$244558 \$244556 \$244814 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28646 VDD|pad|pin1|supply|vdd \$245499 \$244814 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28647 VDD|pad|pin1|supply|vdd \$244577 \$244838 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28648 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$245499
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28649 VDD|pad|pin1|supply|vdd \$244558 \$245499 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28650 \$244838 \$244555 \$244558 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28651 VDD|pad|pin1|supply|vdd \$245499 R[33]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28652 z$29 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$28653 VDD|pad|pin1|supply|vdd cp|i|z$1 \$244559 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28654 VDD|pad|pin1|supply|vdd \$244559 \$244560 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28655 VDD|pad|pin1|supply|vdd \$244839 \$244561 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28656 \$244579 \$244559 \$244561 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28657 VDD|pad|pin1|supply|vdd \$244560 \$244813 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28658 \$244813 d|z$36 \$244579 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28659 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$244561
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28660 \$244562 \$244560 \$244812 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28661 VDD|pad|pin1|supply|vdd \$245500 \$244812 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28662 VDD|pad|pin1|supply|vdd \$244579 \$244839 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28663 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$245500
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28664 VDD|pad|pin1|supply|vdd \$244562 \$245500 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28665 \$244839 \$244559 \$244562 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28666 VDD|pad|pin1|supply|vdd \$245500 R[1]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28667 VDD|pad|pin1|supply|vdd cp|z$4 \$249100 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28668 VDD|pad|pin1|supply|vdd \$249100 \$249101 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28669 \$246601 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28670 VDD|pad|pin1|supply|vdd \$246601 \$246550 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28671 VDD|pad|pin1|supply|vdd \$249189 \$249103 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28672 \$249102 \$249100 \$249103 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28673 VDD|pad|pin1|supply|vdd \$249101 \$249679 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28674 \$249679 d|z$38 \$249102 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28675 VDD|pad|pin1|supply|vdd \$246550 \$248955 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28676 \$248955 d|z$17 \$246602 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28677 \$246602 \$246601 \$248106 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28678 \$248106 \$246603 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28679 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$249103
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28680 \$249104 \$249101 \$249185 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28681 VDD|pad|pin1|supply|vdd \$249190 \$249185 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28682 VDD|pad|pin1|supply|vdd \$249102 \$249189 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28683 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$249190
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28684 VDD|pad|pin1|supply|vdd \$249104 \$249190 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28685 \$249189 \$249100 \$249104 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28686 VDD|pad|pin1|supply|vdd \$249190 R[38]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28687 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$248106
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28688 \$246603 \$246602 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28689 \$246603 \$246601 \$246551 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28690 \$246551 \$246550 \$248959 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28691 VDD|pad|pin1|supply|vdd \$246605 \$248959 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28692 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$246605
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28693 VDD|pad|pin1|supply|vdd \$246551 \$246605 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28694 VDD|pad|pin1|supply|vdd \$246605 R[37]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28695 \$246607 \$246552 \$246606 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28696 \$246607 R[34]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28697 VDD|pad|pin1|supply|vdd i0|i1|q$2 \$246608 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28698 \$246608 s|zn$2 \$246606 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28699 \$249105 \$249094 \$249106 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28700 \$249107 s|zn$4 \$249105 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28701 VDD|pad|pin1|supply|vdd R[15]|i|i0|q \$249107 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28702 \$249106 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28703 VDD|pad|pin1|supply|vdd s|zn$2 \$246552 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28704 VDD|pad|pin1|supply|vdd \$246606 d|z$29 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28705 \$249094 s|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28706 VDD|pad|pin1|supply|vdd \$249105 d|z$45 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28707 \$246610 \$246554 \$246609 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28708 \$246610 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28709 VDD|pad|pin1|supply|vdd R[12]|i|i0|q \$246611 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28710 \$246611 s|zn$4 \$246609 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28711 VDD|pad|pin1|supply|vdd cp|z$4 \$249109 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28712 VDD|pad|pin1|supply|vdd \$249109 \$249110 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28713 VDD|pad|pin1|supply|vdd \$249191 \$249112 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28714 \$249111 \$249109 \$249112 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28715 VDD|pad|pin1|supply|vdd \$249110 \$249686 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28716 \$249686 d|z$45 \$249111 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28717 VDD|pad|pin1|supply|vdd s|zn$4 \$246554 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28718 VDD|pad|pin1|supply|vdd \$246609 d|z$42 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28719 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$249112
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28720 \$249113 \$249110 \$249184 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28721 VDD|pad|pin1|supply|vdd \$249192 \$249184 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28722 VDD|pad|pin1|supply|vdd \$249111 \$249191 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28723 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$249192
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28724 VDD|pad|pin1|supply|vdd \$249113 \$249192 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28725 \$249191 \$249109 \$249113 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28726 VDD|pad|pin1|supply|vdd \$249192 R[15]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28727 VDD|pad|pin1|supply|vdd RD[5]|a2|zn a1|zn$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28728 a1|zn$4 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28729 a1|zn$4 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28730 \$246614 \$246556 \$246613 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28731 \$246614 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28732 VDD|pad|pin1|supply|vdd R[11]|i|i0|q \$246615 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28733 \$246615 s|zn$4 \$246613 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28734 VDD|pad|pin1|supply|vdd cp|i|z$2 \$249114 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28735 VDD|pad|pin1|supply|vdd \$249114 \$249115 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28736 VDD|pad|pin1|supply|vdd s|zn$4 \$246556 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28737 VDD|pad|pin1|supply|vdd \$246613 d|z$43 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28738 VDD|pad|pin1|supply|vdd \$249193 \$249117 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28739 \$249116 \$249114 \$249117 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28740 VDD|pad|pin1|supply|vdd \$249115 \$249690 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28741 \$249690 d|z$43 \$249116 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28742 \$246617 cp|i|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28743 VDD|pad|pin1|supply|vdd \$246617 \$246557 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28744 VDD|pad|pin1|supply|vdd \$246557 \$248981 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28745 \$248981 d|z$32 \$246618 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28746 \$246618 \$246617 \$248107 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28747 \$248107 \$246619 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28748 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$249117
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28749 \$249118 \$249115 \$249183 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28750 VDD|pad|pin1|supply|vdd \$249194 \$249183 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28751 VDD|pad|pin1|supply|vdd \$249116 \$249193 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28752 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$249194
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28753 VDD|pad|pin1|supply|vdd \$249118 \$249194 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28754 \$249193 \$249114 \$249118 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28755 VDD|pad|pin1|supply|vdd \$249194 R[11]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28756 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$248107
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28757 \$246619 \$246618 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28758 \$246619 \$246617 \$246558 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28759 \$246558 \$246557 \$248985 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28760 VDD|pad|pin1|supply|vdd \$246621 \$248985 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28761 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$246621
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28762 VDD|pad|pin1|supply|vdd \$246558 \$246621 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28763 VDD|pad|pin1|supply|vdd \$246621 R[28]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28764 a1|z$15 a1|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$28765 a2|a3|zn$1 a1|i|i0|i1|q \$248996 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$28766 \$248996 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$28767 \$246623 \$246559 \$246622 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28768 \$246623 R[39]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28769 VDD|pad|pin1|supply|vdd i0|i1|q$4 \$246624 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28770 \$246624 s|zn$2 \$246622 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28771 \$249119 \$249095 \$249120 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28772 \$249121 s|z$1 \$249119 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28773 VDD|pad|pin1|supply|vdd R[24]|i0|q \$249121 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28774 \$249120 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28775 VDD|pad|pin1|supply|vdd s|zn$2 \$246559 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28776 VDD|pad|pin1|supply|vdd \$246622 d|z$34 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28777 \$249095 s|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28778 VDD|pad|pin1|supply|vdd \$249119 d|z$46 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28779 \$246626 \$246560 \$246625 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28780 \$246626 R[32]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28781 VDD|pad|pin1|supply|vdd i0|i1|q \$246627 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28782 \$246627 s|zn$2 \$246625 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28783 \$249123 \$249096 \$249124 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28784 \$249125 s|zn$4 \$249123 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28785 VDD|pad|pin1|supply|vdd R[14]|i|i0|q \$249125 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28786 \$249124 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28787 VDD|pad|pin1|supply|vdd s|zn$2 \$246560 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28788 VDD|pad|pin1|supply|vdd \$246625 d|z$40 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28789 \$249096 s|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28790 VDD|pad|pin1|supply|vdd \$249123 d|z$47 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28791 z$30 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$28792 \$249127 \$249097 \$249128 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28793 \$249129 s|z$1 \$249127 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28794 VDD|pad|pin1|supply|vdd R[29]|i0|q \$249129 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28795 \$249128 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28796 cp|i|z$3 \$246629 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$28797 VDD|pad|pin1|supply|vdd i|z$115 \$246629 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$28798 VDD|pad|pin1|supply|vdd a2|a3|z$1 \$246631 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28799 \$246631 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28800 \$249097 s|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28801 VDD|pad|pin1|supply|vdd \$249127 d|z$48 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28802 a2|z$12 \$246631 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28803 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q a2|zn$28 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28804 VDD|pad|pin1|supply|vdd a1|z$15 a2|zn$28 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28805 VDD|pad|pin1|supply|vdd a2|z$12 \$246633 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28806 \$246633 a1|a2|a4|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28807 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$28 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28808 s|z$1 \$246633 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28809 VDD|pad|pin1|supply|vdd a2|z$9 a2|zn$29 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28810 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$29 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28811 VDD|pad|pin1|supply|vdd a1|a3|z a2|zn$29 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28812 \$246635 \$246561 \$246634 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28813 \$246635 R[36]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28814 VDD|pad|pin1|supply|vdd i0|i1|q$3 \$246636 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28815 \$246636 s|zn$2 \$246634 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28816 VDD|pad|pin1|supply|vdd a2|z$11 \$249133 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28817 VDD|pad|pin1|supply|vdd a1|a2|a4|z \$249133 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28818 VDD|pad|pin1|supply|vdd \$249133 s|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$28819 VDD|pad|pin1|supply|vdd s|zn$2 \$246561 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28820 VDD|pad|pin1|supply|vdd \$246634 d|z$44 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28821 \$249134 \$249098 \$249135 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28822 \$249136 s|zn$2 \$249134 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28823 VDD|pad|pin1|supply|vdd i0|i1|q$6 \$249136 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28824 \$249135 R[33]|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28825 \$246638 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28826 VDD|pad|pin1|supply|vdd \$246638 \$246562 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28827 VDD|pad|pin1|supply|vdd \$246562 \$249026 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28828 \$249026 d|z$44 \$246639 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28829 \$246639 \$246638 \$248108 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28830 \$248108 \$246640 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28831 \$249098 s|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28832 VDD|pad|pin1|supply|vdd \$249134 d|z$41 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28833 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$248108
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28834 \$246640 \$246639 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28835 \$246640 \$246638 \$246563 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28836 \$246563 \$246562 \$249029 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28837 VDD|pad|pin1|supply|vdd \$246642 \$249029 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28838 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$246642
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28839 VDD|pad|pin1|supply|vdd \$246563 \$246642 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28840 VDD|pad|pin1|supply|vdd \$246642 R[36]|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28841 \$249137 \$249099 \$249138 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$28842 \$249139 s|zn$4 \$249137 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28843 VDD|pad|pin1|supply|vdd R[9]|i|i0|q \$249139 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28844 \$249138 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28845 \$246644 \$246564 \$246643 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28846 \$246644 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28847 VDD|pad|pin1|supply|vdd R[3]|i|i0|q \$246645 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28848 \$246645 s|z \$246643 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28849 \$249099 s|zn$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$28850 VDD|pad|pin1|supply|vdd \$249137 d|z$49 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28851 VDD|pad|pin1|supply|vdd cp|i|z$1 \$249141 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28852 VDD|pad|pin1|supply|vdd \$249141 \$249142 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28853 VDD|pad|pin1|supply|vdd s|z \$246564 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28854 VDD|pad|pin1|supply|vdd \$246643 d|z$37 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28855 VDD|pad|pin1|supply|vdd \$249197 \$249144 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28856 \$249143 \$249141 \$249144 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28857 VDD|pad|pin1|supply|vdd \$249142 \$249717 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28858 \$249717 d|z$49 \$249143 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28859 cp|i|z$1 \$246646 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$28860 VDD|pad|pin1|supply|vdd i|z$115 \$246646 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$28861 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$249144
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28862 \$249145 \$249142 \$249182 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28863 VDD|pad|pin1|supply|vdd \$249198 \$249182 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28864 VDD|pad|pin1|supply|vdd \$249143 \$249197 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28865 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$249198
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28866 VDD|pad|pin1|supply|vdd \$249145 \$249198 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28867 \$249197 \$249141 \$249145 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28868 VDD|pad|pin1|supply|vdd \$249198 R[9]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28869 \$251080 \$250812 \$251079 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28870 \$251080 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28871 VDD|pad|pin1|supply|vdd R[42]|i0|q \$251081 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28872 \$251081 s|zn$3 \$251079 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28873 VDD|pad|pin1|supply|vdd s|zn$3 \$250812 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28874 VDD|pad|pin1|supply|vdd \$251079 d|z$50 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28875 \$251084 \$250813 \$251083 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28876 \$251084 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28877 VDD|pad|pin1|supply|vdd R[13]|i|i0|q \$251085 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28878 \$251085 s|zn$4 \$251083 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28879 VDD|pad|pin1|supply|vdd s|zn$4 \$250813 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28880 VDD|pad|pin1|supply|vdd \$251083 d|z$51 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28881 \$251087 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28882 VDD|pad|pin1|supply|vdd \$251087 \$250814 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28883 VDD|pad|pin1|supply|vdd \$250814 \$252785 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28884 \$252785 d|z$51 \$251088 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28885 \$251088 \$251087 \$252728 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28886 \$252728 \$251089 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28887 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$252728
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28888 \$251089 \$251088 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28889 \$251089 \$251087 \$250815 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28890 \$250815 \$250814 \$252784 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28891 VDD|pad|pin1|supply|vdd \$251091 \$252784 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28892 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$251091
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28893 VDD|pad|pin1|supply|vdd \$250815 \$251091 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28894 VDD|pad|pin1|supply|vdd \$251091 R[13]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28895 \$251093 \$250816 \$251092 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28896 \$251093 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28897 VDD|pad|pin1|supply|vdd R[44]|i0|q \$251094 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28898 \$251094 s|zn$3 \$251092 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28899 VDD|pad|pin1|supply|vdd s|zn$3 \$250816 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28900 VDD|pad|pin1|supply|vdd \$251092 d|z$52 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28901 VDD|pad|pin1|supply|vdd RD[7]|a2|zn a2|zn$26 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$28902 a2|zn$26 a1|a3|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$28903 a2|zn$26 a2|a3|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$28904 \$251097 \$250818 \$251096 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28905 \$251097 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28906 VDD|pad|pin1|supply|vdd R[8]|i|i0|q \$251098 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28907 \$251098 s|zn$4 \$251096 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28908 VDD|pad|pin1|supply|vdd s|zn$4 \$250818 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28909 VDD|pad|pin1|supply|vdd \$251096 d|z$53 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28910 a1|a3|z a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$28911 a2|z$9 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$28912 \$251101 \$250819 \$251100 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28913 \$251101 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28914 VDD|pad|pin1|supply|vdd R[26]|i0|q \$251102 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28915 \$251102 s|z$1 \$251100 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28916 VDD|pad|pin1|supply|vdd s|z$1 \$250819 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28917 VDD|pad|pin1|supply|vdd \$251100 d|z$54 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28918 \$251104 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28919 VDD|pad|pin1|supply|vdd \$251104 \$250820 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28920 VDD|pad|pin1|supply|vdd \$250820 \$252779 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28921 \$252779 d|z$46 \$251105 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28922 \$251105 \$251104 \$252729 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28923 \$252729 \$251106 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28924 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$252729
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28925 \$251106 \$251105 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28926 \$251106 \$251104 \$250821 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28927 \$250821 \$250820 \$252776 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28928 VDD|pad|pin1|supply|vdd \$251108 \$252776 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28929 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$251108
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28930 VDD|pad|pin1|supply|vdd \$250821 \$251108 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28931 VDD|pad|pin1|supply|vdd \$251108 R[24]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28932 \$251109 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28933 VDD|pad|pin1|supply|vdd \$251109 \$250822 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28934 VDD|pad|pin1|supply|vdd \$250822 \$252775 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28935 \$252775 d|z$48 \$251110 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28936 \$251110 \$251109 \$252730 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28937 \$252730 \$251111 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28938 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$252730
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28939 \$251111 \$251110 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28940 \$251111 \$251109 \$250823 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28941 \$250823 \$250822 \$252773 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28942 VDD|pad|pin1|supply|vdd \$251113 \$252773 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28943 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$251113
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28944 VDD|pad|pin1|supply|vdd \$250823 \$251113 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28945 VDD|pad|pin1|supply|vdd \$251113 R[29]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28946 \$251114 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28947 VDD|pad|pin1|supply|vdd \$251114 \$250824 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28948 VDD|pad|pin1|supply|vdd \$250824 \$252771 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28949 \$252771 d|z$56 \$251115 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28950 \$251115 \$251114 \$252731 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28951 \$252731 \$251116 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28952 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$252731
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28953 \$251116 \$251115 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28954 \$251116 \$251114 \$250825 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28955 \$250825 \$250824 \$252772 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28956 VDD|pad|pin1|supply|vdd \$251118 \$252772 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28957 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$251118
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28958 VDD|pad|pin1|supply|vdd \$250825 \$251118 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28959 VDD|pad|pin1|supply|vdd \$251118 R[41]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28960 \$251120 \$250826 \$251119 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$28961 \$251120 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$28962 VDD|pad|pin1|supply|vdd R[10]|i|i0|q \$251121 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$28963 \$251121 s|zn$4 \$251119 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$28964 VDD|pad|pin1|supply|vdd s|zn$4 \$250826 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$28965 VDD|pad|pin1|supply|vdd \$251119 d|z$55 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$28966 \$251124 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$28967 VDD|pad|pin1|supply|vdd \$251124 \$250827 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28968 VDD|pad|pin1|supply|vdd \$250827 \$252768 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28969 \$252768 d|z$55 \$251125 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28970 \$251125 \$251124 \$252732 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28971 \$252732 \$251126 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$28972 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$252732
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28973 \$251126 \$251125 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$28974 \$251126 \$251124 \$250828 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28975 \$250828 \$250827 \$252764 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28976 VDD|pad|pin1|supply|vdd \$251128 \$252764 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28977 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$251128
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28978 VDD|pad|pin1|supply|vdd \$250828 \$251128 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28979 VDD|pad|pin1|supply|vdd \$251128 R[10]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28980 VDD|pad|pin1|supply|vdd cp|z$4 \$252801 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28981 VDD|pad|pin1|supply|vdd \$252801 \$252802 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28982 VDD|pad|pin1|supply|vdd \$253476 \$252803 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28983 \$253378 \$252801 \$252803 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28984 VDD|pad|pin1|supply|vdd \$252802 \$253472 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28985 \$253472 d|z$39 \$253378 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$28986 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$252803
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$28987 \$252804 \$252802 \$253304 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$28988 VDD|pad|pin1|supply|vdd \$253477 \$253304 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$28989 VDD|pad|pin1|supply|vdd \$253378 \$253476 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$28990 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$253477
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$28991 VDD|pad|pin1|supply|vdd \$252804 \$253477 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$28992 \$253476 \$252801 \$252804 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$28993 VDD|pad|pin1|supply|vdd \$253477 R[45]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$28994 VDD|pad|pin1|supply|vdd cp|z$4 \$252805 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28995 VDD|pad|pin1|supply|vdd \$252805 \$252806 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$28996 VDD|pad|pin1|supply|vdd \$253478 \$252807 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$28997 \$253379 \$252805 \$252807 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$28998 VDD|pad|pin1|supply|vdd \$252806 \$253469 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$28999 \$253469 d|z$42 \$253379 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29000 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$252807
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29001 \$252808 \$252806 \$253319 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29002 VDD|pad|pin1|supply|vdd \$253479 \$253319 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29003 VDD|pad|pin1|supply|vdd \$253379 \$253478 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29004 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$253479
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29005 VDD|pad|pin1|supply|vdd \$252808 \$253479 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29006 \$253478 \$252805 \$252808 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29007 VDD|pad|pin1|supply|vdd \$253479 R[12]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29008 VDD|pad|pin1|supply|vdd cp|i|z$2 \$252809 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29009 VDD|pad|pin1|supply|vdd \$252809 \$252810 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29010 VDD|pad|pin1|supply|vdd \$253480 \$252811 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29011 \$253380 \$252809 \$252811 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29012 VDD|pad|pin1|supply|vdd \$252810 \$253468 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29013 \$253468 d|z$53 \$253380 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29014 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$252811
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29015 \$252812 \$252810 \$253349 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29016 VDD|pad|pin1|supply|vdd \$253481 \$253349 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29017 VDD|pad|pin1|supply|vdd \$253380 \$253480 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29018 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$253481
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29019 VDD|pad|pin1|supply|vdd \$252812 \$253481 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29020 \$253480 \$252809 \$252812 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29021 VDD|pad|pin1|supply|vdd \$253481 R[8]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29022 VDD|pad|pin1|supply|vdd cp|i|z$2 \$252813 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29023 VDD|pad|pin1|supply|vdd \$252813 \$252814 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29024 VDD|pad|pin1|supply|vdd \$253482 \$252815 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29025 \$253381 \$252813 \$252815 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29026 VDD|pad|pin1|supply|vdd \$252814 \$253467 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29027 \$253467 d|z$54 \$253381 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29028 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$252815
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29029 \$252816 \$252814 \$253369 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29030 VDD|pad|pin1|supply|vdd \$253483 \$253369 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29031 VDD|pad|pin1|supply|vdd \$253381 \$253482 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29032 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$253483
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29033 VDD|pad|pin1|supply|vdd \$252816 \$253483 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29034 \$253482 \$252813 \$252816 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29035 VDD|pad|pin1|supply|vdd \$253483 R[26]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29036 VDD|pad|pin1|supply|vdd cp|i|z$3 \$252817 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29037 VDD|pad|pin1|supply|vdd \$252817 \$252818 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29038 VDD|pad|pin1|supply|vdd \$253484 \$252819 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29039 \$253382 \$252817 \$252819 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29040 VDD|pad|pin1|supply|vdd \$252818 \$253466 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29041 \$253466 d|z$47 \$253382 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29042 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$252819
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29043 \$252820 \$252818 \$253374 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29044 VDD|pad|pin1|supply|vdd \$253485 \$253374 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29045 VDD|pad|pin1|supply|vdd \$253382 \$253484 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29046 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$253485
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29047 VDD|pad|pin1|supply|vdd \$252820 \$253485 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29048 \$253484 \$252817 \$252820 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29049 VDD|pad|pin1|supply|vdd \$253485 R[14]|i|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29050 VDD|pad|pin1|supply|vdd a2|z$9 a2|zn$30 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29051 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a2|zn$30 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29052 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a2|zn$30 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29053 \$252821 \$252822 \$253384 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29054 \$253385 s|zn$3 \$252821 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29055 VDD|pad|pin1|supply|vdd R[41]|i0|q \$253385 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29056 \$253384 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29057 \$252822 s|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29058 VDD|pad|pin1|supply|vdd \$252821 d|z$56 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29059 s|zn$3 a1|zn$21 \$253901 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29060 \$253901 a2|zn$30 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29061 VDD|pad|pin1|supply|vdd a1|a3|i|i1|q a3|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29062 VDD|pad|pin1|supply|vdd a2|z$9 a3|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$29063 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q a3|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$29064 VDD|pad|pin1|supply|vdd RD[40]|a4|z a3|zn$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29065 \$253387 a1|zn$17 \$253388 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29066 VDD|pad|pin1|supply|vdd b|z \$253388 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$29067 VDD|pad|pin1|supply|vdd \$253388 d|z$57 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$29068 VDD|pad|pin1|supply|vdd a2|zn$31 \$253387 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29069 \$253390 a1|i0|q \$253486 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29070 \$253486 a2|i|s|zn \$253390 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.4565p AD=0.4565p PS=1.93u PD=1.93u
M$29071 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$253390 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29072 VDD|pad|pin1|supply|vdd \$253486 b|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29073 \$252823 \$252824 \$253391 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29074 \$253392 a2|i|s|zn \$252823 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29075 VDD|pad|pin1|supply|vdd a1|i0|q \$253392 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29076 \$253391 i0|i1|q$8 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29077 \$252824 a2|i|s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29078 VDD|pad|pin1|supply|vdd \$252823 i0|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29079 \$252825 \$252826 \$253394 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29080 \$253395 a1|a2|b|q|s \$252825 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29081 VDD|pad|pin1|supply|vdd i0|z \$253395 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29082 \$253394 i1|zn$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29083 \$252826 a1|a2|b|q|s VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29084 VDD|pad|pin1|supply|vdd \$252825 d|z$58 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29085 \$255088 \$254832 \$255087 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29086 \$255088 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29087 VDD|pad|pin1|supply|vdd R[46]|i0|q \$255090 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29088 \$255090 s|zn$3 \$255087 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29089 i|z$115 \$255097 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$29090 VDD|pad|pin1|supply|vdd CLK|core|i|p2c$1 \$255097
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p
+ PS=2.67u PD=2.23u
M$29091 \$255099 \$254835 \$255098 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29092 \$255099 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29093 VDD|pad|pin1|supply|vdd R[18]|i0|q \$255100 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29094 \$255100 s|zn$6 \$255098 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29095 \$255103 \$254836 \$255102 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29096 \$255103 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29097 VDD|pad|pin1|supply|vdd R[43]|i0|q \$255104 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29098 \$255104 s|zn$3 \$255102 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29099 \$255107 \$254837 \$255106 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29100 \$255107 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29101 VDD|pad|pin1|supply|vdd R[47]|i0|q \$255108 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29102 \$255108 s|zn$3 \$255106 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29103 s|zn$4 a1|zn$21 \$256980 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29104 \$256980 a2|zn$29 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29105 VDD|pad|pin1|supply|vdd a2|zn$27 a2|zn$31 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29106 a2|zn$31 a1|a2|b|q|s VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29107 a2|zn$31 a3|zn$8 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29108 VDD|pad|pin1|supply|vdd \$254828 \$256987 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29109 \$256987 d|z$50 \$255076 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29110 \$255076 \$255075 \$256922 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29111 \$256922 \$255077 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29112 VDD|pad|pin1|supply|vdd \$254830 \$256984 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29113 \$256984 d|z$59 \$255082 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29114 \$255082 \$255080 \$256923 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29115 \$256923 \$255083 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29116 VDD|pad|pin1|supply|vdd \$254833 \$256982 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29117 \$256982 d|z$60 \$255093 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29118 \$255093 \$255092 \$256924 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29119 \$256924 \$255094 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29120 VDD|pad|pin1|supply|vdd \$254839 \$256979 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29121 \$256979 d|z$57 \$255111 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29122 \$255111 \$255110 \$256925 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29123 \$256925 \$255112 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29124 VDD|pad|pin1|supply|vdd \$254841 \$256977 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29125 \$256977 d|z$58 \$255116 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29126 \$255116 \$255115 \$256926 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29127 \$256926 \$255117 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29128 \$255075 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29129 VDD|pad|pin1|supply|vdd \$255075 \$254828 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29130 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$256922
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29131 \$255077 \$255076 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29132 \$255077 \$255075 \$254829 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29133 \$254829 \$254828 \$256986 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29134 VDD|pad|pin1|supply|vdd \$255079 \$256986 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29135 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$255079
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29136 VDD|pad|pin1|supply|vdd \$254829 \$255079 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29137 VDD|pad|pin1|supply|vdd \$255079 R[42]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29138 \$255080 cp|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29139 VDD|pad|pin1|supply|vdd \$255080 \$254830 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29140 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$256923
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29141 \$255083 \$255082 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29142 \$255083 \$255080 \$254831 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29143 \$254831 \$254830 \$256983 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29144 VDD|pad|pin1|supply|vdd \$255085 \$256983 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29145 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$255085
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29146 VDD|pad|pin1|supply|vdd \$254831 \$255085 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29147 VDD|pad|pin1|supply|vdd \$255085 R[40]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29148 VDD|pad|pin1|supply|vdd s|zn$3 \$254832 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29149 VDD|pad|pin1|supply|vdd \$255087 d|z$60 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29150 \$255092 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29151 VDD|pad|pin1|supply|vdd \$255092 \$254833 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29152 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$256924
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29153 \$255094 \$255093 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29154 \$255094 \$255092 \$254834 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29155 \$254834 \$254833 \$256981 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29156 VDD|pad|pin1|supply|vdd \$255096 \$256981 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29157 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$255096
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29158 VDD|pad|pin1|supply|vdd \$254834 \$255096 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29159 VDD|pad|pin1|supply|vdd \$255096 R[46]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29160 VDD|pad|pin1|supply|vdd s|zn$6 \$254835 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29161 VDD|pad|pin1|supply|vdd \$255098 d|z$61 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29162 VDD|pad|pin1|supply|vdd s|zn$3 \$254836 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29163 VDD|pad|pin1|supply|vdd \$255102 d|z$62 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29164 VDD|pad|pin1|supply|vdd s|zn$3 \$254837 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29165 VDD|pad|pin1|supply|vdd \$255106 d|z$63 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29166 \$255110 cp|i|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29167 VDD|pad|pin1|supply|vdd \$255110 \$254839 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29168 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$256925
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29169 \$255112 \$255111 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29170 \$255112 \$255110 \$254840 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29171 \$254840 \$254839 \$256978 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29172 VDD|pad|pin1|supply|vdd \$255114 \$256978 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29173 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$255114
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29174 VDD|pad|pin1|supply|vdd \$254840 \$255114 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29175 VDD|pad|pin1|supply|vdd \$255114 a1|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29176 \$255115 cp|i|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29177 VDD|pad|pin1|supply|vdd \$255115 \$254841 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29178 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$256926
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29179 \$255117 \$255116 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29180 \$255117 \$255115 \$254842 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29181 \$254842 \$254841 \$256976 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29182 VDD|pad|pin1|supply|vdd \$255119 \$256976 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29183 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$255119
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29184 VDD|pad|pin1|supply|vdd \$254842 \$255119 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29185 VDD|pad|pin1|supply|vdd \$255119 i0|i1|q$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29186 VDD|pad|pin1|supply|vdd cp|z$4 \$256998 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29187 VDD|pad|pin1|supply|vdd \$256998 \$256999 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29188 VDD|pad|pin1|supply|vdd \$257748 \$257000 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29189 \$257747 \$256998 \$257000 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29190 VDD|pad|pin1|supply|vdd \$256999 \$257781 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29191 \$257781 d|z$66 \$257747 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29192 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$257000
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29193 \$257001 \$256999 \$257782 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29194 VDD|pad|pin1|supply|vdd \$258009 \$257782 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29195 VDD|pad|pin1|supply|vdd \$257747 \$257748 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29196 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$258009
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29197 VDD|pad|pin1|supply|vdd \$257001 \$258009 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29198 \$257748 \$256998 \$257001 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29199 VDD|pad|pin1|supply|vdd \$258009 i0|i1|q$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29200 \$257002 \$257003 \$257749 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29201 \$257750 s|zn$3 \$257002 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29202 VDD|pad|pin1|supply|vdd R[40]|i0|q \$257750 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29203 \$257749 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29204 \$257003 s|zn$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29205 VDD|pad|pin1|supply|vdd \$257002 d|z$59 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29206 VDD|pad|pin1|supply|vdd cp|i|z$4 \$257004 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29207 VDD|pad|pin1|supply|vdd \$257004 \$257005 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29208 VDD|pad|pin1|supply|vdd \$257752 \$257006 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29209 \$257751 \$257004 \$257006 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29210 VDD|pad|pin1|supply|vdd \$257005 \$257780 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29211 \$257780 d|z$52 \$257751 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29212 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$257006
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29213 \$257007 \$257005 \$257779 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29214 VDD|pad|pin1|supply|vdd \$258011 \$257779 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29215 VDD|pad|pin1|supply|vdd \$257751 \$257752 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29216 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$258011
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29217 VDD|pad|pin1|supply|vdd \$257007 \$258011 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29218 \$257752 \$257004 \$257007 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29219 VDD|pad|pin1|supply|vdd \$258011 R[44]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29220 \$257008 \$257009 \$257753 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29221 \$257754 s|zn$5 \$257008 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29222 VDD|pad|pin1|supply|vdd a2|i|i0|i1|q \$257754 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29223 \$257753 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29224 \$257009 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29225 VDD|pad|pin1|supply|vdd \$257008 d|z$64 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29226 VDD|pad|pin1|supply|vdd cp|i|z$4 \$257010 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29227 VDD|pad|pin1|supply|vdd \$257010 \$257011 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29228 VDD|pad|pin1|supply|vdd \$257757 \$257012 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29229 \$257756 \$257010 \$257012 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29230 VDD|pad|pin1|supply|vdd \$257011 \$257778 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29231 \$257778 d|z$64 \$257756 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29232 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$257012
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29233 \$257013 \$257011 \$257777 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29234 VDD|pad|pin1|supply|vdd \$258012 \$257777 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29235 VDD|pad|pin1|supply|vdd \$257756 \$257757 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29236 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$258012
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29237 VDD|pad|pin1|supply|vdd \$257013 \$258012 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29238 \$257757 \$257010 \$257013 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29239 VDD|pad|pin1|supply|vdd \$258012 a1|a3|i|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29240 VDD|pad|pin1|supply|vdd cp|i|z$5 \$257014 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29241 VDD|pad|pin1|supply|vdd \$257014 \$257015 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29242 VDD|pad|pin1|supply|vdd \$257759 \$257016 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29243 \$257758 \$257014 \$257016 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29244 VDD|pad|pin1|supply|vdd \$257015 \$257776 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29245 \$257776 d|z$61 \$257758 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29246 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$257016
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29247 \$257017 \$257015 \$257775 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29248 VDD|pad|pin1|supply|vdd \$258014 \$257775 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29249 VDD|pad|pin1|supply|vdd \$257758 \$257759 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29250 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$258014
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29251 VDD|pad|pin1|supply|vdd \$257017 \$258014 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29252 \$257759 \$257014 \$257017 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29253 VDD|pad|pin1|supply|vdd \$258014 R[18]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29254 VDD|pad|pin1|supply|vdd cp|i|z$6 \$257018 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29255 VDD|pad|pin1|supply|vdd \$257018 \$257019 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29256 VDD|pad|pin1|supply|vdd \$257761 \$257020 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29257 \$257760 \$257018 \$257020 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29258 VDD|pad|pin1|supply|vdd \$257019 \$257772 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29259 \$257772 d|z$62 \$257760 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29260 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$257020
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29261 \$257021 \$257019 \$257774 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29262 VDD|pad|pin1|supply|vdd \$258015 \$257774 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29263 VDD|pad|pin1|supply|vdd \$257760 \$257761 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29264 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$258015
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29265 VDD|pad|pin1|supply|vdd \$257021 \$258015 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29266 \$257761 \$257018 \$257021 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29267 VDD|pad|pin1|supply|vdd \$258015 R[43]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29268 VDD|pad|pin1|supply|vdd cp|i|z$1 \$257022 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29269 VDD|pad|pin1|supply|vdd \$257022 \$257023 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29270 VDD|pad|pin1|supply|vdd \$257763 \$257024 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29271 \$257762 \$257022 \$257024 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29272 VDD|pad|pin1|supply|vdd \$257023 \$257771 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29273 \$257771 d|z$63 \$257762 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29274 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$257024
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29275 \$257025 \$257023 \$257770 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29276 VDD|pad|pin1|supply|vdd \$258016 \$257770 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29277 VDD|pad|pin1|supply|vdd \$257762 \$257763 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29278 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$258016
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29279 VDD|pad|pin1|supply|vdd \$257025 \$258016 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29280 \$257763 \$257022 \$257025 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29281 VDD|pad|pin1|supply|vdd \$258016 R[47]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29282 \$257026 \$257027 \$257764 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29283 \$257765 a2|i|s|zn \$257026 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29284 VDD|pad|pin1|supply|vdd i0|i1|q$8 \$257765 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29285 \$257764 i0|i1|q$9 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29286 \$257027 a2|i|s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29287 VDD|pad|pin1|supply|vdd \$257026 i0|z$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29288 \$257028 \$257029 \$257767 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29289 \$257768 a1|a2|b|q|s \$257028 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29290 VDD|pad|pin1|supply|vdd i0|z$1 \$257768 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29291 \$257767 i1|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29292 \$257029 a1|a2|b|q|s VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29293 VDD|pad|pin1|supply|vdd \$257028 d|z$65 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29294 \$259368 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29295 VDD|pad|pin1|supply|vdd \$259368 \$259348 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29296 VDD|pad|pin1|supply|vdd \$259348 \$261174 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29297 \$261174 d|z$70 \$259369 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29298 \$259369 \$259368 \$261142 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29299 \$261142 \$259370 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29300 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$261142
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29301 \$259370 \$259369 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29302 \$259370 \$259368 \$259349 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29303 \$259349 \$259348 \$261170 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29304 VDD|pad|pin1|supply|vdd \$259372 \$261170 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29305 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$259372
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29306 VDD|pad|pin1|supply|vdd \$259349 \$259372 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29307 VDD|pad|pin1|supply|vdd \$259372 i0|i1|q$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29308 \$259374 \$259351 \$259373 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29309 \$259374 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29310 VDD|pad|pin1|supply|vdd i0|i1|q$5 \$259375 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29311 \$259375 s|zn$5 \$259373 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29312 VDD|pad|pin1|supply|vdd s|zn$5 \$259351 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29313 VDD|pad|pin1|supply|vdd \$259373 d|z$66 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29314 \$259377 \$259353 \$259376 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29315 \$259377 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29316 VDD|pad|pin1|supply|vdd R[16]|i0|q \$259378 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29317 \$259378 s|zn$6 \$259376 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29318 VDD|pad|pin1|supply|vdd s|zn$6 \$259353 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29319 VDD|pad|pin1|supply|vdd \$259376 d|z$67 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29320 \$259381 \$259354 \$259380 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29321 \$259381 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29322 VDD|pad|pin1|supply|vdd R[23]|i0|q \$259382 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29323 \$259382 s|zn$6 \$259380 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29324 VDD|pad|pin1|supply|vdd s|zn$6 \$259354 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29325 VDD|pad|pin1|supply|vdd \$259380 d|z$68 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29326 \$259384 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29327 VDD|pad|pin1|supply|vdd \$259384 \$259355 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29328 VDD|pad|pin1|supply|vdd \$259355 \$261167 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29329 \$261167 d|z$68 \$259385 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29330 \$259385 \$259384 \$261143 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29331 \$261143 \$259386 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29332 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$261143
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29333 \$259386 \$259385 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29334 \$259386 \$259384 \$259356 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29335 \$259356 \$259355 \$261168 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29336 VDD|pad|pin1|supply|vdd \$259388 \$261168 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29337 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$259388
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29338 VDD|pad|pin1|supply|vdd \$259356 \$259388 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29339 VDD|pad|pin1|supply|vdd \$259388 R[23]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29340 \$259389 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29341 VDD|pad|pin1|supply|vdd \$259389 \$259357 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29342 VDD|pad|pin1|supply|vdd \$259357 \$261166 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29343 \$261166 d|z$71 \$259390 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29344 \$259390 \$259389 \$261144 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29345 \$261144 \$259391 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29346 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$261144
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29347 \$259391 \$259390 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29348 \$259391 \$259389 \$259358 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29349 \$259358 \$259357 \$261162 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29350 VDD|pad|pin1|supply|vdd \$259393 \$261162 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29351 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$259393
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29352 VDD|pad|pin1|supply|vdd \$259358 \$259393 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29353 VDD|pad|pin1|supply|vdd \$259393 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29354 \$259394 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29355 VDD|pad|pin1|supply|vdd \$259394 \$259359 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29356 VDD|pad|pin1|supply|vdd \$259359 \$261160 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29357 \$261160 d|z$72 \$259395 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29358 \$259395 \$259394 \$261145 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29359 \$261145 \$259396 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29360 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$261145
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29361 \$259396 \$259395 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29362 \$259396 \$259394 \$259360 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29363 \$259360 \$259359 \$261161 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29364 VDD|pad|pin1|supply|vdd \$259398 \$261161 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29365 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$259398
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29366 VDD|pad|pin1|supply|vdd \$259360 \$259398 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29367 VDD|pad|pin1|supply|vdd \$259398 R[21]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29368 s|zn$6 a1|zn$21 \$261157 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29369 \$261157 a2|zn$28 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29370 \$259399 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29371 VDD|pad|pin1|supply|vdd \$259399 \$259361 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29372 VDD|pad|pin1|supply|vdd \$259361 \$261159 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29373 \$261159 d|z$73 \$259400 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29374 \$259400 \$259399 \$261146 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29375 \$261146 \$259401 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29376 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$261146
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29377 \$259401 \$259400 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29378 \$259401 \$259399 \$259362 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29379 \$259362 \$259361 \$261152 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29380 VDD|pad|pin1|supply|vdd \$259403 \$261152 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29381 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$259403
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29382 VDD|pad|pin1|supply|vdd \$259362 \$259403 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29383 VDD|pad|pin1|supply|vdd \$259403 R[22]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29384 \$259405 \$259363 \$259404 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29385 \$259405 i1|z$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29386 VDD|pad|pin1|supply|vdd i0|z$2 \$259406 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29387 \$259406 a1|a2|b|q|s \$259404 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29388 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$259363 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29389 VDD|pad|pin1|supply|vdd \$259404 d|z$69 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29390 \$259408 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29391 VDD|pad|pin1|supply|vdd \$259408 \$259364 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29392 VDD|pad|pin1|supply|vdd \$259364 \$261149 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29393 \$261149 d|z$65 \$259409 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29394 \$259409 \$259408 \$261147 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29395 \$261147 \$259410 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29396 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$261147
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29397 \$259410 \$259409 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29398 \$259410 \$259408 \$259365 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29399 \$259365 \$259364 \$261148 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29400 VDD|pad|pin1|supply|vdd \$259412 \$261148 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29401 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$259412
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29402 VDD|pad|pin1|supply|vdd \$259365 \$259412 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29403 VDD|pad|pin1|supply|vdd \$259412 i0|i1|q$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29404 CLK|core|i|p2c$1 \$258894 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$29405 \$261262 \$261217 \$261263 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29406 \$261264 s|zn$5 \$261262 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29407 VDD|pad|pin1|supply|vdd i0|i1|q$3 \$261264 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29408 \$261263 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29409 \$261217 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29410 VDD|pad|pin1|supply|vdd \$261262 d|z$70 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29411 \$261265 \$261218 \$261266 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29412 \$261267 s|zn$5 \$261265 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29413 VDD|pad|pin1|supply|vdd i0|i1|q$7 \$261267 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29414 \$261266 i0|i1|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29415 \$261218 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29416 VDD|pad|pin1|supply|vdd \$261265 d|z$74 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29417 VDD|pad|pin1|supply|vdd cp|i|z$7 \$261269 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29418 VDD|pad|pin1|supply|vdd \$261269 \$261270 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29419 VDD|pad|pin1|supply|vdd \$261847 \$261272 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29420 \$261271 \$261269 \$261272 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29421 VDD|pad|pin1|supply|vdd \$261270 \$262077 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29422 \$262077 d|z$74 \$261271 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29423 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$261272
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29424 \$261273 \$261270 \$261844 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29425 VDD|pad|pin1|supply|vdd \$262081 \$261844 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29426 VDD|pad|pin1|supply|vdd \$261271 \$261847 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29427 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$262081
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29428 VDD|pad|pin1|supply|vdd \$261273 \$262081 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29429 \$261847 \$261269 \$261273 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29430 VDD|pad|pin1|supply|vdd \$262081 i0|i1|q$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29431 VDD|pad|pin1|supply|vdd cp|i|z$4 \$261274 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29432 VDD|pad|pin1|supply|vdd \$261274 \$261275 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29433 VDD|pad|pin1|supply|vdd \$261848 \$261277 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29434 \$261276 \$261274 \$261277 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29435 VDD|pad|pin1|supply|vdd \$261275 \$262080 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29436 \$262080 d|z$78 \$261276 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29437 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$261277
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29438 \$261278 \$261275 \$261839 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29439 VDD|pad|pin1|supply|vdd \$262082 \$261839 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29440 VDD|pad|pin1|supply|vdd \$261276 \$261848 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29441 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$262082
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29442 VDD|pad|pin1|supply|vdd \$261278 \$262082 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29443 \$261848 \$261274 \$261278 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29444 VDD|pad|pin1|supply|vdd \$262082 a1|i|i0|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29445 \$261279 \$261219 \$261280 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29446 \$261281 s|zn$5 \$261279 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29447 VDD|pad|pin1|supply|vdd a1|i|i0|i1|q \$261281 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29448 \$261280 a2|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29449 \$261219 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29450 VDD|pad|pin1|supply|vdd \$261279 d|z$71 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29451 \$261282 \$261220 \$261283 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29452 \$261284 s|zn$6 \$261282 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29453 VDD|pad|pin1|supply|vdd R[21]|i0|q \$261284 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29454 \$261283 i0|i1|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29455 \$261220 s|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29456 VDD|pad|pin1|supply|vdd \$261282 d|z$72 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29457 \$261285 \$261221 \$261286 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29458 \$261287 s|zn$6 \$261285 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29459 VDD|pad|pin1|supply|vdd R[20]|i0|q \$261287 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29460 \$261286 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29461 \$261221 s|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29462 VDD|pad|pin1|supply|vdd \$261285 d|z$75 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29463 \$261289 \$261222 \$261290 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29464 \$261291 s|zn$6 \$261289 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29465 VDD|pad|pin1|supply|vdd R[19]|i0|q \$261291 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29466 \$261290 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29467 \$261222 s|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29468 VDD|pad|pin1|supply|vdd \$261289 d|z$76 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29469 \$261293 \$261223 \$261294 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29470 \$261295 s|zn$6 \$261293 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29471 VDD|pad|pin1|supply|vdd R[22]|i0|q \$261295 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29472 \$261294 i0|i1|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29473 \$261223 s|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29474 VDD|pad|pin1|supply|vdd \$261293 d|z$73 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29475 \$261296 \$261224 \$261297 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29476 \$261298 a1|a2|b|q|s \$261296 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29477 VDD|pad|pin1|supply|vdd i0|z$3 \$261298 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29478 \$261297 i1|z$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29479 \$261224 a1|a2|b|q|s VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29480 VDD|pad|pin1|supply|vdd \$261296 d|z$77 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29481 VDD|pad|pin1|supply|vdd cp|i|z$6 \$261300 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29482 VDD|pad|pin1|supply|vdd \$261300 \$261301 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29483 VDD|pad|pin1|supply|vdd \$261851 \$261303 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29484 \$261302 \$261300 \$261303 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29485 VDD|pad|pin1|supply|vdd \$261301 \$262079 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29486 \$262079 d|z$69 \$261302 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29487 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$261303
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29488 \$261304 \$261301 \$261768 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29489 VDD|pad|pin1|supply|vdd \$262083 \$261768 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29490 VDD|pad|pin1|supply|vdd \$261302 \$261851 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29491 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$262083
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29492 VDD|pad|pin1|supply|vdd \$261304 \$262083 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29493 \$261851 \$261300 \$261304 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29494 VDD|pad|pin1|supply|vdd \$262083 i0|i1|q$10 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29495 \$263506 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29496 VDD|pad|pin1|supply|vdd \$263506 \$263439 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29497 VDD|pad|pin1|supply|vdd \$263439 \$265332 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29498 \$265332 d|z$81 \$263507 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29499 \$263507 \$263506 \$264486 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29500 \$264486 \$263508 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29501 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$264486
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29502 \$263508 \$263507 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29503 \$263508 \$263506 \$263440 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29504 \$263440 \$263439 \$265328 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29505 VDD|pad|pin1|supply|vdd \$263510 \$265328 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29506 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$263510
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29507 VDD|pad|pin1|supply|vdd \$263440 \$263510 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29508 VDD|pad|pin1|supply|vdd \$263510 i0|i1|q$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29509 \$263511 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29510 VDD|pad|pin1|supply|vdd \$263511 \$263441 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29511 VDD|pad|pin1|supply|vdd \$263441 \$265329 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29512 \$265329 d|z$67 \$263512 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29513 \$263512 \$263511 \$264487 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29514 \$264487 \$263513 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29515 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$264487
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29516 \$263513 \$263512 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29517 \$263513 \$263511 \$263442 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29518 \$263442 \$263441 \$265327 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29519 VDD|pad|pin1|supply|vdd \$263515 \$265327 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29520 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$263515
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29521 VDD|pad|pin1|supply|vdd \$263442 \$263515 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29522 VDD|pad|pin1|supply|vdd \$263515 R[16]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29523 \$263517 \$263443 \$263516 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29524 \$263517 a1|i|i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29525 VDD|pad|pin1|supply|vdd i0|i1|q$4 \$263518 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29526 \$263518 s|zn$5 \$263516 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29527 VDD|pad|pin1|supply|vdd s|zn$5 \$263443 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29528 VDD|pad|pin1|supply|vdd \$263516 d|z$78 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29529 \$263520 \$263444 \$263519 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29530 \$263520 i1|zn$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29531 VDD|pad|pin1|supply|vdd i0|z$4 \$263521 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29532 \$263521 a1|a2|b|q|s \$263519 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29533 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$263444 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29534 VDD|pad|pin1|supply|vdd \$263519 d|z$79 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29535 \$263524 \$263445 \$263523 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29536 \$263524 i1|z$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29537 VDD|pad|pin1|supply|vdd i0|z$5 \$263525 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29538 \$263525 a1|a2|b|q|s \$263523 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29539 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$263445 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29540 VDD|pad|pin1|supply|vdd \$263523 d|z$80 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29541 \$263528 \$263446 \$263527 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29542 \$263528 i0|i1|q$11 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29543 VDD|pad|pin1|supply|vdd i0|i1|q$12 \$263529 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29544 \$263529 a2|i|s|zn \$263527 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29545 VDD|pad|pin1|supply|vdd a2|i|s|zn \$263446 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29546 VDD|pad|pin1|supply|vdd \$263527 i0|z$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29547 \$263530 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29548 VDD|pad|pin1|supply|vdd \$263530 \$263447 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29549 VDD|pad|pin1|supply|vdd \$263447 \$265325 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29550 \$265325 d|z$75 \$263531 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29551 \$263531 \$263530 \$264488 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29552 \$264488 \$263532 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29553 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$264488
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29554 \$263532 \$263531 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29555 \$263532 \$263530 \$263448 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29556 \$263448 \$263447 \$265326 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29557 VDD|pad|pin1|supply|vdd \$263534 \$265326 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29558 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$263534
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29559 VDD|pad|pin1|supply|vdd \$263448 \$263534 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29560 VDD|pad|pin1|supply|vdd \$263534 R[20]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29561 \$263535 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29562 VDD|pad|pin1|supply|vdd \$263535 \$263449 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29563 VDD|pad|pin1|supply|vdd \$263449 \$265323 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29564 \$265323 d|z$76 \$263536 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29565 \$263536 \$263535 \$264489 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29566 \$264489 \$263537 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29567 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$264489
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29568 \$263537 \$263536 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29569 \$263537 \$263535 \$263450 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29570 \$263450 \$263449 \$265324 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29571 VDD|pad|pin1|supply|vdd \$263539 \$265324 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29572 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$263539
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29573 VDD|pad|pin1|supply|vdd \$263450 \$263539 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29574 VDD|pad|pin1|supply|vdd \$263539 R[19]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29575 \$263540 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29576 VDD|pad|pin1|supply|vdd \$263540 \$263451 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29577 VDD|pad|pin1|supply|vdd \$263451 \$265321 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29578 \$265321 d|z$77 \$263541 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29579 \$263541 \$263540 \$264490 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29580 \$264490 \$263542 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29581 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$264490
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29582 \$263542 \$263541 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29583 \$263542 \$263540 \$263452 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29584 \$263452 \$263451 \$265322 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29585 VDD|pad|pin1|supply|vdd \$263544 \$265322 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29586 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$263544
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29587 VDD|pad|pin1|supply|vdd \$263452 \$263544 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29588 VDD|pad|pin1|supply|vdd \$263544 i0|i1|q$12 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29589 \$263546 \$263453 \$263545 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29590 \$263546 i0|i1|q$10 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29591 VDD|pad|pin1|supply|vdd i0|i1|q$9 \$263547 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29592 \$263547 a2|i|s|zn \$263545 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29593 VDD|pad|pin1|supply|vdd a2|i|s|zn \$263453 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29594 VDD|pad|pin1|supply|vdd \$263545 i0|z$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29595 VDD|pad|pin1|supply|vdd cp|i|z$7 \$265338 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29596 VDD|pad|pin1|supply|vdd \$265338 \$265339 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29597 VDD|pad|pin1|supply|vdd \$266387 \$265340 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29598 \$265479 \$265338 \$265340 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29599 VDD|pad|pin1|supply|vdd \$265339 \$266262 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29600 \$266262 d|z$83 \$265479 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29601 \$267881 \$267883 \$267880 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29602 \$267881 i0|i1|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29603 VDD|pad|pin1|supply|vdd i0|i1|q$2 \$267882 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29604 \$267882 s|zn$5 \$267880 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29605 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$265340
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29606 \$265341 \$265339 \$266273 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29607 VDD|pad|pin1|supply|vdd \$266428 \$266273 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29608 VDD|pad|pin1|supply|vdd \$265479 \$266387 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29609 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$266428
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29610 VDD|pad|pin1|supply|vdd \$265341 \$266428 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29611 \$266387 \$265338 \$265341 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29612 VDD|pad|pin1|supply|vdd \$266428 i0|i1|q$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29613 \$267885 \$267887 \$267884 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29614 \$267885 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29615 VDD|pad|pin1|supply|vdd i0|i1|q \$267886 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29616 \$267886 s|zn$5 \$267884 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29617 VDD|pad|pin1|supply|vdd cp|i|z$7 \$265342 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29618 VDD|pad|pin1|supply|vdd \$265342 \$265343 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29619 VDD|pad|pin1|supply|vdd \$266388 \$265344 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29620 \$265480 \$265342 \$265344 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29621 VDD|pad|pin1|supply|vdd \$265343 \$266280 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29622 \$266280 d|z$84 \$265480 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29623 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$265344
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29624 \$265345 \$265343 \$266275 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29625 VDD|pad|pin1|supply|vdd \$266429 \$266275 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29626 VDD|pad|pin1|supply|vdd \$265480 \$266388 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29627 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$266429
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29628 VDD|pad|pin1|supply|vdd \$265345 \$266429 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29629 \$266388 \$265342 \$265345 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29630 VDD|pad|pin1|supply|vdd \$266429 i0|i1|q$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29631 VDD|pad|pin1|supply|vdd cp|i|z$7 \$265346 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29632 VDD|pad|pin1|supply|vdd \$265346 \$265347 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29633 VDD|pad|pin1|supply|vdd \$266389 \$265348 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29634 \$265481 \$265346 \$265348 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29635 VDD|pad|pin1|supply|vdd \$265347 \$266282 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29636 \$266282 d|z$85 \$265481 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29637 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$265348
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29638 \$265349 \$265347 \$266285 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29639 VDD|pad|pin1|supply|vdd \$266430 \$266285 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29640 VDD|pad|pin1|supply|vdd \$265481 \$266389 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29641 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$266430
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29642 VDD|pad|pin1|supply|vdd \$265349 \$266430 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29643 \$266389 \$265346 \$265349 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29644 VDD|pad|pin1|supply|vdd \$266430 R[17]|i0|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29645 VDD|pad|pin1|supply|vdd cp|i|z$4 \$265350 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29646 VDD|pad|pin1|supply|vdd \$265350 \$265351 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29647 VDD|pad|pin1|supply|vdd \$266390 \$265352 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29648 \$265482 \$265350 \$265352 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29649 VDD|pad|pin1|supply|vdd \$265351 \$266289 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29650 \$266289 d|z$79 \$265482 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29651 z$32 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29652 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$265352
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29653 \$265353 \$265351 \$266296 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29654 VDD|pad|pin1|supply|vdd \$266431 \$266296 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29655 VDD|pad|pin1|supply|vdd \$265482 \$266390 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29656 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$266431
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29657 VDD|pad|pin1|supply|vdd \$265353 \$266431 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29658 \$266390 \$265350 \$265353 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29659 VDD|pad|pin1|supply|vdd \$266431 i0|i1|q$13 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29660 VDD|pad|pin1|supply|vdd a1|b|d|z s|zn$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29661 s|zn$5 a1|zn$22 \$269781 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.4565p AD=0.4565p PS=1.93u PD=1.93u
M$29662 \$269781 a2|zn$32 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29663 \$267906 \$267908 \$267905 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29664 \$267906 a1|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29665 VDD|pad|pin1|supply|vdd i0|i1|q$13 \$267907 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29666 \$267907 a2|i|s|zn \$267905 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29667 VDD|pad|pin1|supply|vdd cp|i|z$4 \$265354 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29668 VDD|pad|pin1|supply|vdd \$265354 \$265355 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29669 VDD|pad|pin1|supply|vdd \$266391 \$265356 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29670 \$265484 \$265354 \$265356 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29671 VDD|pad|pin1|supply|vdd \$265355 \$266300 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29672 \$266300 d|z$80 \$265484 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29673 \$267911 \$267913 \$267910 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29674 \$267911 i0|i1|q$13 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29675 VDD|pad|pin1|supply|vdd i0|i1|q$11 \$267912 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29676 \$267912 a2|i|s|zn \$267910 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29677 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$265356
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29678 \$265357 \$265355 \$266307 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29679 VDD|pad|pin1|supply|vdd \$266432 \$266307 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29680 VDD|pad|pin1|supply|vdd \$265484 \$266391 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29681 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$266432
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29682 VDD|pad|pin1|supply|vdd \$265357 \$266432 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29683 \$266391 \$265354 \$265357 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29684 VDD|pad|pin1|supply|vdd \$266432 i0|i1|q$11 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29685 VDD|pad|pin1|supply|vdd a2|q \$267914 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29686 \$267914 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29687 DOUT_EN|z \$267914 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29688 cp|i|z$4 \$267916 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.494625p PS=3.33u PD=2.67u
M$29689 VDD|pad|pin1|supply|vdd i|z$115 \$267916 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$29690 VDD|pad|pin1|supply|vdd a1|a2|q$2 a1|zn$21 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29691 a1|zn$21 a1|i0|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29692 \$267919 \$267921 \$267917 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29693 \$267919 DATA|core|i0|i1|p2c VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p
+ PS=1.93u PD=1.93u
M$29694 VDD|pad|pin1|supply|vdd a1|i0|q$1 \$267920 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29695 \$267920 d|s|zn \$267917 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29696 VDD|pad|pin1|supply|vdd a1|a2|q$2 \$267923 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29697 \$267923 a1|i0|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29698 a1|a2|a4|z \$267923 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$29699 \$265358 \$265359 \$265485 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29700 \$265486 a2|i|s|zn \$265358 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29701 VDD|pad|pin1|supply|vdd i0|i1|q$10 \$265486 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29702 \$265485 i0|i1|q$12 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29703 \$265359 a2|i|s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29704 VDD|pad|pin1|supply|vdd \$265358 i0|z$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29705 a1|b|d|z CEB|a1|core|i|p2c VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p
+ PS=3.33u PD=3.33u
M$29706 z$31 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29707 VDD|pad|pin1|supply|vdd a1|a2|q \$265488 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29708 VDD|pad|pin1|supply|vdd a1|b|d|z \$265488 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29709 VDD|pad|pin1|supply|vdd \$265488 d|z$82 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29710 VDD|pad|pin1|supply|vdd s|zn$5 \$267883 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29711 VDD|pad|pin1|supply|vdd \$267880 d|z$81 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29712 VDD|pad|pin1|supply|vdd s|zn$5 \$267887 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29713 VDD|pad|pin1|supply|vdd \$267884 d|z$86 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29714 VDD|pad|pin1|supply|vdd \$267890 \$269865 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29715 \$269865 d|z$86 \$267891 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29716 \$267891 \$267889 \$269389 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29717 \$269389 \$267892 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29718 VDD|pad|pin1|supply|vdd \$267897 \$269847 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29719 \$269847 d|z$88 \$267898 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29720 \$267898 \$267896 \$269390 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29721 \$269390 \$267899 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29722 VDD|pad|pin1|supply|vdd a2|i|s|zn \$267908 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29723 VDD|pad|pin1|supply|vdd \$267905 i0|z$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29724 VDD|pad|pin1|supply|vdd a2|i|s|zn \$267913 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29725 VDD|pad|pin1|supply|vdd \$267910 i0|z$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29726 VDD|pad|pin1|supply|vdd d|s|zn \$267921 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29727 VDD|pad|pin1|supply|vdd \$267917 d|z$87 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29728 VDD|pad|pin1|supply|vdd \$267925 \$269726 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29729 \$269726 a1|b|d|z \$267926 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29730 \$267926 \$267924 \$269391 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29731 \$269391 \$267927 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29732 VDD|pad|pin1|supply|vdd \$267933 \$269657 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29733 \$269657 d|z$82 \$267934 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29734 \$267934 \$267932 \$269392 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29735 \$269392 \$267935 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29736 \$269998 \$269910 \$270063 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29737 \$270064 s|zn$5 \$269998 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29738 VDD|pad|pin1|supply|vdd i0|i1|q$1 \$270064 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29739 \$270063 i0|i1|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29740 \$269910 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29741 VDD|pad|pin1|supply|vdd \$269998 d|z$83 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29742 \$269999 \$269911 \$270065 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29743 \$270066 s|zn$5 \$269999 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29744 VDD|pad|pin1|supply|vdd i0|i1|q$6 \$270066 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29745 \$270065 i0|i1|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29746 \$269911 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29747 VDD|pad|pin1|supply|vdd \$269999 d|z$84 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29748 \$267889 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29749 VDD|pad|pin1|supply|vdd \$267889 \$267890 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29750 z$33 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29751 VDD|pad|pin1|supply|vdd i|z$115 \$270000 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$29752 VDD|pad|pin1|supply|vdd \$270000 cp|i|z$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$29753 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$269389
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29754 \$267892 \$267891 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29755 \$267892 \$267889 \$267893 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29756 \$267893 \$267890 \$269824 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29757 VDD|pad|pin1|supply|vdd \$267895 \$269824 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29758 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$267895
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29759 VDD|pad|pin1|supply|vdd \$267893 \$267895 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29760 VDD|pad|pin1|supply|vdd \$267895 i0|i1|q$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29761 \$270001 \$269912 \$270068 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29762 \$270069 s|zn$5 \$270001 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29763 VDD|pad|pin1|supply|vdd DATA|core|i0|i1|p2c \$270069
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p
+ PS=1.93u PD=1.74u
M$29764 \$270068 i0|i1|q VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29765 \$269912 s|zn$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29766 VDD|pad|pin1|supply|vdd \$270001 d|z$88 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29767 \$270002 \$269913 \$270070 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29768 \$270071 s|zn$6 \$270002 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29769 VDD|pad|pin1|supply|vdd R[17]|i0|q \$270071 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29770 \$270070 i0|i1|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29771 \$267896 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29772 VDD|pad|pin1|supply|vdd \$267896 \$267897 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29773 \$269913 s|zn$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29774 VDD|pad|pin1|supply|vdd \$270002 d|z$85 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29775 VDD|pad|pin1|supply|vdd cp|i|z$4 \$270003 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29776 VDD|pad|pin1|supply|vdd \$270003 \$270004 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29777 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$269390
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29778 \$267899 \$267898 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29779 \$267899 \$267896 \$267900 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29780 \$267900 \$267897 \$269813 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29781 VDD|pad|pin1|supply|vdd \$267902 \$269813 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29782 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$267902
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29783 VDD|pad|pin1|supply|vdd \$267900 \$267902 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29784 VDD|pad|pin1|supply|vdd \$267902 i0|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29785 VDD|pad|pin1|supply|vdd \$270779 \$270005 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29786 \$270072 \$270003 \$270005 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29787 VDD|pad|pin1|supply|vdd \$270004 \$270744 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29788 \$270744 d|z$90 \$270072 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29789 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$270005
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29790 \$270006 \$270004 \$270059 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29791 VDD|pad|pin1|supply|vdd \$270780 \$270059 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29792 VDD|pad|pin1|supply|vdd \$270072 \$270779 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29793 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$270780
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29794 VDD|pad|pin1|supply|vdd \$270006 \$270780 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29795 \$270779 \$270003 \$270006 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29796 VDD|pad|pin1|supply|vdd \$270780 a1|i1|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29797 VDD|pad|pin1|supply|vdd cp|i|z$4 \$270007 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29798 VDD|pad|pin1|supply|vdd \$270007 \$270008 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29799 VDD|pad|pin1|supply|vdd \$270781 \$270009 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29800 \$270074 \$270007 \$270009 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29801 VDD|pad|pin1|supply|vdd \$270008 \$270749 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29802 \$270749 d|z$91 \$270074 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29803 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$270009
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29804 \$270010 \$270008 \$270058 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29805 VDD|pad|pin1|supply|vdd \$270782 \$270058 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29806 VDD|pad|pin1|supply|vdd \$270074 \$270781 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29807 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$270782
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29808 VDD|pad|pin1|supply|vdd \$270010 \$270782 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29809 \$270781 \$270007 \$270010 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29810 VDD|pad|pin1|supply|vdd \$270782 DOUT_DAT|c2p|core|i|q
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p
+ PS=2.67u PD=3.33u
M$29811 VDD|pad|pin1|supply|vdd cp|i|z$5 \$270011 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29812 VDD|pad|pin1|supply|vdd \$270011 \$270012 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29813 VDD|pad|pin1|supply|vdd \$270783 \$270013 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29814 \$270075 \$270011 \$270013 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29815 VDD|pad|pin1|supply|vdd \$270012 \$270771 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29816 \$270771 d|z$87 \$270075 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29817 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$270013
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29818 \$270014 \$270012 \$270057 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29819 VDD|pad|pin1|supply|vdd \$270784 \$270057 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29820 VDD|pad|pin1|supply|vdd \$270075 \$270783 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29821 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$270784
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29822 VDD|pad|pin1|supply|vdd \$270014 \$270784 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29823 \$270783 \$270011 \$270014 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29824 VDD|pad|pin1|supply|vdd \$270784 a1|i0|q$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29825 VDD|pad|pin1|supply|vdd cp|i|z$5 \$270015 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29826 VDD|pad|pin1|supply|vdd \$270015 \$270016 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29827 VDD|pad|pin1|supply|vdd \$270785 \$270017 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29828 \$270076 \$270015 \$270017 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29829 VDD|pad|pin1|supply|vdd \$270016 \$270774 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29830 \$270774 d|s|zn \$270076 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29831 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$270017
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29832 \$270787 \$270016 \$270056 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29833 VDD|pad|pin1|supply|vdd \$270786 \$270056 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29834 VDD|pad|pin1|supply|vdd \$270076 \$270785 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29835 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$270786
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29836 VDD|pad|pin1|supply|vdd \$270787 \$270786 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29837 \$270785 \$270015 \$270787 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29838 VDD|pad|pin1|supply|vdd \$270786 a2|i|q$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29839 \$267924 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29840 VDD|pad|pin1|supply|vdd \$267924 \$267925 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29841 a2|z$13 a2|i|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29842 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$269391
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29843 \$267927 \$267926 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29844 \$267927 \$267924 \$267928 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29845 \$267928 \$267925 \$269690 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29846 VDD|pad|pin1|supply|vdd \$267930 \$269690 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29847 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$267930
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29848 VDD|pad|pin1|supply|vdd \$267928 \$267930 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29849 VDD|pad|pin1|supply|vdd \$267930 a1|a2|q$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29850 VDD|pad|pin1|supply|vdd a2|q$1 \$270079 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29851 VDD|pad|pin1|supply|vdd a1|b|d|z \$270079 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29852 VDD|pad|pin1|supply|vdd \$270079 d|z$89 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29853 VDD|pad|pin1|supply|vdd a3|zn$10 a1|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29854 VDD|pad|pin1|supply|vdd a2|z$13 a1|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$29855 VDD|pad|pin1|supply|vdd a1|a2|q$1 a1|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$29856 VDD|pad|pin1|supply|vdd a4|zn$6 a1|zn$22 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29857 VDD|pad|pin1|supply|vdd i|z$115 \$270018 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$29858 VDD|pad|pin1|supply|vdd \$270018 cp|i|z$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$29859 \$267932 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29860 VDD|pad|pin1|supply|vdd \$267932 \$267933 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29861 VDD|pad|pin1|supply|vdd cp|i|z$6 \$270019 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29862 VDD|pad|pin1|supply|vdd \$270019 \$270020 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29863 VDD|pad|pin1|supply|vdd \$270788 \$270021 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29864 \$270081 \$270019 \$270021 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29865 VDD|pad|pin1|supply|vdd \$270020 \$270763 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29866 \$270763 d|z$89 \$270081 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29867 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$269392
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29868 \$267935 \$267934 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29869 \$267935 \$267932 \$267936 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29870 \$267936 \$267933 \$269679 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29871 VDD|pad|pin1|supply|vdd \$267938 \$269679 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29872 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$267938
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29873 VDD|pad|pin1|supply|vdd \$267936 \$267938 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29874 VDD|pad|pin1|supply|vdd \$267938 a1|a2|b|q|s VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29875 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$270021
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29876 \$270022 \$270020 \$270055 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29877 VDD|pad|pin1|supply|vdd \$270789 \$270055 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29878 VDD|pad|pin1|supply|vdd \$270081 \$270788 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29879 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$270789
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29880 VDD|pad|pin1|supply|vdd \$270022 \$270789 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29881 \$270788 \$270019 \$270022 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29882 VDD|pad|pin1|supply|vdd \$270789 a1|a2|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29883 VDD|pad|pin1|supply|vdd cp|i|z$7 \$274510 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29884 VDD|pad|pin1|supply|vdd \$274510 \$274511 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29885 \$272012 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29886 VDD|pad|pin1|supply|vdd \$272012 \$272013 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29887 VDD|pad|pin1|supply|vdd \$274520 \$274512 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$29888 \$274519 \$274510 \$274512 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29889 VDD|pad|pin1|supply|vdd \$274511 \$275183 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29890 \$275183 d|z$98 \$274519 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29891 VDD|pad|pin1|supply|vdd \$272013 \$274053 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29892 \$274053 d|z$92 \$272014 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29893 \$272014 \$272012 \$273661 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29894 \$273661 \$272015 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29895 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$274512
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29896 \$274513 \$274511 \$275179 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29897 VDD|pad|pin1|supply|vdd \$275260 \$275179 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29898 VDD|pad|pin1|supply|vdd \$274519 \$274520 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$29899 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$275260
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29900 VDD|pad|pin1|supply|vdd \$274513 \$275260 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29901 \$274520 \$274510 \$274513 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29902 VDD|pad|pin1|supply|vdd \$275260 a2|q$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29903 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$273661
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29904 \$272015 \$272014 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29905 \$272015 \$272012 \$272016 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29906 \$272016 \$272013 \$274057 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29907 VDD|pad|pin1|supply|vdd \$272018 \$274057 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29908 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$272018
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29909 VDD|pad|pin1|supply|vdd \$272016 \$272018 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29910 VDD|pad|pin1|supply|vdd \$272018 a1|a2|q$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29911 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$274521 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29912 VDD|pad|pin1|supply|vdd a1|b|d|z \$274521 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29913 a3|zn$9 a1|a2|q$3 \$274054 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29914 \$274054 a2|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$29915 VDD|pad|pin1|supply|vdd \$274521 d|z$92 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29916 VDD|pad|pin1|supply|vdd a1|a2|q$3 \$274522 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29917 VDD|pad|pin1|supply|vdd a1|b|d|z \$274522 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29918 \$272022 \$272024 \$272021 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.383625p AD=0.31075p PS=1.93u PD=2.23u
M$29919 \$272022 i1|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p PS=1.93u PD=1.93u
M$29920 VDD|pad|pin1|supply|vdd i0|z$6 \$272023 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29921 \$272023 a1|a2|b|q|s \$272021 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29922 VDD|pad|pin1|supply|vdd \$274522 d|z$98 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29923 VDD|pad|pin1|supply|vdd a1|a2|b|q|s \$272024 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.2904p AD=0.31075p PS=1.6u PD=2.23u
M$29924 VDD|pad|pin1|supply|vdd \$272021 d|z$90 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29925 VDD|pad|pin1|supply|vdd a1|a2|q$5 \$274523 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29926 VDD|pad|pin1|supply|vdd a1|b|d|z \$274523 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29927 VDD|pad|pin1|supply|vdd \$274523 d|z$95 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29928 \$272025 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29929 VDD|pad|pin1|supply|vdd \$272025 \$272026 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29930 a1|z$17 a2|i|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29931 VDD|pad|pin1|supply|vdd \$272026 \$274063 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29932 \$274063 a2|d|z \$272027 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29933 \$272027 \$272025 \$273662 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29934 \$273662 \$272028 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29935 VDD|pad|pin1|supply|vdd a2|d|z \$274526 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29936 VDD|pad|pin1|supply|vdd a1|i1|q \$274526 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29937 VDD|pad|pin1|supply|vdd \$274526 d|z$91 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29938 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$273662
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29939 \$272028 \$272027 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29940 \$272028 \$272025 \$272029 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29941 \$272029 \$272026 \$274071 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29942 VDD|pad|pin1|supply|vdd \$272031 \$274071 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29943 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$272031
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29944 VDD|pad|pin1|supply|vdd \$272029 \$272031 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29945 VDD|pad|pin1|supply|vdd \$272031 a2|q VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29946 a2|d|z a2|i|s|zn VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29947 VDD|pad|pin1|supply|vdd a2|i|q$2 \$274527 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29948 VDD|pad|pin1|supply|vdd a1|b|d|z \$274527 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29949 VDD|pad|pin1|supply|vdd \$274527 d|z$96 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29950 VDD|pad|pin1|supply|vdd a1|a2|q$2 \$274529 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29951 VDD|pad|pin1|supply|vdd a1|b|d|z \$274529 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29952 z$34 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.6215p PS=3.33u PD=3.33u
M$29953 VDD|pad|pin1|supply|vdd \$274529 d|z$97 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29954 \$272033 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29955 VDD|pad|pin1|supply|vdd \$272033 \$272034 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29956 VDD|pad|pin1|supply|vdd \$272034 \$274075 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29957 \$274075 d|z$93 \$272035 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29958 \$272035 \$272033 \$273663 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29959 \$273663 \$272036 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29960 VDD|pad|pin1|supply|vdd i|z$115 \$274531 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.494625p AD=0.31075p PS=2.67u PD=2.23u
M$29961 VDD|pad|pin1|supply|vdd \$274531 cp|i|z$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.494625p AD=0.6215p PS=2.67u PD=3.33u
M$29962 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$273663
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29963 \$272036 \$272035 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29964 \$272036 \$272033 \$272037 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29965 \$272037 \$272034 \$274087 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29966 VDD|pad|pin1|supply|vdd \$272039 \$274087 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29967 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$272039
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29968 VDD|pad|pin1|supply|vdd \$272037 \$272039 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29969 VDD|pad|pin1|supply|vdd \$272039 a1|i0|q$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29970 \$274514 \$274424 \$274532 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.31075p AD=0.383625p PS=2.23u PD=1.93u
M$29971 \$274533 d|s|z \$274514 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.55u AS=0.32995p AD=0.31075p PS=1.74u PD=2.23u
M$29972 VDD|pad|pin1|supply|vdd a1|i0|q$2 \$274533 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.91u AS=0.431325p AD=0.32995p PS=1.93u PD=1.74u
M$29973 \$274532 DATA|core|i0|i1|p2c VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=1.1u AS=0.383625p AD=0.431325p
+ PS=1.93u PD=1.93u
M$29974 VDD|pad|pin1|supply|vdd a2|zn$33 a2|i|s|zn VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$29975 a2|i|s|zn a1|i0|q$2 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$29976 \$274424 d|s|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.2904p PS=2.23u PD=1.6u
M$29977 VDD|pad|pin1|supply|vdd \$274514 d|z$93 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.77u AS=0.2904p AD=0.43505p PS=1.6u PD=2.67u
M$29978 VDD|pad|pin1|supply|vdd a3|zn$11 a2|zn$33 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29979 VDD|pad|pin1|supply|vdd a2|zn$34 a2|zn$33 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.4565p PS=2.67u PD=1.93u
M$29980 VDD|pad|pin1|supply|vdd a1|zn$23 a2|zn$33 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$29981 \$272042 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$29982 VDD|pad|pin1|supply|vdd \$272042 \$272043 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$29983 VDD|pad|pin1|supply|vdd \$272043 \$274118 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$29984 \$274118 d|s|z \$272044 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$29985 \$272044 \$272042 \$273664 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$29986 \$273664 \$272045 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$29987 VDD|pad|pin1|supply|vdd a4|zn$7 a2|zn$33 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29988 VDD|pad|pin1|supply|vdd a2|i|q$1 \$274535 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29989 VDD|pad|pin1|supply|vdd a1|b|d|z \$274535 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$29990 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$273664
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$29991 \$272045 \$272044 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$29992 \$272045 \$272042 \$272046 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$29993 \$272046 \$272043 \$274110 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$29994 VDD|pad|pin1|supply|vdd \$272048 \$274110 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$29995 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$272048
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$29996 VDD|pad|pin1|supply|vdd \$272046 \$272048 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$29997 VDD|pad|pin1|supply|vdd \$272048 a1|a2|q$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$29998 VDD|pad|pin1|supply|vdd \$274535 d|s|z VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$29999 a3|zn$10 a1|a2|q$4 \$275191 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30000 \$275191 a2|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$30001 d|s|zn CEB|a1|core|i|p2c \$275192 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30002 \$275192 a1|a2|q$1 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$30003 VDD|pad|pin1|supply|vdd a1|a2|q$4 \$274537 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30004 VDD|pad|pin1|supply|vdd a1|b|d|z \$274537 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30005 \$272050 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30006 VDD|pad|pin1|supply|vdd \$272050 \$272051 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30007 VDD|pad|pin1|supply|vdd \$274537 d|z$94 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30008 VDD|pad|pin1|supply|vdd \$272051 \$274120 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30009 \$274120 d|z$94 \$272052 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30010 \$272052 \$272050 \$273665 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30011 \$273665 \$272053 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30012 VDD|pad|pin1|supply|vdd cp|i|z$6 \$274515 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30013 VDD|pad|pin1|supply|vdd \$274515 \$274516 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30014 VDD|pad|pin1|supply|vdd \$274539 \$274517 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30015 \$274538 \$274515 \$274517 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30016 VDD|pad|pin1|supply|vdd \$274516 \$275193 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30017 \$275193 d|z$99 \$274538 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30018 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$273665
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30019 \$272053 \$272052 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30020 \$272053 \$272050 \$272054 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30021 \$272054 \$272051 \$274121 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30022 VDD|pad|pin1|supply|vdd \$272056 \$274121 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30023 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$272056
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30024 VDD|pad|pin1|supply|vdd \$272054 \$272056 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30025 VDD|pad|pin1|supply|vdd \$272056 a2|q$1 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30026 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$274517
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30027 \$274518 \$274516 \$275197 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30028 VDD|pad|pin1|supply|vdd \$275263 \$275197 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30029 VDD|pad|pin1|supply|vdd \$274538 \$274539 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30030 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$275263
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30031 VDD|pad|pin1|supply|vdd \$274518 \$275263 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30032 \$274539 \$274515 \$274518 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30033 VDD|pad|pin1|supply|vdd \$275263 a2|q$3 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30034 a4|zn$6 a1|a2|q \$274094 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30035 \$274094 a1|a2|b|q|s VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$30036 \$276915 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30037 VDD|pad|pin1|supply|vdd \$276915 \$276166 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30038 VDD|pad|pin1|supply|vdd \$276166 \$278681 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30039 \$278681 d|z$101 \$276916 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30040 \$276916 \$276915 \$277709 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30041 \$277709 \$276917 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30042 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$277709
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30043 \$276917 \$276916 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30044 \$276917 \$276915 \$276167 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30045 \$276167 \$276166 \$278688 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30046 VDD|pad|pin1|supply|vdd \$276919 \$278688 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30047 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$276919
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30048 VDD|pad|pin1|supply|vdd \$276167 \$276919 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30049 VDD|pad|pin1|supply|vdd \$276919 a1|a2|q$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30050 VDD|pad|pin1|supply|vdd a2|q$6 \$276921 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30051 \$276921 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30052 d|z$100 \$276921 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30053 a4|zn$8 a1|a2|q$6 \$278698 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30054 \$278698 a2|q$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$30055 VDD|pad|pin1|supply|vdd a3|zn$9 a2|zn$32 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30056 a2|zn$32 a2|zn$35 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.5675p PS=1.93u PD=2.67u
M$30057 VDD|pad|pin1|supply|vdd a1|z$17 a2|zn$32 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.5675p AD=0.6215p PS=2.67u PD=3.33u
M$30058 a2|zn$32 a4|zn$8 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30059 a2|zn$35 a1|a2|q$5 \$278706 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30060 \$278706 a2|q$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$30061 \$276924 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30062 VDD|pad|pin1|supply|vdd \$276924 \$276169 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30063 VDD|pad|pin1|supply|vdd \$276169 \$278719 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30064 \$278719 d|z$96 \$276925 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30065 \$276925 \$276924 \$277710 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30066 \$277710 \$276926 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30067 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$277710
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30068 \$276926 \$276925 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30069 \$276926 \$276924 \$276170 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30070 \$276170 \$276169 \$278732 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30071 VDD|pad|pin1|supply|vdd \$276928 \$278732 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30072 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$276928
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30073 VDD|pad|pin1|supply|vdd \$276170 \$276928 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30074 VDD|pad|pin1|supply|vdd \$276928 a1|a2|q$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30075 \$276929 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30076 VDD|pad|pin1|supply|vdd \$276929 \$276171 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30077 VDD|pad|pin1|supply|vdd \$276171 \$278741 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30078 \$278741 d|z$102 \$276930 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30079 \$276930 \$276929 \$277711 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30080 \$277711 \$276931 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30081 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$277711
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30082 \$276931 \$276930 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30083 \$276931 \$276929 \$276172 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30084 \$276172 \$276171 \$278751 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30085 VDD|pad|pin1|supply|vdd \$276933 \$278751 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30086 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$276933
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30087 VDD|pad|pin1|supply|vdd \$276172 \$276933 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30088 VDD|pad|pin1|supply|vdd \$276933 a2|q$4 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30089 \$276935 cp|i|z$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30090 VDD|pad|pin1|supply|vdd \$276935 \$276173 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30091 VDD|pad|pin1|supply|vdd \$276173 \$278759 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30092 \$278759 d|z$103 \$276936 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30093 \$276936 \$276935 \$277712 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30094 \$277712 \$276937 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30095 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$277712
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30096 \$276937 \$276936 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30097 \$276937 \$276935 \$276174 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30098 \$276174 \$276173 \$278771 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30099 VDD|pad|pin1|supply|vdd \$276939 \$278771 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30100 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$276939
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30101 VDD|pad|pin1|supply|vdd \$276174 \$276939 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30102 VDD|pad|pin1|supply|vdd \$276939 a1|a2|q$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30103 \$276941 cp|i|z$6 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30104 VDD|pad|pin1|supply|vdd \$276941 \$276175 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30105 VDD|pad|pin1|supply|vdd \$276175 \$278782 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30106 \$278782 d|z$104 \$276942 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30107 \$276942 \$276941 \$277713 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30108 \$277713 \$276943 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30109 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$277713
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30110 \$276943 \$276942 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30111 \$276943 \$276941 \$276176 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30112 \$276176 \$276175 \$278773 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30113 VDD|pad|pin1|supply|vdd \$276945 \$278773 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30114 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$276945
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30115 VDD|pad|pin1|supply|vdd \$276176 \$276945 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30116 VDD|pad|pin1|supply|vdd \$276945 a2|q$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30117 VDD|pad|pin1|supply|vdd a1|a2|q$6 \$279198 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30118 VDD|pad|pin1|supply|vdd a1|b|d|z \$279198 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30119 VDD|pad|pin1|supply|vdd \$279198 d|z$105 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30120 VDD|pad|pin1|supply|vdd a2|q$2 \$279200 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30121 VDD|pad|pin1|supply|vdd a1|b|d|z \$279200 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30122 VDD|pad|pin1|supply|vdd \$279200 d|z$101 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30123 VDD|pad|pin1|supply|vdd cp|i|z$7 \$279142 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30124 VDD|pad|pin1|supply|vdd \$279142 \$279143 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30125 VDD|pad|pin1|supply|vdd \$279255 \$279144 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30126 \$279201 \$279142 \$279144 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30127 VDD|pad|pin1|supply|vdd \$279143 \$279251 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30128 \$279251 d|z$100 \$279201 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30129 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$279144
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30130 \$279145 \$279143 \$279250 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30131 VDD|pad|pin1|supply|vdd \$279556 \$279250 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30132 VDD|pad|pin1|supply|vdd \$279201 \$279255 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30133 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$279556
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30134 VDD|pad|pin1|supply|vdd \$279145 \$279556 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30135 \$279255 \$279142 \$279145 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30136 VDD|pad|pin1|supply|vdd \$279556 a1|a2|q$5 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30137 VDD|pad|pin1|supply|vdd cp|i|z$5 \$279146 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30138 VDD|pad|pin1|supply|vdd \$279146 \$279147 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30139 VDD|pad|pin1|supply|vdd \$279256 \$279148 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30140 \$279202 \$279146 \$279148 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30141 VDD|pad|pin1|supply|vdd \$279147 \$279249 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30142 \$279249 d|z$106 \$279202 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30143 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$279148
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30144 \$279149 \$279147 \$279248 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30145 VDD|pad|pin1|supply|vdd \$279557 \$279248 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30146 VDD|pad|pin1|supply|vdd \$279202 \$279256 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30147 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$279557
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30148 VDD|pad|pin1|supply|vdd \$279149 \$279557 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30149 \$279256 \$279146 \$279149 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30150 VDD|pad|pin1|supply|vdd \$279557 a2|i|q$2 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30151 VDD|pad|pin1|supply|vdd cp|i|z$5 \$279150 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30152 VDD|pad|pin1|supply|vdd \$279150 \$279151 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30153 VDD|pad|pin1|supply|vdd \$279257 \$279152 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30154 \$279203 \$279150 \$279152 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30155 VDD|pad|pin1|supply|vdd \$279151 \$279246 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30156 \$279246 d|z$97 \$279203 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30157 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$279152
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30158 \$279153 \$279151 \$279247 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30159 VDD|pad|pin1|supply|vdd \$279558 \$279247 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30160 VDD|pad|pin1|supply|vdd \$279203 \$279257 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30161 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$279558
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30162 VDD|pad|pin1|supply|vdd \$279153 \$279558 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30163 \$279257 \$279150 \$279153 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30164 VDD|pad|pin1|supply|vdd \$279558 a1|a2|q$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30165 VDD|pad|pin1|supply|vdd cp|i|z$5 \$279154 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30166 VDD|pad|pin1|supply|vdd \$279154 \$279155 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30167 VDD|pad|pin1|supply|vdd \$279258 \$279156 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30168 \$279205 \$279154 \$279156 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30169 VDD|pad|pin1|supply|vdd \$279155 \$279245 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30170 \$279245 d|z$107 \$279205 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30171 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$279156
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30172 \$279157 \$279155 \$279244 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30173 VDD|pad|pin1|supply|vdd \$279559 \$279244 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30174 VDD|pad|pin1|supply|vdd \$279205 \$279258 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30175 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$279559
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30176 VDD|pad|pin1|supply|vdd \$279157 \$279559 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30177 \$279258 \$279154 \$279157 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30178 VDD|pad|pin1|supply|vdd \$279559 a2|q$8 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30179 a4|zn$7 a1|a2|q$2 \$279534 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30180 \$279534 a2|q$8 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$30181 VDD|pad|pin1|supply|vdd cp|i|z$6 \$279158 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30182 VDD|pad|pin1|supply|vdd \$279158 \$279159 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30183 VDD|pad|pin1|supply|vdd \$279259 \$279160 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.394325p AD=0.1336375p PS=3.22u PD=1.16u
M$30184 \$279207 \$279158 \$279160 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30185 VDD|pad|pin1|supply|vdd \$279159 \$279243 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30186 \$279243 d|z$108 \$279207 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30187 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$279160
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30188 \$279161 \$279159 \$279242 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30189 VDD|pad|pin1|supply|vdd \$279560 \$279242 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30190 VDD|pad|pin1|supply|vdd \$279207 \$279259 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.349425p AD=0.3857125p PS=2.285u PD=1.86u
M$30191 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$279560
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30192 VDD|pad|pin1|supply|vdd \$279161 \$279560 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30193 \$279259 \$279158 \$279161 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30194 VDD|pad|pin1|supply|vdd \$279560 a1|a2|q$9 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30195 VDD|pad|pin1|supply|vdd a1|a2|q$9 \$279208 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30196 VDD|pad|pin1|supply|vdd a1|b|d|z \$279208 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30197 VDD|pad|pin1|supply|vdd \$279208 d|z$104 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30198 VDD|pad|pin1|supply|vdd a2|q$5 \$279209 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30199 VDD|pad|pin1|supply|vdd a1|b|d|z \$279209 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30200 VDD|pad|pin1|supply|vdd \$279209 d|z$99 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.6215p PS=4.81u PD=3.33u
M$30201 \$280738 cp|i|z$7 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30202 VDD|pad|pin1|supply|vdd \$280738 \$280723 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30203 VDD|pad|pin1|supply|vdd \$280723 \$282471 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30204 \$282471 d|z$105 \$280739 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30205 \$280739 \$280738 \$282153 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30206 \$282153 \$280740 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30207 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$282153
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30208 \$280740 \$280739 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30209 \$280740 \$280738 \$280724 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30210 \$280724 \$280723 \$282483 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30211 VDD|pad|pin1|supply|vdd \$280742 \$282483 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30212 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$280742
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30213 VDD|pad|pin1|supply|vdd \$280724 \$280742 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30214 VDD|pad|pin1|supply|vdd \$280742 a2|q$6 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30215 \$280743 cp|i|z$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.31075p AD=0.33925p PS=2.23u PD=2.12u
M$30216 VDD|pad|pin1|supply|vdd \$280743 \$280725 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.55u AS=0.33925p AD=0.31075p PS=2.12u PD=2.23u
M$30217 VDD|pad|pin1|supply|vdd \$280725 \$282463 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.81u AS=0.67965p AD=0.33615p PS=4.23u PD=1.64u
M$30218 \$282463 d|z$95 \$280744 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.81u AS=0.33615p AD=0.27255p PS=1.64u PD=1.64u
M$30219 \$280744 \$280743 \$282154 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.33u AS=0.27255p AD=0.1336375p PS=1.64u PD=1.16u
M$30220 \$282154 \$280745 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.305u AS=0.1336375p AD=0.394325p PS=1.16u PD=3.22u
M$30221 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$282154
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.275u AS=0.349425p
+ AD=0.162875p PS=2.285u PD=1.73u
M$30222 \$280745 \$280744 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.715u AS=0.3857125p AD=0.349425p PS=1.86u PD=2.285u
M$30223 \$280745 \$280743 \$280726 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=1.03u AS=0.3857125p AD=0.3274125p PS=1.86u PD=1.86u
M$30224 \$280726 \$280725 \$282425 VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u
+ W=0.275u AS=0.3274125p AD=0.114125p PS=1.86u PD=1.105u
M$30225 VDD|pad|pin1|supply|vdd \$280747 \$282425 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.275u AS=0.4271125p AD=0.114125p PS=2.56u PD=1.105u
M$30226 VDD|pad|pin1|supply|vdd RST|a1|b|cdn|core|i|p2c \$280747
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=0.99u AS=0.4271125p
+ AD=0.41085p PS=2.56u PD=1.82u
M$30227 VDD|pad|pin1|supply|vdd \$280726 \$280747 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=0.99u AS=0.552925p AD=0.41085p PS=2.67u PD=1.82u
M$30228 VDD|pad|pin1|supply|vdd \$280747 a2|q$7 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.552925p AD=0.6215p PS=2.67u PD=3.33u
M$30229 VDD|pad|pin1|supply|vdd a2|q$7 \$280748 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30230 \$280748 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30231 d|z$106 \$280748 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30232 VDD|pad|pin1|supply|vdd a1|a2|q$8 \$280749 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30233 \$280749 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30234 d|z$102 \$280749 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30235 VDD|pad|pin1|supply|vdd a2|q$4 \$280750 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30236 \$280750 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30237 d|z$107 \$280750 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30238 a3|zn$11 a1|a2|q$8 \$282412 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30239 \$282412 a2|q$4 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$30240 VDD|pad|pin1|supply|vdd a2|q$8 \$280751 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30241 \$280751 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30242 d|z$103 \$280751 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30243 a2|zn$34 a1|a2|q$7 \$282375 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30244 \$282375 a2|q$3 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$30245 VDD|pad|pin1|supply|vdd a1|a2|q$7 \$280752 VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.8435p AD=0.4565p PS=4.81u PD=1.93u
M$30246 \$280752 a1|b|d|z VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.8435p PS=1.93u PD=4.81u
M$30247 d|z$108 \$280752 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.6215p AD=0.8435p PS=3.33u PD=4.81u
M$30248 a1|zn$23 a1|a2|q$9 \$282333 VDD|pad|pin1|supply|vdd sg13_lv_pmos
+ L=0.13u W=1.1u AS=0.6215p AD=0.4565p PS=3.33u PD=1.93u
M$30249 \$282333 a2|q$5 VDD|pad|pin1|supply|vdd VDD|pad|pin1|supply|vdd
+ sg13_lv_pmos L=0.13u W=1.1u AS=0.4565p AD=0.6215p PS=1.93u PD=3.33u
M$30250 CEB|a1|core|i|p2c \$286830 VDD|pad|pin1|supply|vdd
+ VDD|pad|pin1|supply|vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p
+ PS=10.18u PD=10.18u
M$30251 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$50381
+ AVDD|anode|cathode|pad|vdd VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30271 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate
+ anode|cathode|pad|pad_adc_result_0_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$30279 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$1
+ anode|cathode|pad|pad_adc_result_1_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$30287 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$2
+ anode|cathode|pad|pad_adc_result_2_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$30295 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$3
+ anode|cathode|pad|pad_adc_result_3_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$30303 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$4
+ anode|cathode|pad|pad_adc_result_4_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$30311 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$5
+ anode|cathode|pad|pad_adc_valid_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=106.56u AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$30319 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$6
+ anode|cathode|pad|pad_adc_sample_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=106.56u
+ AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$30403 VDD|pad|pin1|supply|vdd core \$64423 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$30404 VDD|pad|pin1|supply|vdd core$1 \$64425 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$30405 \$63424 \$63425 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30406 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63424 \$63425
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30407 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63425 gate|ngate|o
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30408 \$63426 \$63427 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30409 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63426 \$63427
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30410 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63427 gate|o|pgate
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30411 \$63428 \$63429 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30412 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63428 \$63429
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30413 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63429 gate|ngate|o$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30414 \$63430 \$63431 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30415 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63430 \$63431
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30416 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63431 gate|o|pgate$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30417 \$63432 \$63433 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30418 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63432 \$63433
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30419 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63433 gate|ngate|o$2
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30420 \$63434 \$63435 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30421 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63434 \$63435
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30422 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63435 gate|o|pgate$2
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30423 \$63436 \$63437 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30424 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63436 \$63437
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30425 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63437 gate|ngate|o$3
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30426 \$63438 \$63439 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30427 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63438 \$63439
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30428 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63439 gate|o|pgate$3
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30429 \$63440 \$63441 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30430 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63440 \$63441
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30431 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63441 gate|ngate|o$4
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30432 \$63442 \$63443 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30433 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63442 \$63443
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30434 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63443 gate|o|pgate$4
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30435 \$63444 \$63445 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30436 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63444 \$63445
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30437 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63445 gate|ngate|o$5
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30438 \$63446 \$63447 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30439 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63446 \$63447
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30440 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63447 gate|o|pgate$5
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30441 \$63448 \$63449 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30442 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63448 \$63449
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30443 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63449 gate|ngate|o$6
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30444 \$63450 \$63451 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30445 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63450 \$63451
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30446 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$63451 gate|o|pgate$6
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30447 VDD|pad|pin1|supply|vdd core$2 \$90574 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$30448 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$104194
+ anode|cathode|pad|pad_adc_vrefp_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30488 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$123894
+ anode|cathode|pad|pad_adc_vrefn_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30508 VDD|pad|pin1|supply|vdd in|pin2 gate|out VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.5u W=350u AS=67.55p AD=67.55p PS=376.3u PD=376.3u
M$30578 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$148329
+ anode|cathode|pad|pad_adc_vin_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30618 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$166060
+ anode|cathode|pad|pad_adc_vip_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=266.4u AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30658 VDDIO|cathode|guard|iovdd|pad|pin1|supply in|pin2$1 gate|out$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.5u W=350u
+ AS=67.55p AD=67.55p PS=376.3u PD=376.3u
M$30708 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$192134 anode|cathode|pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30748 VDDIO|cathode|guard|iovdd|pad|pin1|supply gate|o|pgate$7
+ anode|cathode|pad|pad_miso_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ sg13_hv_pmos L=0.6u W=106.56u AS=50.4828p AD=50.4828p PS=135.04u PD=135.04u
M$30764 \$200627 \$201363 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30765 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$200627 \$201363
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30766 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$201363 gate|ngate|o$7
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30767 \$202320 \$202581 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$30768 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$202320 \$202581
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$30769 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$202581 gate|o|pgate$7
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.45u W=3.9u
+ AS=1.326p AD=1.326p PS=8.48u PD=8.48u
M$30770 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$220269 anode|cathode|pad$1
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30810 VDD|pad|pin1|supply|vdd core$3 \$231093 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$30811 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$252800 anode|cathode|pad$2
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30851 VDD|pad|pin1|supply|vdd core$4 \$258894 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$30852 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$276914 anode|cathode|pad$3
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30892 VDD|pad|pin1|supply|vdd core$5 \$286830 VDD|pad|pin1|supply|vdd
+ sg13_hv_pmos L=0.45u W=4.65u AS=1.581p AD=1.581p PS=9.98u PD=9.98u
M$30893 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$323983 anode|cathode|pad$4
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30913 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$323984 anode|cathode|pad$5
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30933 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$323985 anode|cathode|pad$6
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30953 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$323986 anode|cathode|pad$7
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30973 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$323987 anode|cathode|pad$8
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$30993 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$323988 anode|cathode|pad$9
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$31013 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$323989 anode|cathode|pad$10
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$31033 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$323990 anode|cathode|pad$11
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$31053 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$323991 anode|cathode|pad$12
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
M$31073 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$323992 anode|cathode|pad$13
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply sg13_hv_pmos L=0.6u W=266.4u
+ AS=123.21p AD=123.21p PS=316.72u PD=316.72u
D$31293 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_rst_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31295 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_clk_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31297 VSS|anode|cathode|vss gate|ngate|o dantenna A=0.6084p P=3.12u m=1
D$31298 VSS|anode|cathode|vss gate|ngate|o$1 dantenna A=0.6084p P=3.12u m=1
D$31299 VSS|anode|cathode|vss gate|ngate|o$2 dantenna A=0.6084p P=3.12u m=1
D$31300 VSS|anode|cathode|vss gate|ngate|o$3 dantenna A=0.6084p P=3.12u m=1
D$31301 VSS|anode|cathode|vss gate|ngate|o$4 dantenna A=0.6084p P=3.12u m=1
D$31302 VSS|anode|cathode|vss gate|ngate|o$5 dantenna A=0.6084p P=3.12u m=1
D$31303 VSS|anode|cathode|vss gate|ngate|o$6 dantenna A=0.6084p P=3.12u m=1
D$31304 VSS|anode|cathode|vss AVDD|anode|cathode|pad|vdd dantenna A=35.0028p
+ P=58.08u m=2
D$31305 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_result_0_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31306 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_result_1_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31307 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_result_2_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31308 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_result_3_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31309 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_result_4_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31310 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_valid_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31311 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_sample_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31313 VSS|anode|cathode|vss core|padres dantenna A=1.984p P=7.48u m=1
D$31314 VSS|anode|cathode|vss core dantenna A=1.984p P=7.48u m=1
D$31315 VSS|anode|cathode|vss core$1 dantenna A=1.984p P=7.48u m=1
D$31323 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_go_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31325 VSS|anode|cathode|vss core$2 dantenna A=1.984p P=7.48u m=1
D$31326 VSS|anode|cathode|vss VSS|anode|cathode|vss dantenna A=35.0028p
+ P=58.08u m=4
D$31330 VSS|anode|cathode|vss VREFH|core|padres dantenna A=1.984p P=7.48u m=1
D$31331 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_vrefp_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31333 VSS|anode|cathode|vss VREFL|core|padres dantenna A=1.984p P=7.48u m=1
D$31334 VSS|anode|cathode|vss gate|out dantenna A=0.2304p P=1.92u m=1
D$31335 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_vrefn_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31337 VSS|anode|cathode|vss VSSIO|anode|cathode|guard|iovss dantenna
+ A=35.0028p P=58.08u m=2
D$31339 VSS|anode|cathode|vss VIN|core|padres dantenna A=1.984p P=7.48u m=1
D$31340 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_vin_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31342 VSS|anode|cathode|vss VALID|a3|c2p|core|i|z dantenna A=1.44045p P=4.91u
+ m=2
D$31343 VSS|anode|cathode|vss SAMPLE|a1|c2p|core|i|z dantenna A=1.44045p
+ P=4.91u m=2
D$31344 VSS|anode|cathode|vss VIP|core|padres dantenna A=1.984p P=7.48u m=1
D$31347 VSS|anode|cathode|vss gate|out$1 dantenna A=0.2304p P=1.92u m=1
D$31348 VSS|anode|cathode|vss anode|cathode|pad|pad_adc_vip_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31350 VSS|anode|cathode|vss core|padres$1 dantenna A=1.984p P=7.48u m=1
D$31351 VSS|anode|cathode|vss gate|ngate|o$7 dantenna A=0.6084p P=3.12u m=1
D$31352 VSS|anode|cathode|vss anode|cathode|pad dantenna A=35.0028p P=58.08u m=2
D$31354 VSS|anode|cathode|vss anode|cathode|pad|pad_miso_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31356 VSS|anode|cathode|vss core|padres$2 dantenna A=1.984p P=7.48u m=1
D$31357 VSS|anode|cathode|vss anode|cathode|pad|pad_mosi_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31359 VSS|anode|cathode|vss anode|cathode|pad$1 dantenna A=35.0028p P=58.08u
+ m=2
D$31361 VSS|anode|cathode|vss core$3 dantenna A=1.984p P=7.48u m=1
D$31362 VSS|anode|cathode|vss anode|cathode|pad|pad_sclk_pad dantenna
+ A=35.0028p P=58.08u m=2
D$31364 VSS|anode|cathode|vss core|padres$3 dantenna A=1.984p P=7.48u m=1
D$31365 VSS|anode|cathode|vss anode|cathode|pad$2 dantenna A=35.0028p P=58.08u
+ m=2
D$31367 VSS|anode|cathode|vss core$4 dantenna A=1.984p P=7.48u m=1
D$31368 VSS|anode|cathode|vss anode|cathode|pad|pad_cs_pad dantenna A=35.0028p
+ P=58.08u m=2
D$31370 VSS|anode|cathode|vss core|padres$4 dantenna A=1.984p P=7.48u m=1
D$31371 VSS|anode|cathode|vss anode|cathode|pad$3 dantenna A=35.0028p P=58.08u
+ m=2
D$31373 VSS|anode|cathode|vss core$5 dantenna A=1.984p P=7.48u m=1
D$31374 VSS|anode|cathode|vss core|padres$5 dantenna A=1.984p P=7.48u m=1
D$31375 VSS|anode|cathode|vss core|padres$6 dantenna A=1.984p P=7.48u m=1
D$31376 VSS|anode|cathode|vss core|padres$7 dantenna A=1.984p P=7.48u m=1
D$31377 VSS|anode|cathode|vss core|padres$8 dantenna A=1.984p P=7.48u m=1
D$31378 VSS|anode|cathode|vss core|padres$9 dantenna A=1.984p P=7.48u m=1
D$31379 VSS|anode|cathode|vss core|padres$10 dantenna A=1.984p P=7.48u m=1
D$31380 VSS|anode|cathode|vss core|padres$11 dantenna A=1.984p P=7.48u m=1
D$31381 VSS|anode|cathode|vss core|padres$12 dantenna A=1.984p P=7.48u m=1
D$31382 VSS|anode|cathode|vss core|padres$13 dantenna A=1.984p P=7.48u m=1
D$31383 VSS|anode|cathode|vss core|padres$14 dantenna A=1.984p P=7.48u m=1
D$31384 VSS|anode|cathode|vss anode|cathode|pad$4 dantenna A=35.0028p P=58.08u
+ m=2
D$31385 VSS|anode|cathode|vss anode|cathode|pad$5 dantenna A=35.0028p P=58.08u
+ m=2
D$31386 VSS|anode|cathode|vss anode|cathode|pad$6 dantenna A=35.0028p P=58.08u
+ m=2
D$31387 VSS|anode|cathode|vss anode|cathode|pad$7 dantenna A=35.0028p P=58.08u
+ m=2
D$31388 VSS|anode|cathode|vss anode|cathode|pad$8 dantenna A=35.0028p P=58.08u
+ m=2
D$31389 VSS|anode|cathode|vss anode|cathode|pad$9 dantenna A=35.0028p P=58.08u
+ m=2
D$31390 VSS|anode|cathode|vss anode|cathode|pad$10 dantenna A=35.0028p P=58.08u
+ m=2
D$31391 VSS|anode|cathode|vss anode|cathode|pad$11 dantenna A=35.0028p P=58.08u
+ m=2
D$31392 VSS|anode|cathode|vss anode|cathode|pad$12 dantenna A=35.0028p P=58.08u
+ m=2
D$31393 VSS|anode|cathode|vss anode|cathode|pad$13 dantenna A=35.0028p P=58.08u
+ m=2
D$31404 AVDD|anode|cathode|pad|vdd VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=35.0028p P=58.08u m=2
D$31405 anode|cathode|pad|pad_adc_result_0_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31406 anode|cathode|pad|pad_adc_result_1_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31407 anode|cathode|pad|pad_adc_result_2_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31408 anode|cathode|pad|pad_adc_result_3_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31409 anode|cathode|pad|pad_adc_result_4_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31410 anode|cathode|pad|pad_adc_valid_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31411 anode|cathode|pad|pad_adc_sample_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31420 anode|cathode|pad|pad_adc_rst_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31422 anode|cathode|pad|pad_adc_clk_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31424 gate|o|pgate VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$31425 gate|o|pgate$1 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$31426 gate|o|pgate$2 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$31427 gate|o|pgate$3 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$31428 gate|o|pgate$4 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$31429 gate|o|pgate$5 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$31430 gate|o|pgate$6 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$31431 VSS|anode|cathode|vss VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=35.0028p P=58.08u m=4
D$31433 VREFH|core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31434 core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31435 core VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$31436 core$1 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$31437 core$2 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$31438 anode|cathode|pad|pad_adc_go_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31442 anode|cathode|pad|pad_adc_vrefp_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31444 anode|cathode|pad|pad_adc_vrefn_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31446 VREFL|core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31447 VIN|core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31448 VSSIO|anode|cathode|guard|iovss
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31450 anode|cathode|pad|pad_adc_vin_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31452 VALID|a3|c2p|core|i|z VDD|pad|pin1|supply|vdd dpantenna A=1.44045p
+ P=4.91u m=2
D$31454 SAMPLE|a1|c2p|core|i|z VDD|pad|pin1|supply|vdd dpantenna A=1.44045p
+ P=4.91u m=2
D$31456 anode|cathode|pad|pad_adc_vip_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31458 VIP|core|padres VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31459 anode|cathode|pad VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=35.0028p P=58.08u m=2
D$31461 core|padres$1 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31462 gate|o|pgate$7 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=0.2304p P=1.92u m=1
D$31463 anode|cathode|pad|pad_miso_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31465 anode|cathode|pad$1 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=35.0028p P=58.08u m=2
D$31467 core|padres$2 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31468 anode|cathode|pad|pad_mosi_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31470 core$3 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$31471 anode|cathode|pad|pad_sclk_pad
+ VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=35.0028p P=58.08u m=2
D$31473 core|padres$3 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31474 anode|cathode|pad$2 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=35.0028p P=58.08u m=2
D$31476 core$4 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$31477 anode|cathode|pad|pad_cs_pad VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=35.0028p P=58.08u m=2
D$31479 core|padres$4 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31480 anode|cathode|pad$3 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=35.0028p P=58.08u m=2
D$31482 core|padres$5 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31483 core|padres$6 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31484 core|padres$7 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31485 core|padres$8 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31486 core|padres$9 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31487 core|padres$10 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31488 core|padres$11 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31489 core|padres$12 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31490 core|padres$13 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31491 core|padres$14 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=3.1872p P=11.24u m=1
D$31492 core$5 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna A=3.1872p
+ P=11.24u m=1
D$31493 anode|cathode|pad$4 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=35.0028p P=58.08u m=2
D$31494 anode|cathode|pad$5 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=35.0028p P=58.08u m=2
D$31495 anode|cathode|pad$6 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=35.0028p P=58.08u m=2
D$31496 anode|cathode|pad$7 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=35.0028p P=58.08u m=2
D$31497 anode|cathode|pad$8 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=35.0028p P=58.08u m=2
D$31498 anode|cathode|pad$9 VDDIO|cathode|guard|iovdd|pad|pin1|supply dpantenna
+ A=35.0028p P=58.08u m=2
D$31499 anode|cathode|pad$10 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=35.0028p P=58.08u m=2
D$31500 anode|cathode|pad$11 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=35.0028p P=58.08u m=2
D$31501 anode|cathode|pad$12 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=35.0028p P=58.08u m=2
D$31502 anode|cathode|pad$13 VDDIO|cathode|guard|iovdd|pad|pin1|supply
+ dpantenna A=35.0028p P=58.08u m=2
R$31513 VSSIO|anode|cathode|guard|iovss \$40710 rppd w=0.5u l=3.54u ps=0 b=0 m=1
R$31514 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$50381 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31515 AVDD|anode|cathode|pad|vdd core|padres rppd w=1u l=2u ps=0 b=0 m=1
R$31516 anode|cathode|pad|pad_adc_rst_pad core rppd w=1u l=2u ps=0 b=0 m=1
R$31517 anode|cathode|pad|pad_adc_clk_pad core$1 rppd w=1u l=2u ps=0 b=0 m=1
R$31518 VSSIO|anode|cathode|guard|iovss \$104193 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31519 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$104194 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31520 core$2 anode|cathode|pad|pad_adc_go_pad rppd w=1u l=2u ps=0 b=0 m=1
R$31521 VSSIO|anode|cathode|guard|iovss \$123893 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31522 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$123894 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31523 anode|cathode|pad|pad_adc_vrefp_pad VREFH|core|padres rppd w=1u l=2u
+ ps=0 b=0 m=1
R$31529 anode|cathode|pad|pad_adc_vrefn_pad VREFL|core|padres rppd w=1u l=2u
+ ps=0 b=0 m=1
R$31549 VDD|pad|pin1|supply|vdd in|pin2 rppd w=1u l=520u ps=0 b=0 m=1
R$31551 VSSIO|anode|cathode|guard|iovss \$144910 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31552 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$148329 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31553 VSSIO|anode|cathode|guard|iovss \$166059 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31554 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$166060 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31555 anode|cathode|pad|pad_adc_vin_pad VIN|core|padres rppd w=1u l=2u ps=0
+ b=0 m=1
R$31561 anode|cathode|pad|pad_adc_vip_pad VIP|core|padres rppd w=1u l=2u ps=0
+ b=0 m=1
R$31582 in|pin2$1 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=1u l=520u
+ ps=0 b=0 m=1
R$31583 VSSIO|anode|cathode|guard|iovss \$192133 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31584 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$192134 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31585 VSSIO|anode|cathode|guard|iovss \$220268 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31586 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$220269 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31587 anode|cathode|pad core|padres$1 rppd w=1u l=2u ps=0 b=0 m=1
R$31588 anode|cathode|pad$1 core|padres$2 rppd w=1u l=2u ps=0 b=0 m=1
R$31589 core$3 anode|cathode|pad|pad_mosi_pad rppd w=1u l=2u ps=0 b=0 m=1
R$31590 VSSIO|anode|cathode|guard|iovss \$249093 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31591 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$252800 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31592 anode|cathode|pad$2 core|padres$3 rppd w=1u l=2u ps=0 b=0 m=1
R$31593 core$4 anode|cathode|pad|pad_sclk_pad rppd w=1u l=2u ps=0 b=0 m=1
R$31594 VSSIO|anode|cathode|guard|iovss \$276913 rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31595 VDDIO|cathode|guard|iovdd|pad|pin1|supply \$276914 rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31596 anode|cathode|pad$3 core|padres$4 rppd w=1u l=2u ps=0 b=0 m=1
R$31597 core$5 anode|cathode|pad|pad_cs_pad rppd w=1u l=2u ps=0 b=0 m=1
R$31598 core|padres$5 anode|cathode|pad$4 rppd w=1u l=2u ps=0 b=0 m=1
R$31599 core|padres$6 anode|cathode|pad$5 rppd w=1u l=2u ps=0 b=0 m=1
R$31600 core|padres$7 anode|cathode|pad$6 rppd w=1u l=2u ps=0 b=0 m=1
R$31601 core|padres$8 anode|cathode|pad$7 rppd w=1u l=2u ps=0 b=0 m=1
R$31602 core|padres$9 anode|cathode|pad$8 rppd w=1u l=2u ps=0 b=0 m=1
R$31603 core|padres$10 anode|cathode|pad$9 rppd w=1u l=2u ps=0 b=0 m=1
R$31604 core|padres$11 anode|cathode|pad$10 rppd w=1u l=2u ps=0 b=0 m=1
R$31605 core|padres$12 anode|cathode|pad$11 rppd w=1u l=2u ps=0 b=0 m=1
R$31606 core|padres$13 anode|cathode|pad$12 rppd w=1u l=2u ps=0 b=0 m=1
R$31607 core|padres$14 anode|cathode|pad$13 rppd w=1u l=2u ps=0 b=0 m=1
R$31608 \$323983 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31609 \$323984 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31610 \$323985 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31611 \$323986 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31612 \$323987 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31613 \$323988 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31614 \$323989 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31615 \$323990 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31616 \$323991 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31617 \$323992 VDDIO|cathode|guard|iovdd|pad|pin1|supply rppd w=0.5u l=12.9u
+ ps=0 b=0 m=1
R$31618 \$335158 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31619 \$335159 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31620 \$335160 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31621 \$335161 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31622 \$335162 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31623 \$335163 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31624 \$335164 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31625 \$335165 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31626 \$335166 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
R$31627 \$335167 VSSIO|anode|cathode|guard|iovss rppd w=0.5u l=3.54u ps=0 b=0
+ m=1
.ENDS asicone_202508
