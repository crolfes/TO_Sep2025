magic
tech ihp-sg13g2
magscale 1 2
timestamp 1756453207
<< metal1 >>
rect 4000 300 10800 400
rect 4000 -100 4120 300
rect 4260 161 10800 200
rect 4260 160 4981 161
rect 4260 42 4380 160
rect 4500 42 4981 160
rect 4260 41 4981 42
rect 5103 41 5585 161
rect 5707 41 6189 161
rect 6311 41 6793 161
rect 6915 41 7397 161
rect 7519 41 8001 161
rect 8123 41 8605 161
rect 8727 41 9209 161
rect 9331 41 9813 161
rect 9935 41 10800 161
rect 4260 0 10800 41
rect 4000 -115 10800 -100
rect 4000 -203 4220 -115
rect 4310 -203 4570 -115
rect 4000 -205 4570 -203
rect 4660 -205 4820 -115
rect 4910 -205 5180 -115
rect 5270 -205 5430 -115
rect 5520 -205 5780 -115
rect 5870 -205 6030 -115
rect 6120 -205 6390 -115
rect 6480 -205 6640 -115
rect 6730 -205 6990 -115
rect 7080 -205 7240 -115
rect 7330 -205 7590 -115
rect 7680 -205 7840 -115
rect 7930 -205 8200 -115
rect 8290 -205 8450 -115
rect 8540 -205 8800 -115
rect 8890 -205 9050 -115
rect 9140 -205 9410 -115
rect 9500 -205 9660 -115
rect 9750 -205 10010 -115
rect 10100 -205 10800 -115
rect 4000 -240 10800 -205
rect -840 -2220 2000 -2200
rect -840 -2280 -820 -2220
rect 1980 -2280 2000 -2220
rect -840 -2300 2000 -2280
rect 2200 -2460 4080 -2440
rect 2200 -2580 2220 -2460
rect 4060 -2580 4080 -2460
rect 2200 -2600 4080 -2580
<< via1 >>
rect 4380 42 4500 160
rect 4981 41 5103 161
rect 5585 41 5707 161
rect 6189 41 6311 161
rect 6793 41 6915 161
rect 7397 41 7519 161
rect 8001 41 8123 161
rect 8605 41 8727 161
rect 9209 41 9331 161
rect 9813 41 9935 161
rect 4220 -203 4310 -115
rect 4570 -205 4660 -115
rect 4820 -205 4910 -115
rect 5180 -205 5270 -115
rect 5430 -205 5520 -115
rect 5780 -205 5870 -115
rect 6030 -205 6120 -115
rect 6390 -205 6480 -115
rect 6640 -205 6730 -115
rect 6990 -205 7080 -115
rect 7240 -205 7330 -115
rect 7590 -205 7680 -115
rect 7840 -205 7930 -115
rect 8200 -205 8290 -115
rect 8450 -205 8540 -115
rect 8800 -205 8890 -115
rect 9050 -205 9140 -115
rect 9410 -205 9500 -115
rect 9660 -205 9750 -115
rect 10010 -205 10100 -115
rect -820 -2280 1980 -2220
rect 2220 -2580 4060 -2460
<< metal2 >>
rect 4600 394 4910 400
rect 5200 397 5520 400
rect 4060 -80 4320 320
rect 4220 -115 4320 -80
rect 4310 -120 4320 -115
rect 4380 160 4500 169
rect 4220 -345 4310 -203
rect 4380 -320 4500 42
rect 4570 -60 4910 394
rect 4570 -115 4660 -60
rect 4820 -115 4910 -60
rect 4981 161 5103 170
rect 4561 -205 4570 -115
rect 4660 -205 4669 -115
rect 4811 -205 4820 -115
rect 4910 -205 4919 -115
rect 4570 -304 4660 -205
rect 4820 -325 4910 -205
rect 4981 -361 5103 41
rect 5180 -60 5520 397
rect 5180 -115 5270 -60
rect 5430 -115 5520 -60
rect 5585 161 5707 170
rect 5171 -205 5180 -115
rect 5270 -205 5279 -115
rect 5421 -205 5430 -115
rect 5520 -205 5529 -115
rect 5180 -290 5270 -205
rect 5430 -305 5520 -205
rect 5585 -361 5707 41
rect 5780 -60 6120 400
rect 5780 -115 5870 -60
rect 6030 -115 6120 -60
rect 6189 161 6311 170
rect 5771 -205 5780 -115
rect 5870 -205 5879 -115
rect 6021 -205 6030 -115
rect 6120 -205 6129 -115
rect 5780 -325 5870 -205
rect 6030 -305 6120 -205
rect 6189 -361 6311 41
rect 6390 -60 6730 400
rect 6390 -115 6480 -60
rect 6640 -115 6730 -60
rect 6793 161 6915 170
rect 6381 -205 6390 -115
rect 6480 -205 6489 -115
rect 6631 -205 6640 -115
rect 6730 -205 6739 -115
rect 6390 -330 6480 -205
rect 6640 -309 6730 -205
rect 6793 -361 6915 41
rect 6990 -60 7330 400
rect 6990 -115 7080 -60
rect 7240 -115 7330 -60
rect 7397 161 7519 170
rect 6981 -205 6990 -115
rect 7080 -205 7089 -115
rect 7231 -205 7240 -115
rect 7330 -205 7339 -115
rect 6990 -325 7080 -205
rect 7240 -301 7330 -205
rect 7397 -361 7519 41
rect 7590 -60 7930 400
rect 7590 -115 7680 -60
rect 7840 -115 7930 -60
rect 8001 161 8123 170
rect 7581 -205 7590 -115
rect 7680 -205 7689 -115
rect 7831 -205 7840 -115
rect 7930 -205 7939 -115
rect 7590 -301 7680 -205
rect 7840 -290 7930 -205
rect 8001 -361 8123 41
rect 8200 -60 8540 400
rect 8200 -115 8290 -60
rect 8450 -115 8540 -60
rect 8605 161 8727 170
rect 8191 -205 8200 -115
rect 8290 -205 8299 -115
rect 8441 -205 8450 -115
rect 8540 -205 8549 -115
rect 8200 -290 8290 -205
rect 8450 -290 8540 -205
rect 8605 -361 8727 41
rect 8800 -60 9140 400
rect 8800 -115 8890 -60
rect 9050 -115 9140 -60
rect 9209 161 9331 170
rect 8791 -205 8800 -115
rect 8890 -205 8899 -115
rect 9041 -205 9050 -115
rect 9140 -205 9149 -115
rect 8800 -290 8890 -205
rect 9050 -304 9140 -205
rect 9209 -361 9331 41
rect 9410 -60 9750 400
rect 9410 -115 9500 -60
rect 9660 -115 9750 -60
rect 9813 161 9935 170
rect 9401 -205 9410 -115
rect 9500 -205 9509 -115
rect 9651 -205 9660 -115
rect 9750 -205 9759 -115
rect 9410 -325 9500 -205
rect 9660 -325 9750 -205
rect 9813 -361 9935 41
rect 10010 -115 10260 400
rect 10001 -205 10010 -115
rect 10100 -205 10260 -115
rect 10010 -240 10260 -205
rect 10010 -296 10100 -240
rect -840 -2220 2000 -2200
rect -840 -2280 -820 -2220
rect 1980 -2280 2000 -2220
rect -840 -2300 2000 -2280
rect 2200 -2460 4080 -2440
rect 2200 -2580 2220 -2460
rect 4060 -2580 4080 -2460
rect 2200 -2600 4080 -2580
<< via2 >>
rect 4570 -205 4660 -115
rect 4820 -205 4910 -115
rect 5180 -205 5270 -115
rect 5430 -205 5520 -115
rect 5780 -205 5870 -115
rect 6030 -205 6120 -115
rect 6390 -205 6480 -115
rect 6640 -205 6730 -115
rect 6990 -205 7080 -115
rect 7240 -205 7330 -115
rect 7590 -205 7680 -115
rect 7840 -205 7930 -115
rect 8200 -205 8290 -115
rect 8450 -205 8540 -115
rect 8800 -205 8890 -115
rect 9050 -205 9140 -115
rect 9410 -205 9500 -115
rect 9660 -205 9750 -115
rect 10010 -205 10100 -115
rect -820 -2280 1980 -2220
rect 2220 -2580 4060 -2460
<< metal3 >>
rect 4116 340 10200 460
rect 4116 -200 4156 340
rect -1000 -480 4156 -200
rect 4570 -115 4660 -106
rect 4570 -325 4660 -205
rect 4720 -480 4760 340
rect 4820 -115 4910 -106
rect 4820 -325 4910 -205
rect 5180 -115 5270 -106
rect 5180 -325 5270 -205
rect 5324 -460 5364 340
rect 5430 -115 5520 -106
rect 5430 -325 5520 -205
rect 5780 -115 5870 -106
rect 5780 -305 5870 -205
rect -1000 -1980 4140 -480
rect 5928 -500 5968 340
rect 6030 -115 6120 -106
rect 6030 -305 6120 -205
rect 6390 -115 6480 -106
rect 6390 -305 6480 -205
rect 6532 -440 6572 340
rect 6640 -115 6730 -106
rect 6640 -305 6730 -205
rect 6990 -115 7080 -106
rect 6990 -305 7080 -205
rect 7136 -500 7176 340
rect 7240 -115 7330 -106
rect 7240 -290 7330 -205
rect 7590 -115 7680 -106
rect 7590 -325 7680 -205
rect 7740 -460 7780 340
rect 7840 -115 7930 -106
rect 7840 -305 7930 -205
rect 8200 -115 8290 -106
rect 8200 -305 8290 -205
rect 8344 -420 8384 340
rect 8450 -115 8540 -106
rect 8450 -325 8540 -205
rect 8800 -115 8890 -106
rect 8800 -305 8890 -205
rect 8948 -440 8988 340
rect 9050 -115 9140 -106
rect 9050 -325 9140 -205
rect 9410 -115 9500 -106
rect 9410 -305 9500 -205
rect 9552 -440 9592 340
rect 9660 -115 9750 -106
rect 9660 -325 9750 -205
rect 10010 -115 10100 -106
rect 10010 -305 10100 -205
rect 10156 -440 10196 340
rect -1000 -2000 4160 -1980
rect -1000 -2220 2000 -2200
rect -1000 -2280 -820 -2220
rect 1980 -2280 2000 -2220
rect -1000 -6400 2000 -2280
rect 2200 -2280 4160 -2000
rect 2200 -2460 4100 -2280
rect 2200 -2580 2220 -2460
rect 4060 -2580 4100 -2460
rect 2200 -2600 4100 -2580
use sg13g2_Clamp_N20N0D  sg13g2_Clamp_N20N0D_0
timestamp 1756394914
transform -1 0 15156 0 -1 -296
box -124 -124 16124 2104
use sg13g2_Clamp_P20N0D  sg13g2_Clamp_P20N0D_0
timestamp 1756453207
transform 1 0 -844 0 1 -6334
box -56 -26 16026 3980
<< labels >>
rlabel metal1 10700 100 10700 100 0 pad
port 3 nsew
rlabel metal1 10700 340 10700 340 0 guard
port 4 nsew
rlabel metal3 -900 -1200 -900 -1200 0 VDD
port 1 nsew
rlabel metal3 -900 -4500 -900 -4500 0 VSS
port 2 nsew
<< end >>
