magic
tech ihp-sg13g2
magscale 1 2
timestamp 1756394914
<< nwell >>
rect -124 1788 16124 2104
rect -124 192 192 1788
rect 15808 192 16124 1788
rect -124 -124 16124 192
<< pwell >>
rect 334 1536 15666 1656
rect 334 464 454 1536
rect 4924 464 11076 1536
rect 15546 464 15666 1536
rect 334 344 15666 464
<< hvnmos >>
rect 5044 550 5164 1430
rect 5400 550 5520 1430
rect 5648 550 5768 1430
rect 6004 550 6124 1430
rect 6252 550 6372 1430
rect 6608 550 6728 1430
rect 6856 550 6976 1430
rect 7212 550 7332 1430
rect 7460 550 7580 1430
rect 7816 550 7936 1430
rect 8064 550 8184 1430
rect 8420 550 8540 1430
rect 8668 550 8788 1430
rect 9024 550 9144 1430
rect 9272 550 9392 1430
rect 9628 550 9748 1430
rect 9876 550 9996 1430
rect 10232 550 10352 1430
rect 10480 550 10600 1430
rect 10836 550 10956 1430
<< hvndiff >>
rect 4950 1414 5044 1430
rect 4950 1382 4964 1414
rect 4996 1382 5044 1414
rect 4950 1346 5044 1382
rect 4950 1314 4964 1346
rect 4996 1314 5044 1346
rect 4950 1278 5044 1314
rect 4950 1246 4964 1278
rect 4996 1246 5044 1278
rect 4950 1210 5044 1246
rect 4950 1178 4964 1210
rect 4996 1178 5044 1210
rect 4950 1142 5044 1178
rect 4950 1110 4964 1142
rect 4996 1110 5044 1142
rect 4950 1074 5044 1110
rect 4950 1042 4964 1074
rect 4996 1042 5044 1074
rect 4950 1006 5044 1042
rect 4950 974 4964 1006
rect 4996 974 5044 1006
rect 4950 938 5044 974
rect 4950 906 4964 938
rect 4996 906 5044 938
rect 4950 870 5044 906
rect 4950 838 4964 870
rect 4996 838 5044 870
rect 4950 802 5044 838
rect 4950 770 4964 802
rect 4996 770 5044 802
rect 4950 734 5044 770
rect 4950 702 4964 734
rect 4996 702 5044 734
rect 4950 666 5044 702
rect 4950 634 4964 666
rect 4996 634 5044 666
rect 4950 598 5044 634
rect 4950 566 4964 598
rect 4996 566 5044 598
rect 4950 550 5044 566
rect 5164 1414 5400 1430
rect 5164 1382 5266 1414
rect 5298 1382 5400 1414
rect 5164 1346 5400 1382
rect 5164 1314 5266 1346
rect 5298 1314 5400 1346
rect 5164 1278 5400 1314
rect 5164 1246 5266 1278
rect 5298 1246 5400 1278
rect 5164 1210 5400 1246
rect 5164 1178 5266 1210
rect 5298 1178 5400 1210
rect 5164 1142 5400 1178
rect 5164 1110 5266 1142
rect 5298 1110 5400 1142
rect 5164 1074 5400 1110
rect 5164 1042 5266 1074
rect 5298 1042 5400 1074
rect 5164 1006 5400 1042
rect 5164 974 5266 1006
rect 5298 974 5400 1006
rect 5164 938 5400 974
rect 5164 906 5266 938
rect 5298 906 5400 938
rect 5164 870 5400 906
rect 5164 838 5266 870
rect 5298 838 5400 870
rect 5164 802 5400 838
rect 5164 770 5266 802
rect 5298 770 5400 802
rect 5164 734 5400 770
rect 5164 702 5266 734
rect 5298 702 5400 734
rect 5164 666 5400 702
rect 5164 634 5266 666
rect 5298 634 5400 666
rect 5164 598 5400 634
rect 5164 566 5266 598
rect 5298 566 5400 598
rect 5164 550 5400 566
rect 5520 1414 5648 1430
rect 5520 1382 5568 1414
rect 5600 1382 5648 1414
rect 5520 1346 5648 1382
rect 5520 1314 5568 1346
rect 5600 1314 5648 1346
rect 5520 1278 5648 1314
rect 5520 1246 5568 1278
rect 5600 1246 5648 1278
rect 5520 1210 5648 1246
rect 5520 1178 5568 1210
rect 5600 1178 5648 1210
rect 5520 1142 5648 1178
rect 5520 1110 5568 1142
rect 5600 1110 5648 1142
rect 5520 1074 5648 1110
rect 5520 1042 5568 1074
rect 5600 1042 5648 1074
rect 5520 1006 5648 1042
rect 5520 974 5568 1006
rect 5600 974 5648 1006
rect 5520 938 5648 974
rect 5520 906 5568 938
rect 5600 906 5648 938
rect 5520 870 5648 906
rect 5520 838 5568 870
rect 5600 838 5648 870
rect 5520 802 5648 838
rect 5520 770 5568 802
rect 5600 770 5648 802
rect 5520 734 5648 770
rect 5520 702 5568 734
rect 5600 702 5648 734
rect 5520 666 5648 702
rect 5520 634 5568 666
rect 5600 634 5648 666
rect 5520 598 5648 634
rect 5520 566 5568 598
rect 5600 566 5648 598
rect 5520 550 5648 566
rect 5768 1414 6004 1430
rect 5768 1382 5870 1414
rect 5902 1382 6004 1414
rect 5768 1346 6004 1382
rect 5768 1314 5870 1346
rect 5902 1314 6004 1346
rect 5768 1278 6004 1314
rect 5768 1246 5870 1278
rect 5902 1246 6004 1278
rect 5768 1210 6004 1246
rect 5768 1178 5870 1210
rect 5902 1178 6004 1210
rect 5768 1142 6004 1178
rect 5768 1110 5870 1142
rect 5902 1110 6004 1142
rect 5768 1074 6004 1110
rect 5768 1042 5870 1074
rect 5902 1042 6004 1074
rect 5768 1006 6004 1042
rect 5768 974 5870 1006
rect 5902 974 6004 1006
rect 5768 938 6004 974
rect 5768 906 5870 938
rect 5902 906 6004 938
rect 5768 870 6004 906
rect 5768 838 5870 870
rect 5902 838 6004 870
rect 5768 802 6004 838
rect 5768 770 5870 802
rect 5902 770 6004 802
rect 5768 734 6004 770
rect 5768 702 5870 734
rect 5902 702 6004 734
rect 5768 666 6004 702
rect 5768 634 5870 666
rect 5902 634 6004 666
rect 5768 598 6004 634
rect 5768 566 5870 598
rect 5902 566 6004 598
rect 5768 550 6004 566
rect 6124 1414 6252 1430
rect 6124 1382 6172 1414
rect 6204 1382 6252 1414
rect 6124 1346 6252 1382
rect 6124 1314 6172 1346
rect 6204 1314 6252 1346
rect 6124 1278 6252 1314
rect 6124 1246 6172 1278
rect 6204 1246 6252 1278
rect 6124 1210 6252 1246
rect 6124 1178 6172 1210
rect 6204 1178 6252 1210
rect 6124 1142 6252 1178
rect 6124 1110 6172 1142
rect 6204 1110 6252 1142
rect 6124 1074 6252 1110
rect 6124 1042 6172 1074
rect 6204 1042 6252 1074
rect 6124 1006 6252 1042
rect 6124 974 6172 1006
rect 6204 974 6252 1006
rect 6124 938 6252 974
rect 6124 906 6172 938
rect 6204 906 6252 938
rect 6124 870 6252 906
rect 6124 838 6172 870
rect 6204 838 6252 870
rect 6124 802 6252 838
rect 6124 770 6172 802
rect 6204 770 6252 802
rect 6124 734 6252 770
rect 6124 702 6172 734
rect 6204 702 6252 734
rect 6124 666 6252 702
rect 6124 634 6172 666
rect 6204 634 6252 666
rect 6124 598 6252 634
rect 6124 566 6172 598
rect 6204 566 6252 598
rect 6124 550 6252 566
rect 6372 1414 6608 1430
rect 6372 1382 6474 1414
rect 6506 1382 6608 1414
rect 6372 1346 6608 1382
rect 6372 1314 6474 1346
rect 6506 1314 6608 1346
rect 6372 1278 6608 1314
rect 6372 1246 6474 1278
rect 6506 1246 6608 1278
rect 6372 1210 6608 1246
rect 6372 1178 6474 1210
rect 6506 1178 6608 1210
rect 6372 1142 6608 1178
rect 6372 1110 6474 1142
rect 6506 1110 6608 1142
rect 6372 1074 6608 1110
rect 6372 1042 6474 1074
rect 6506 1042 6608 1074
rect 6372 1006 6608 1042
rect 6372 974 6474 1006
rect 6506 974 6608 1006
rect 6372 938 6608 974
rect 6372 906 6474 938
rect 6506 906 6608 938
rect 6372 870 6608 906
rect 6372 838 6474 870
rect 6506 838 6608 870
rect 6372 802 6608 838
rect 6372 770 6474 802
rect 6506 770 6608 802
rect 6372 734 6608 770
rect 6372 702 6474 734
rect 6506 702 6608 734
rect 6372 666 6608 702
rect 6372 634 6474 666
rect 6506 634 6608 666
rect 6372 598 6608 634
rect 6372 566 6474 598
rect 6506 566 6608 598
rect 6372 550 6608 566
rect 6728 1414 6856 1430
rect 6728 1382 6776 1414
rect 6808 1382 6856 1414
rect 6728 1346 6856 1382
rect 6728 1314 6776 1346
rect 6808 1314 6856 1346
rect 6728 1278 6856 1314
rect 6728 1246 6776 1278
rect 6808 1246 6856 1278
rect 6728 1210 6856 1246
rect 6728 1178 6776 1210
rect 6808 1178 6856 1210
rect 6728 1142 6856 1178
rect 6728 1110 6776 1142
rect 6808 1110 6856 1142
rect 6728 1074 6856 1110
rect 6728 1042 6776 1074
rect 6808 1042 6856 1074
rect 6728 1006 6856 1042
rect 6728 974 6776 1006
rect 6808 974 6856 1006
rect 6728 938 6856 974
rect 6728 906 6776 938
rect 6808 906 6856 938
rect 6728 870 6856 906
rect 6728 838 6776 870
rect 6808 838 6856 870
rect 6728 802 6856 838
rect 6728 770 6776 802
rect 6808 770 6856 802
rect 6728 734 6856 770
rect 6728 702 6776 734
rect 6808 702 6856 734
rect 6728 666 6856 702
rect 6728 634 6776 666
rect 6808 634 6856 666
rect 6728 598 6856 634
rect 6728 566 6776 598
rect 6808 566 6856 598
rect 6728 550 6856 566
rect 6976 1414 7212 1430
rect 6976 1382 7078 1414
rect 7110 1382 7212 1414
rect 6976 1346 7212 1382
rect 6976 1314 7078 1346
rect 7110 1314 7212 1346
rect 6976 1278 7212 1314
rect 6976 1246 7078 1278
rect 7110 1246 7212 1278
rect 6976 1210 7212 1246
rect 6976 1178 7078 1210
rect 7110 1178 7212 1210
rect 6976 1142 7212 1178
rect 6976 1110 7078 1142
rect 7110 1110 7212 1142
rect 6976 1074 7212 1110
rect 6976 1042 7078 1074
rect 7110 1042 7212 1074
rect 6976 1006 7212 1042
rect 6976 974 7078 1006
rect 7110 974 7212 1006
rect 6976 938 7212 974
rect 6976 906 7078 938
rect 7110 906 7212 938
rect 6976 870 7212 906
rect 6976 838 7078 870
rect 7110 838 7212 870
rect 6976 802 7212 838
rect 6976 770 7078 802
rect 7110 770 7212 802
rect 6976 734 7212 770
rect 6976 702 7078 734
rect 7110 702 7212 734
rect 6976 666 7212 702
rect 6976 634 7078 666
rect 7110 634 7212 666
rect 6976 598 7212 634
rect 6976 566 7078 598
rect 7110 566 7212 598
rect 6976 550 7212 566
rect 7332 1414 7460 1430
rect 7332 1382 7380 1414
rect 7412 1382 7460 1414
rect 7332 1346 7460 1382
rect 7332 1314 7380 1346
rect 7412 1314 7460 1346
rect 7332 1278 7460 1314
rect 7332 1246 7380 1278
rect 7412 1246 7460 1278
rect 7332 1210 7460 1246
rect 7332 1178 7380 1210
rect 7412 1178 7460 1210
rect 7332 1142 7460 1178
rect 7332 1110 7380 1142
rect 7412 1110 7460 1142
rect 7332 1074 7460 1110
rect 7332 1042 7380 1074
rect 7412 1042 7460 1074
rect 7332 1006 7460 1042
rect 7332 974 7380 1006
rect 7412 974 7460 1006
rect 7332 938 7460 974
rect 7332 906 7380 938
rect 7412 906 7460 938
rect 7332 870 7460 906
rect 7332 838 7380 870
rect 7412 838 7460 870
rect 7332 802 7460 838
rect 7332 770 7380 802
rect 7412 770 7460 802
rect 7332 734 7460 770
rect 7332 702 7380 734
rect 7412 702 7460 734
rect 7332 666 7460 702
rect 7332 634 7380 666
rect 7412 634 7460 666
rect 7332 598 7460 634
rect 7332 566 7380 598
rect 7412 566 7460 598
rect 7332 550 7460 566
rect 7580 1414 7816 1430
rect 7580 1382 7682 1414
rect 7714 1382 7816 1414
rect 7580 1346 7816 1382
rect 7580 1314 7682 1346
rect 7714 1314 7816 1346
rect 7580 1278 7816 1314
rect 7580 1246 7682 1278
rect 7714 1246 7816 1278
rect 7580 1210 7816 1246
rect 7580 1178 7682 1210
rect 7714 1178 7816 1210
rect 7580 1142 7816 1178
rect 7580 1110 7682 1142
rect 7714 1110 7816 1142
rect 7580 1074 7816 1110
rect 7580 1042 7682 1074
rect 7714 1042 7816 1074
rect 7580 1006 7816 1042
rect 7580 974 7682 1006
rect 7714 974 7816 1006
rect 7580 938 7816 974
rect 7580 906 7682 938
rect 7714 906 7816 938
rect 7580 870 7816 906
rect 7580 838 7682 870
rect 7714 838 7816 870
rect 7580 802 7816 838
rect 7580 770 7682 802
rect 7714 770 7816 802
rect 7580 734 7816 770
rect 7580 702 7682 734
rect 7714 702 7816 734
rect 7580 666 7816 702
rect 7580 634 7682 666
rect 7714 634 7816 666
rect 7580 598 7816 634
rect 7580 566 7682 598
rect 7714 566 7816 598
rect 7580 550 7816 566
rect 7936 1414 8064 1430
rect 7936 1382 7984 1414
rect 8016 1382 8064 1414
rect 7936 1346 8064 1382
rect 7936 1314 7984 1346
rect 8016 1314 8064 1346
rect 7936 1278 8064 1314
rect 7936 1246 7984 1278
rect 8016 1246 8064 1278
rect 7936 1210 8064 1246
rect 7936 1178 7984 1210
rect 8016 1178 8064 1210
rect 7936 1142 8064 1178
rect 7936 1110 7984 1142
rect 8016 1110 8064 1142
rect 7936 1074 8064 1110
rect 7936 1042 7984 1074
rect 8016 1042 8064 1074
rect 7936 1006 8064 1042
rect 7936 974 7984 1006
rect 8016 974 8064 1006
rect 7936 938 8064 974
rect 7936 906 7984 938
rect 8016 906 8064 938
rect 7936 870 8064 906
rect 7936 838 7984 870
rect 8016 838 8064 870
rect 7936 802 8064 838
rect 7936 770 7984 802
rect 8016 770 8064 802
rect 7936 734 8064 770
rect 7936 702 7984 734
rect 8016 702 8064 734
rect 7936 666 8064 702
rect 7936 634 7984 666
rect 8016 634 8064 666
rect 7936 598 8064 634
rect 7936 566 7984 598
rect 8016 566 8064 598
rect 7936 550 8064 566
rect 8184 1414 8420 1430
rect 8184 1382 8286 1414
rect 8318 1382 8420 1414
rect 8184 1346 8420 1382
rect 8184 1314 8286 1346
rect 8318 1314 8420 1346
rect 8184 1278 8420 1314
rect 8184 1246 8286 1278
rect 8318 1246 8420 1278
rect 8184 1210 8420 1246
rect 8184 1178 8286 1210
rect 8318 1178 8420 1210
rect 8184 1142 8420 1178
rect 8184 1110 8286 1142
rect 8318 1110 8420 1142
rect 8184 1074 8420 1110
rect 8184 1042 8286 1074
rect 8318 1042 8420 1074
rect 8184 1006 8420 1042
rect 8184 974 8286 1006
rect 8318 974 8420 1006
rect 8184 938 8420 974
rect 8184 906 8286 938
rect 8318 906 8420 938
rect 8184 870 8420 906
rect 8184 838 8286 870
rect 8318 838 8420 870
rect 8184 802 8420 838
rect 8184 770 8286 802
rect 8318 770 8420 802
rect 8184 734 8420 770
rect 8184 702 8286 734
rect 8318 702 8420 734
rect 8184 666 8420 702
rect 8184 634 8286 666
rect 8318 634 8420 666
rect 8184 598 8420 634
rect 8184 566 8286 598
rect 8318 566 8420 598
rect 8184 550 8420 566
rect 8540 1414 8668 1430
rect 8540 1382 8588 1414
rect 8620 1382 8668 1414
rect 8540 1346 8668 1382
rect 8540 1314 8588 1346
rect 8620 1314 8668 1346
rect 8540 1278 8668 1314
rect 8540 1246 8588 1278
rect 8620 1246 8668 1278
rect 8540 1210 8668 1246
rect 8540 1178 8588 1210
rect 8620 1178 8668 1210
rect 8540 1142 8668 1178
rect 8540 1110 8588 1142
rect 8620 1110 8668 1142
rect 8540 1074 8668 1110
rect 8540 1042 8588 1074
rect 8620 1042 8668 1074
rect 8540 1006 8668 1042
rect 8540 974 8588 1006
rect 8620 974 8668 1006
rect 8540 938 8668 974
rect 8540 906 8588 938
rect 8620 906 8668 938
rect 8540 870 8668 906
rect 8540 838 8588 870
rect 8620 838 8668 870
rect 8540 802 8668 838
rect 8540 770 8588 802
rect 8620 770 8668 802
rect 8540 734 8668 770
rect 8540 702 8588 734
rect 8620 702 8668 734
rect 8540 666 8668 702
rect 8540 634 8588 666
rect 8620 634 8668 666
rect 8540 598 8668 634
rect 8540 566 8588 598
rect 8620 566 8668 598
rect 8540 550 8668 566
rect 8788 1414 9024 1430
rect 8788 1382 8890 1414
rect 8922 1382 9024 1414
rect 8788 1346 9024 1382
rect 8788 1314 8890 1346
rect 8922 1314 9024 1346
rect 8788 1278 9024 1314
rect 8788 1246 8890 1278
rect 8922 1246 9024 1278
rect 8788 1210 9024 1246
rect 8788 1178 8890 1210
rect 8922 1178 9024 1210
rect 8788 1142 9024 1178
rect 8788 1110 8890 1142
rect 8922 1110 9024 1142
rect 8788 1074 9024 1110
rect 8788 1042 8890 1074
rect 8922 1042 9024 1074
rect 8788 1006 9024 1042
rect 8788 974 8890 1006
rect 8922 974 9024 1006
rect 8788 938 9024 974
rect 8788 906 8890 938
rect 8922 906 9024 938
rect 8788 870 9024 906
rect 8788 838 8890 870
rect 8922 838 9024 870
rect 8788 802 9024 838
rect 8788 770 8890 802
rect 8922 770 9024 802
rect 8788 734 9024 770
rect 8788 702 8890 734
rect 8922 702 9024 734
rect 8788 666 9024 702
rect 8788 634 8890 666
rect 8922 634 9024 666
rect 8788 598 9024 634
rect 8788 566 8890 598
rect 8922 566 9024 598
rect 8788 550 9024 566
rect 9144 1414 9272 1430
rect 9144 1382 9192 1414
rect 9224 1382 9272 1414
rect 9144 1346 9272 1382
rect 9144 1314 9192 1346
rect 9224 1314 9272 1346
rect 9144 1278 9272 1314
rect 9144 1246 9192 1278
rect 9224 1246 9272 1278
rect 9144 1210 9272 1246
rect 9144 1178 9192 1210
rect 9224 1178 9272 1210
rect 9144 1142 9272 1178
rect 9144 1110 9192 1142
rect 9224 1110 9272 1142
rect 9144 1074 9272 1110
rect 9144 1042 9192 1074
rect 9224 1042 9272 1074
rect 9144 1006 9272 1042
rect 9144 974 9192 1006
rect 9224 974 9272 1006
rect 9144 938 9272 974
rect 9144 906 9192 938
rect 9224 906 9272 938
rect 9144 870 9272 906
rect 9144 838 9192 870
rect 9224 838 9272 870
rect 9144 802 9272 838
rect 9144 770 9192 802
rect 9224 770 9272 802
rect 9144 734 9272 770
rect 9144 702 9192 734
rect 9224 702 9272 734
rect 9144 666 9272 702
rect 9144 634 9192 666
rect 9224 634 9272 666
rect 9144 598 9272 634
rect 9144 566 9192 598
rect 9224 566 9272 598
rect 9144 550 9272 566
rect 9392 1414 9628 1430
rect 9392 1382 9494 1414
rect 9526 1382 9628 1414
rect 9392 1346 9628 1382
rect 9392 1314 9494 1346
rect 9526 1314 9628 1346
rect 9392 1278 9628 1314
rect 9392 1246 9494 1278
rect 9526 1246 9628 1278
rect 9392 1210 9628 1246
rect 9392 1178 9494 1210
rect 9526 1178 9628 1210
rect 9392 1142 9628 1178
rect 9392 1110 9494 1142
rect 9526 1110 9628 1142
rect 9392 1074 9628 1110
rect 9392 1042 9494 1074
rect 9526 1042 9628 1074
rect 9392 1006 9628 1042
rect 9392 974 9494 1006
rect 9526 974 9628 1006
rect 9392 938 9628 974
rect 9392 906 9494 938
rect 9526 906 9628 938
rect 9392 870 9628 906
rect 9392 838 9494 870
rect 9526 838 9628 870
rect 9392 802 9628 838
rect 9392 770 9494 802
rect 9526 770 9628 802
rect 9392 734 9628 770
rect 9392 702 9494 734
rect 9526 702 9628 734
rect 9392 666 9628 702
rect 9392 634 9494 666
rect 9526 634 9628 666
rect 9392 598 9628 634
rect 9392 566 9494 598
rect 9526 566 9628 598
rect 9392 550 9628 566
rect 9748 1414 9876 1430
rect 9748 1382 9796 1414
rect 9828 1382 9876 1414
rect 9748 1346 9876 1382
rect 9748 1314 9796 1346
rect 9828 1314 9876 1346
rect 9748 1278 9876 1314
rect 9748 1246 9796 1278
rect 9828 1246 9876 1278
rect 9748 1210 9876 1246
rect 9748 1178 9796 1210
rect 9828 1178 9876 1210
rect 9748 1142 9876 1178
rect 9748 1110 9796 1142
rect 9828 1110 9876 1142
rect 9748 1074 9876 1110
rect 9748 1042 9796 1074
rect 9828 1042 9876 1074
rect 9748 1006 9876 1042
rect 9748 974 9796 1006
rect 9828 974 9876 1006
rect 9748 938 9876 974
rect 9748 906 9796 938
rect 9828 906 9876 938
rect 9748 870 9876 906
rect 9748 838 9796 870
rect 9828 838 9876 870
rect 9748 802 9876 838
rect 9748 770 9796 802
rect 9828 770 9876 802
rect 9748 734 9876 770
rect 9748 702 9796 734
rect 9828 702 9876 734
rect 9748 666 9876 702
rect 9748 634 9796 666
rect 9828 634 9876 666
rect 9748 598 9876 634
rect 9748 566 9796 598
rect 9828 566 9876 598
rect 9748 550 9876 566
rect 9996 1414 10232 1430
rect 9996 1382 10098 1414
rect 10130 1382 10232 1414
rect 9996 1346 10232 1382
rect 9996 1314 10098 1346
rect 10130 1314 10232 1346
rect 9996 1278 10232 1314
rect 9996 1246 10098 1278
rect 10130 1246 10232 1278
rect 9996 1210 10232 1246
rect 9996 1178 10098 1210
rect 10130 1178 10232 1210
rect 9996 1142 10232 1178
rect 9996 1110 10098 1142
rect 10130 1110 10232 1142
rect 9996 1074 10232 1110
rect 9996 1042 10098 1074
rect 10130 1042 10232 1074
rect 9996 1006 10232 1042
rect 9996 974 10098 1006
rect 10130 974 10232 1006
rect 9996 938 10232 974
rect 9996 906 10098 938
rect 10130 906 10232 938
rect 9996 870 10232 906
rect 9996 838 10098 870
rect 10130 838 10232 870
rect 9996 802 10232 838
rect 9996 770 10098 802
rect 10130 770 10232 802
rect 9996 734 10232 770
rect 9996 702 10098 734
rect 10130 702 10232 734
rect 9996 666 10232 702
rect 9996 634 10098 666
rect 10130 634 10232 666
rect 9996 598 10232 634
rect 9996 566 10098 598
rect 10130 566 10232 598
rect 9996 550 10232 566
rect 10352 1414 10480 1430
rect 10352 1382 10400 1414
rect 10432 1382 10480 1414
rect 10352 1346 10480 1382
rect 10352 1314 10400 1346
rect 10432 1314 10480 1346
rect 10352 1278 10480 1314
rect 10352 1246 10400 1278
rect 10432 1246 10480 1278
rect 10352 1210 10480 1246
rect 10352 1178 10400 1210
rect 10432 1178 10480 1210
rect 10352 1142 10480 1178
rect 10352 1110 10400 1142
rect 10432 1110 10480 1142
rect 10352 1074 10480 1110
rect 10352 1042 10400 1074
rect 10432 1042 10480 1074
rect 10352 1006 10480 1042
rect 10352 974 10400 1006
rect 10432 974 10480 1006
rect 10352 938 10480 974
rect 10352 906 10400 938
rect 10432 906 10480 938
rect 10352 870 10480 906
rect 10352 838 10400 870
rect 10432 838 10480 870
rect 10352 802 10480 838
rect 10352 770 10400 802
rect 10432 770 10480 802
rect 10352 734 10480 770
rect 10352 702 10400 734
rect 10432 702 10480 734
rect 10352 666 10480 702
rect 10352 634 10400 666
rect 10432 634 10480 666
rect 10352 598 10480 634
rect 10352 566 10400 598
rect 10432 566 10480 598
rect 10352 550 10480 566
rect 10600 1414 10836 1430
rect 10600 1382 10702 1414
rect 10734 1382 10836 1414
rect 10600 1346 10836 1382
rect 10600 1314 10702 1346
rect 10734 1314 10836 1346
rect 10600 1278 10836 1314
rect 10600 1246 10702 1278
rect 10734 1246 10836 1278
rect 10600 1210 10836 1246
rect 10600 1178 10702 1210
rect 10734 1178 10836 1210
rect 10600 1142 10836 1178
rect 10600 1110 10702 1142
rect 10734 1110 10836 1142
rect 10600 1074 10836 1110
rect 10600 1042 10702 1074
rect 10734 1042 10836 1074
rect 10600 1006 10836 1042
rect 10600 974 10702 1006
rect 10734 974 10836 1006
rect 10600 938 10836 974
rect 10600 906 10702 938
rect 10734 906 10836 938
rect 10600 870 10836 906
rect 10600 838 10702 870
rect 10734 838 10836 870
rect 10600 802 10836 838
rect 10600 770 10702 802
rect 10734 770 10836 802
rect 10600 734 10836 770
rect 10600 702 10702 734
rect 10734 702 10836 734
rect 10600 666 10836 702
rect 10600 634 10702 666
rect 10734 634 10836 666
rect 10600 598 10836 634
rect 10600 566 10702 598
rect 10734 566 10836 598
rect 10600 550 10836 566
rect 10956 1414 11050 1430
rect 10956 1382 11004 1414
rect 11036 1382 11050 1414
rect 10956 1346 11050 1382
rect 10956 1314 11004 1346
rect 11036 1314 11050 1346
rect 10956 1278 11050 1314
rect 10956 1246 11004 1278
rect 11036 1246 11050 1278
rect 10956 1210 11050 1246
rect 10956 1178 11004 1210
rect 11036 1178 11050 1210
rect 10956 1142 11050 1178
rect 10956 1110 11004 1142
rect 11036 1110 11050 1142
rect 10956 1074 11050 1110
rect 10956 1042 11004 1074
rect 11036 1042 11050 1074
rect 10956 1006 11050 1042
rect 10956 974 11004 1006
rect 11036 974 11050 1006
rect 10956 938 11050 974
rect 10956 906 11004 938
rect 11036 906 11050 938
rect 10956 870 11050 906
rect 10956 838 11004 870
rect 11036 838 11050 870
rect 10956 802 11050 838
rect 10956 770 11004 802
rect 11036 770 11050 802
rect 10956 734 11050 770
rect 10956 702 11004 734
rect 11036 702 11050 734
rect 10956 666 11050 702
rect 10956 634 11004 666
rect 11036 634 11050 666
rect 10956 598 11050 634
rect 10956 566 11004 598
rect 11036 566 11050 598
rect 10956 550 11050 566
<< hvndiffc >>
rect 4964 1382 4996 1414
rect 4964 1314 4996 1346
rect 4964 1246 4996 1278
rect 4964 1178 4996 1210
rect 4964 1110 4996 1142
rect 4964 1042 4996 1074
rect 4964 974 4996 1006
rect 4964 906 4996 938
rect 4964 838 4996 870
rect 4964 770 4996 802
rect 4964 702 4996 734
rect 4964 634 4996 666
rect 4964 566 4996 598
rect 5266 1382 5298 1414
rect 5266 1314 5298 1346
rect 5266 1246 5298 1278
rect 5266 1178 5298 1210
rect 5266 1110 5298 1142
rect 5266 1042 5298 1074
rect 5266 974 5298 1006
rect 5266 906 5298 938
rect 5266 838 5298 870
rect 5266 770 5298 802
rect 5266 702 5298 734
rect 5266 634 5298 666
rect 5266 566 5298 598
rect 5568 1382 5600 1414
rect 5568 1314 5600 1346
rect 5568 1246 5600 1278
rect 5568 1178 5600 1210
rect 5568 1110 5600 1142
rect 5568 1042 5600 1074
rect 5568 974 5600 1006
rect 5568 906 5600 938
rect 5568 838 5600 870
rect 5568 770 5600 802
rect 5568 702 5600 734
rect 5568 634 5600 666
rect 5568 566 5600 598
rect 5870 1382 5902 1414
rect 5870 1314 5902 1346
rect 5870 1246 5902 1278
rect 5870 1178 5902 1210
rect 5870 1110 5902 1142
rect 5870 1042 5902 1074
rect 5870 974 5902 1006
rect 5870 906 5902 938
rect 5870 838 5902 870
rect 5870 770 5902 802
rect 5870 702 5902 734
rect 5870 634 5902 666
rect 5870 566 5902 598
rect 6172 1382 6204 1414
rect 6172 1314 6204 1346
rect 6172 1246 6204 1278
rect 6172 1178 6204 1210
rect 6172 1110 6204 1142
rect 6172 1042 6204 1074
rect 6172 974 6204 1006
rect 6172 906 6204 938
rect 6172 838 6204 870
rect 6172 770 6204 802
rect 6172 702 6204 734
rect 6172 634 6204 666
rect 6172 566 6204 598
rect 6474 1382 6506 1414
rect 6474 1314 6506 1346
rect 6474 1246 6506 1278
rect 6474 1178 6506 1210
rect 6474 1110 6506 1142
rect 6474 1042 6506 1074
rect 6474 974 6506 1006
rect 6474 906 6506 938
rect 6474 838 6506 870
rect 6474 770 6506 802
rect 6474 702 6506 734
rect 6474 634 6506 666
rect 6474 566 6506 598
rect 6776 1382 6808 1414
rect 6776 1314 6808 1346
rect 6776 1246 6808 1278
rect 6776 1178 6808 1210
rect 6776 1110 6808 1142
rect 6776 1042 6808 1074
rect 6776 974 6808 1006
rect 6776 906 6808 938
rect 6776 838 6808 870
rect 6776 770 6808 802
rect 6776 702 6808 734
rect 6776 634 6808 666
rect 6776 566 6808 598
rect 7078 1382 7110 1414
rect 7078 1314 7110 1346
rect 7078 1246 7110 1278
rect 7078 1178 7110 1210
rect 7078 1110 7110 1142
rect 7078 1042 7110 1074
rect 7078 974 7110 1006
rect 7078 906 7110 938
rect 7078 838 7110 870
rect 7078 770 7110 802
rect 7078 702 7110 734
rect 7078 634 7110 666
rect 7078 566 7110 598
rect 7380 1382 7412 1414
rect 7380 1314 7412 1346
rect 7380 1246 7412 1278
rect 7380 1178 7412 1210
rect 7380 1110 7412 1142
rect 7380 1042 7412 1074
rect 7380 974 7412 1006
rect 7380 906 7412 938
rect 7380 838 7412 870
rect 7380 770 7412 802
rect 7380 702 7412 734
rect 7380 634 7412 666
rect 7380 566 7412 598
rect 7682 1382 7714 1414
rect 7682 1314 7714 1346
rect 7682 1246 7714 1278
rect 7682 1178 7714 1210
rect 7682 1110 7714 1142
rect 7682 1042 7714 1074
rect 7682 974 7714 1006
rect 7682 906 7714 938
rect 7682 838 7714 870
rect 7682 770 7714 802
rect 7682 702 7714 734
rect 7682 634 7714 666
rect 7682 566 7714 598
rect 7984 1382 8016 1414
rect 7984 1314 8016 1346
rect 7984 1246 8016 1278
rect 7984 1178 8016 1210
rect 7984 1110 8016 1142
rect 7984 1042 8016 1074
rect 7984 974 8016 1006
rect 7984 906 8016 938
rect 7984 838 8016 870
rect 7984 770 8016 802
rect 7984 702 8016 734
rect 7984 634 8016 666
rect 7984 566 8016 598
rect 8286 1382 8318 1414
rect 8286 1314 8318 1346
rect 8286 1246 8318 1278
rect 8286 1178 8318 1210
rect 8286 1110 8318 1142
rect 8286 1042 8318 1074
rect 8286 974 8318 1006
rect 8286 906 8318 938
rect 8286 838 8318 870
rect 8286 770 8318 802
rect 8286 702 8318 734
rect 8286 634 8318 666
rect 8286 566 8318 598
rect 8588 1382 8620 1414
rect 8588 1314 8620 1346
rect 8588 1246 8620 1278
rect 8588 1178 8620 1210
rect 8588 1110 8620 1142
rect 8588 1042 8620 1074
rect 8588 974 8620 1006
rect 8588 906 8620 938
rect 8588 838 8620 870
rect 8588 770 8620 802
rect 8588 702 8620 734
rect 8588 634 8620 666
rect 8588 566 8620 598
rect 8890 1382 8922 1414
rect 8890 1314 8922 1346
rect 8890 1246 8922 1278
rect 8890 1178 8922 1210
rect 8890 1110 8922 1142
rect 8890 1042 8922 1074
rect 8890 974 8922 1006
rect 8890 906 8922 938
rect 8890 838 8922 870
rect 8890 770 8922 802
rect 8890 702 8922 734
rect 8890 634 8922 666
rect 8890 566 8922 598
rect 9192 1382 9224 1414
rect 9192 1314 9224 1346
rect 9192 1246 9224 1278
rect 9192 1178 9224 1210
rect 9192 1110 9224 1142
rect 9192 1042 9224 1074
rect 9192 974 9224 1006
rect 9192 906 9224 938
rect 9192 838 9224 870
rect 9192 770 9224 802
rect 9192 702 9224 734
rect 9192 634 9224 666
rect 9192 566 9224 598
rect 9494 1382 9526 1414
rect 9494 1314 9526 1346
rect 9494 1246 9526 1278
rect 9494 1178 9526 1210
rect 9494 1110 9526 1142
rect 9494 1042 9526 1074
rect 9494 974 9526 1006
rect 9494 906 9526 938
rect 9494 838 9526 870
rect 9494 770 9526 802
rect 9494 702 9526 734
rect 9494 634 9526 666
rect 9494 566 9526 598
rect 9796 1382 9828 1414
rect 9796 1314 9828 1346
rect 9796 1246 9828 1278
rect 9796 1178 9828 1210
rect 9796 1110 9828 1142
rect 9796 1042 9828 1074
rect 9796 974 9828 1006
rect 9796 906 9828 938
rect 9796 838 9828 870
rect 9796 770 9828 802
rect 9796 702 9828 734
rect 9796 634 9828 666
rect 9796 566 9828 598
rect 10098 1382 10130 1414
rect 10098 1314 10130 1346
rect 10098 1246 10130 1278
rect 10098 1178 10130 1210
rect 10098 1110 10130 1142
rect 10098 1042 10130 1074
rect 10098 974 10130 1006
rect 10098 906 10130 938
rect 10098 838 10130 870
rect 10098 770 10130 802
rect 10098 702 10130 734
rect 10098 634 10130 666
rect 10098 566 10130 598
rect 10400 1382 10432 1414
rect 10400 1314 10432 1346
rect 10400 1246 10432 1278
rect 10400 1178 10432 1210
rect 10400 1110 10432 1142
rect 10400 1042 10432 1074
rect 10400 974 10432 1006
rect 10400 906 10432 938
rect 10400 838 10432 870
rect 10400 770 10432 802
rect 10400 702 10432 734
rect 10400 634 10432 666
rect 10400 566 10432 598
rect 10702 1382 10734 1414
rect 10702 1314 10734 1346
rect 10702 1246 10734 1278
rect 10702 1178 10734 1210
rect 10702 1110 10734 1142
rect 10702 1042 10734 1074
rect 10702 974 10734 1006
rect 10702 906 10734 938
rect 10702 838 10734 870
rect 10702 770 10734 802
rect 10702 702 10734 734
rect 10702 634 10734 666
rect 10702 566 10734 598
rect 11004 1382 11036 1414
rect 11004 1314 11036 1346
rect 11004 1246 11036 1278
rect 11004 1178 11036 1210
rect 11004 1110 11036 1142
rect 11004 1042 11036 1074
rect 11004 974 11036 1006
rect 11004 906 11036 938
rect 11004 838 11036 870
rect 11004 770 11036 802
rect 11004 702 11036 734
rect 11004 634 11036 666
rect 11004 566 11036 598
<< psubdiff >>
rect 360 1612 15640 1630
rect 360 1580 402 1612
rect 434 1580 470 1612
rect 502 1580 538 1612
rect 570 1580 606 1612
rect 638 1580 674 1612
rect 706 1580 742 1612
rect 774 1580 810 1612
rect 842 1580 878 1612
rect 910 1580 946 1612
rect 978 1580 1014 1612
rect 1046 1580 1082 1612
rect 1114 1580 1150 1612
rect 1182 1580 1218 1612
rect 1250 1580 1286 1612
rect 1318 1580 1354 1612
rect 1386 1580 1422 1612
rect 1454 1580 1490 1612
rect 1522 1580 1558 1612
rect 1590 1580 1626 1612
rect 1658 1580 1694 1612
rect 1726 1580 1762 1612
rect 1794 1580 1830 1612
rect 1862 1580 1898 1612
rect 1930 1580 1966 1612
rect 1998 1580 2034 1612
rect 2066 1580 2102 1612
rect 2134 1580 2170 1612
rect 2202 1580 2238 1612
rect 2270 1580 2306 1612
rect 2338 1580 2374 1612
rect 2406 1580 2442 1612
rect 2474 1580 2510 1612
rect 2542 1580 2578 1612
rect 2610 1580 2646 1612
rect 2678 1580 2714 1612
rect 2746 1580 2782 1612
rect 2814 1580 2850 1612
rect 2882 1580 2918 1612
rect 2950 1580 2986 1612
rect 3018 1580 3054 1612
rect 3086 1580 3122 1612
rect 3154 1580 3190 1612
rect 3222 1580 3258 1612
rect 3290 1580 3326 1612
rect 3358 1580 3394 1612
rect 3426 1580 3462 1612
rect 3494 1580 3530 1612
rect 3562 1580 3598 1612
rect 3630 1580 3666 1612
rect 3698 1580 3734 1612
rect 3766 1580 3802 1612
rect 3834 1580 3870 1612
rect 3902 1580 3938 1612
rect 3970 1580 4006 1612
rect 4038 1580 4074 1612
rect 4106 1580 4142 1612
rect 4174 1580 4210 1612
rect 4242 1580 4278 1612
rect 4310 1580 4346 1612
rect 4378 1580 4414 1612
rect 4446 1580 4482 1612
rect 4514 1580 4550 1612
rect 4582 1580 4618 1612
rect 4650 1580 4686 1612
rect 4718 1580 4754 1612
rect 4786 1580 4822 1612
rect 4854 1580 4890 1612
rect 4922 1580 4958 1612
rect 4990 1580 5026 1612
rect 5058 1580 5094 1612
rect 5126 1580 5162 1612
rect 5194 1580 5230 1612
rect 5262 1580 5298 1612
rect 5330 1580 5366 1612
rect 5398 1580 5434 1612
rect 5466 1580 5502 1612
rect 5534 1580 5570 1612
rect 5602 1580 5638 1612
rect 5670 1580 5706 1612
rect 5738 1580 5774 1612
rect 5806 1580 5842 1612
rect 5874 1580 5910 1612
rect 5942 1580 5978 1612
rect 6010 1580 6046 1612
rect 6078 1580 6114 1612
rect 6146 1580 6182 1612
rect 6214 1580 6250 1612
rect 6282 1580 6318 1612
rect 6350 1580 6386 1612
rect 6418 1580 6454 1612
rect 6486 1580 6522 1612
rect 6554 1580 6590 1612
rect 6622 1580 6658 1612
rect 6690 1580 6726 1612
rect 6758 1580 6794 1612
rect 6826 1580 6862 1612
rect 6894 1580 6930 1612
rect 6962 1580 6998 1612
rect 7030 1580 7066 1612
rect 7098 1580 7134 1612
rect 7166 1580 7202 1612
rect 7234 1580 7270 1612
rect 7302 1580 7338 1612
rect 7370 1580 7406 1612
rect 7438 1580 7474 1612
rect 7506 1580 7542 1612
rect 7574 1580 7610 1612
rect 7642 1580 7678 1612
rect 7710 1580 7746 1612
rect 7778 1580 7814 1612
rect 7846 1580 7882 1612
rect 7914 1580 7950 1612
rect 7982 1580 8018 1612
rect 8050 1580 8086 1612
rect 8118 1580 8154 1612
rect 8186 1580 8222 1612
rect 8254 1580 8290 1612
rect 8322 1580 8358 1612
rect 8390 1580 8426 1612
rect 8458 1580 8494 1612
rect 8526 1580 8562 1612
rect 8594 1580 8630 1612
rect 8662 1580 8698 1612
rect 8730 1580 8766 1612
rect 8798 1580 8834 1612
rect 8866 1580 8902 1612
rect 8934 1580 8970 1612
rect 9002 1580 9038 1612
rect 9070 1580 9106 1612
rect 9138 1580 9174 1612
rect 9206 1580 9242 1612
rect 9274 1580 9310 1612
rect 9342 1580 9378 1612
rect 9410 1580 9446 1612
rect 9478 1580 9514 1612
rect 9546 1580 9582 1612
rect 9614 1580 9650 1612
rect 9682 1580 9718 1612
rect 9750 1580 9786 1612
rect 9818 1580 9854 1612
rect 9886 1580 9922 1612
rect 9954 1580 9990 1612
rect 10022 1580 10058 1612
rect 10090 1580 10126 1612
rect 10158 1580 10194 1612
rect 10226 1580 10262 1612
rect 10294 1580 10330 1612
rect 10362 1580 10398 1612
rect 10430 1580 10466 1612
rect 10498 1580 10534 1612
rect 10566 1580 10602 1612
rect 10634 1580 10670 1612
rect 10702 1580 10738 1612
rect 10770 1580 10806 1612
rect 10838 1580 10874 1612
rect 10906 1580 10942 1612
rect 10974 1580 11010 1612
rect 11042 1580 11078 1612
rect 11110 1580 11146 1612
rect 11178 1580 11214 1612
rect 11246 1580 11282 1612
rect 11314 1580 11350 1612
rect 11382 1580 11418 1612
rect 11450 1580 11486 1612
rect 11518 1580 11554 1612
rect 11586 1580 11622 1612
rect 11654 1580 11690 1612
rect 11722 1580 11758 1612
rect 11790 1580 11826 1612
rect 11858 1580 11894 1612
rect 11926 1580 11962 1612
rect 11994 1580 12030 1612
rect 12062 1580 12098 1612
rect 12130 1580 12166 1612
rect 12198 1580 12234 1612
rect 12266 1580 12302 1612
rect 12334 1580 12370 1612
rect 12402 1580 12438 1612
rect 12470 1580 12506 1612
rect 12538 1580 12574 1612
rect 12606 1580 12642 1612
rect 12674 1580 12710 1612
rect 12742 1580 12778 1612
rect 12810 1580 12846 1612
rect 12878 1580 12914 1612
rect 12946 1580 12982 1612
rect 13014 1580 13050 1612
rect 13082 1580 13118 1612
rect 13150 1580 13186 1612
rect 13218 1580 13254 1612
rect 13286 1580 13322 1612
rect 13354 1580 13390 1612
rect 13422 1580 13458 1612
rect 13490 1580 13526 1612
rect 13558 1580 13594 1612
rect 13626 1580 13662 1612
rect 13694 1580 13730 1612
rect 13762 1580 13798 1612
rect 13830 1580 13866 1612
rect 13898 1580 13934 1612
rect 13966 1580 14002 1612
rect 14034 1580 14070 1612
rect 14102 1580 14138 1612
rect 14170 1580 14206 1612
rect 14238 1580 14274 1612
rect 14306 1580 14342 1612
rect 14374 1580 14410 1612
rect 14442 1580 14478 1612
rect 14510 1580 14546 1612
rect 14578 1580 14614 1612
rect 14646 1580 14682 1612
rect 14714 1580 14750 1612
rect 14782 1580 14818 1612
rect 14850 1580 14886 1612
rect 14918 1580 14954 1612
rect 14986 1580 15022 1612
rect 15054 1580 15090 1612
rect 15122 1580 15158 1612
rect 15190 1580 15226 1612
rect 15258 1580 15294 1612
rect 15326 1580 15362 1612
rect 15394 1580 15430 1612
rect 15462 1580 15498 1612
rect 15530 1580 15566 1612
rect 15598 1580 15640 1612
rect 360 1562 15640 1580
rect 360 1526 428 1562
rect 360 1494 378 1526
rect 410 1494 428 1526
rect 15572 1526 15640 1562
rect 360 1458 428 1494
rect 360 1426 378 1458
rect 410 1426 428 1458
rect 15572 1494 15590 1526
rect 15622 1494 15640 1526
rect 15572 1458 15640 1494
rect 360 1390 428 1426
rect 360 1358 378 1390
rect 410 1358 428 1390
rect 360 1322 428 1358
rect 360 1290 378 1322
rect 410 1290 428 1322
rect 360 1254 428 1290
rect 360 1222 378 1254
rect 410 1222 428 1254
rect 360 1186 428 1222
rect 360 1154 378 1186
rect 410 1154 428 1186
rect 360 1118 428 1154
rect 360 1086 378 1118
rect 410 1086 428 1118
rect 360 1050 428 1086
rect 360 1018 378 1050
rect 410 1018 428 1050
rect 360 982 428 1018
rect 360 950 378 982
rect 410 950 428 982
rect 360 914 428 950
rect 360 882 378 914
rect 410 882 428 914
rect 360 846 428 882
rect 360 814 378 846
rect 410 814 428 846
rect 360 778 428 814
rect 360 746 378 778
rect 410 746 428 778
rect 360 710 428 746
rect 360 678 378 710
rect 410 678 428 710
rect 360 642 428 678
rect 360 610 378 642
rect 410 610 428 642
rect 360 574 428 610
rect 360 542 378 574
rect 410 542 428 574
rect 15572 1426 15590 1458
rect 15622 1426 15640 1458
rect 15572 1390 15640 1426
rect 15572 1358 15590 1390
rect 15622 1358 15640 1390
rect 15572 1322 15640 1358
rect 15572 1290 15590 1322
rect 15622 1290 15640 1322
rect 15572 1254 15640 1290
rect 15572 1222 15590 1254
rect 15622 1222 15640 1254
rect 15572 1186 15640 1222
rect 15572 1154 15590 1186
rect 15622 1154 15640 1186
rect 15572 1118 15640 1154
rect 15572 1086 15590 1118
rect 15622 1086 15640 1118
rect 15572 1050 15640 1086
rect 15572 1018 15590 1050
rect 15622 1018 15640 1050
rect 15572 982 15640 1018
rect 15572 950 15590 982
rect 15622 950 15640 982
rect 15572 914 15640 950
rect 15572 882 15590 914
rect 15622 882 15640 914
rect 15572 846 15640 882
rect 15572 814 15590 846
rect 15622 814 15640 846
rect 15572 778 15640 814
rect 15572 746 15590 778
rect 15622 746 15640 778
rect 15572 710 15640 746
rect 15572 678 15590 710
rect 15622 678 15640 710
rect 15572 642 15640 678
rect 15572 610 15590 642
rect 15622 610 15640 642
rect 15572 574 15640 610
rect 360 506 428 542
rect 360 474 378 506
rect 410 474 428 506
rect 15572 542 15590 574
rect 15622 542 15640 574
rect 15572 506 15640 542
rect 360 438 428 474
rect 15572 474 15590 506
rect 15622 474 15640 506
rect 15572 438 15640 474
rect 360 420 15640 438
rect 360 388 402 420
rect 434 388 470 420
rect 502 388 538 420
rect 570 388 606 420
rect 638 388 674 420
rect 706 388 742 420
rect 774 388 810 420
rect 842 388 878 420
rect 910 388 946 420
rect 978 388 1014 420
rect 1046 388 1082 420
rect 1114 388 1150 420
rect 1182 388 1218 420
rect 1250 388 1286 420
rect 1318 388 1354 420
rect 1386 388 1422 420
rect 1454 388 1490 420
rect 1522 388 1558 420
rect 1590 388 1626 420
rect 1658 388 1694 420
rect 1726 388 1762 420
rect 1794 388 1830 420
rect 1862 388 1898 420
rect 1930 388 1966 420
rect 1998 388 2034 420
rect 2066 388 2102 420
rect 2134 388 2170 420
rect 2202 388 2238 420
rect 2270 388 2306 420
rect 2338 388 2374 420
rect 2406 388 2442 420
rect 2474 388 2510 420
rect 2542 388 2578 420
rect 2610 388 2646 420
rect 2678 388 2714 420
rect 2746 388 2782 420
rect 2814 388 2850 420
rect 2882 388 2918 420
rect 2950 388 2986 420
rect 3018 388 3054 420
rect 3086 388 3122 420
rect 3154 388 3190 420
rect 3222 388 3258 420
rect 3290 388 3326 420
rect 3358 388 3394 420
rect 3426 388 3462 420
rect 3494 388 3530 420
rect 3562 388 3598 420
rect 3630 388 3666 420
rect 3698 388 3734 420
rect 3766 388 3802 420
rect 3834 388 3870 420
rect 3902 388 3938 420
rect 3970 388 4006 420
rect 4038 388 4074 420
rect 4106 388 4142 420
rect 4174 388 4210 420
rect 4242 388 4278 420
rect 4310 388 4346 420
rect 4378 388 4414 420
rect 4446 388 4482 420
rect 4514 388 4550 420
rect 4582 388 4618 420
rect 4650 388 4686 420
rect 4718 388 4754 420
rect 4786 388 4822 420
rect 4854 388 4890 420
rect 4922 388 4958 420
rect 4990 388 5026 420
rect 5058 388 5094 420
rect 5126 388 5162 420
rect 5194 388 5230 420
rect 5262 388 5298 420
rect 5330 388 5366 420
rect 5398 388 5434 420
rect 5466 388 5502 420
rect 5534 388 5570 420
rect 5602 388 5638 420
rect 5670 388 5706 420
rect 5738 388 5774 420
rect 5806 388 5842 420
rect 5874 388 5910 420
rect 5942 388 5978 420
rect 6010 388 6046 420
rect 6078 388 6114 420
rect 6146 388 6182 420
rect 6214 388 6250 420
rect 6282 388 6318 420
rect 6350 388 6386 420
rect 6418 388 6454 420
rect 6486 388 6522 420
rect 6554 388 6590 420
rect 6622 388 6658 420
rect 6690 388 6726 420
rect 6758 388 6794 420
rect 6826 388 6862 420
rect 6894 388 6930 420
rect 6962 388 6998 420
rect 7030 388 7066 420
rect 7098 388 7134 420
rect 7166 388 7202 420
rect 7234 388 7270 420
rect 7302 388 7338 420
rect 7370 388 7406 420
rect 7438 388 7474 420
rect 7506 388 7542 420
rect 7574 388 7610 420
rect 7642 388 7678 420
rect 7710 388 7746 420
rect 7778 388 7814 420
rect 7846 388 7882 420
rect 7914 388 7950 420
rect 7982 388 8018 420
rect 8050 388 8086 420
rect 8118 388 8154 420
rect 8186 388 8222 420
rect 8254 388 8290 420
rect 8322 388 8358 420
rect 8390 388 8426 420
rect 8458 388 8494 420
rect 8526 388 8562 420
rect 8594 388 8630 420
rect 8662 388 8698 420
rect 8730 388 8766 420
rect 8798 388 8834 420
rect 8866 388 8902 420
rect 8934 388 8970 420
rect 9002 388 9038 420
rect 9070 388 9106 420
rect 9138 388 9174 420
rect 9206 388 9242 420
rect 9274 388 9310 420
rect 9342 388 9378 420
rect 9410 388 9446 420
rect 9478 388 9514 420
rect 9546 388 9582 420
rect 9614 388 9650 420
rect 9682 388 9718 420
rect 9750 388 9786 420
rect 9818 388 9854 420
rect 9886 388 9922 420
rect 9954 388 9990 420
rect 10022 388 10058 420
rect 10090 388 10126 420
rect 10158 388 10194 420
rect 10226 388 10262 420
rect 10294 388 10330 420
rect 10362 388 10398 420
rect 10430 388 10466 420
rect 10498 388 10534 420
rect 10566 388 10602 420
rect 10634 388 10670 420
rect 10702 388 10738 420
rect 10770 388 10806 420
rect 10838 388 10874 420
rect 10906 388 10942 420
rect 10974 388 11010 420
rect 11042 388 11078 420
rect 11110 388 11146 420
rect 11178 388 11214 420
rect 11246 388 11282 420
rect 11314 388 11350 420
rect 11382 388 11418 420
rect 11450 388 11486 420
rect 11518 388 11554 420
rect 11586 388 11622 420
rect 11654 388 11690 420
rect 11722 388 11758 420
rect 11790 388 11826 420
rect 11858 388 11894 420
rect 11926 388 11962 420
rect 11994 388 12030 420
rect 12062 388 12098 420
rect 12130 388 12166 420
rect 12198 388 12234 420
rect 12266 388 12302 420
rect 12334 388 12370 420
rect 12402 388 12438 420
rect 12470 388 12506 420
rect 12538 388 12574 420
rect 12606 388 12642 420
rect 12674 388 12710 420
rect 12742 388 12778 420
rect 12810 388 12846 420
rect 12878 388 12914 420
rect 12946 388 12982 420
rect 13014 388 13050 420
rect 13082 388 13118 420
rect 13150 388 13186 420
rect 13218 388 13254 420
rect 13286 388 13322 420
rect 13354 388 13390 420
rect 13422 388 13458 420
rect 13490 388 13526 420
rect 13558 388 13594 420
rect 13626 388 13662 420
rect 13694 388 13730 420
rect 13762 388 13798 420
rect 13830 388 13866 420
rect 13898 388 13934 420
rect 13966 388 14002 420
rect 14034 388 14070 420
rect 14102 388 14138 420
rect 14170 388 14206 420
rect 14238 388 14274 420
rect 14306 388 14342 420
rect 14374 388 14410 420
rect 14442 388 14478 420
rect 14510 388 14546 420
rect 14578 388 14614 420
rect 14646 388 14682 420
rect 14714 388 14750 420
rect 14782 388 14818 420
rect 14850 388 14886 420
rect 14918 388 14954 420
rect 14986 388 15022 420
rect 15054 388 15090 420
rect 15122 388 15158 420
rect 15190 388 15226 420
rect 15258 388 15294 420
rect 15326 388 15362 420
rect 15394 388 15430 420
rect 15462 388 15498 420
rect 15530 388 15566 420
rect 15598 388 15640 420
rect 360 370 15640 388
<< nsubdiff >>
rect 0 1962 16000 1980
rect 0 1930 28 1962
rect 60 1930 96 1962
rect 128 1930 164 1962
rect 196 1930 232 1962
rect 264 1930 300 1962
rect 332 1930 368 1962
rect 400 1930 436 1962
rect 468 1930 504 1962
rect 536 1930 572 1962
rect 604 1930 640 1962
rect 672 1930 708 1962
rect 740 1930 776 1962
rect 808 1930 844 1962
rect 876 1930 912 1962
rect 944 1930 980 1962
rect 1012 1930 1048 1962
rect 1080 1930 1116 1962
rect 1148 1930 1184 1962
rect 1216 1930 1252 1962
rect 1284 1930 1320 1962
rect 1352 1930 1388 1962
rect 1420 1930 1456 1962
rect 1488 1930 1524 1962
rect 1556 1930 1592 1962
rect 1624 1930 1660 1962
rect 1692 1930 1728 1962
rect 1760 1930 1796 1962
rect 1828 1930 1864 1962
rect 1896 1930 1932 1962
rect 1964 1930 2000 1962
rect 2032 1930 2068 1962
rect 2100 1930 2136 1962
rect 2168 1930 2204 1962
rect 2236 1930 2272 1962
rect 2304 1930 2340 1962
rect 2372 1930 2408 1962
rect 2440 1930 2476 1962
rect 2508 1930 2544 1962
rect 2576 1930 2612 1962
rect 2644 1930 2680 1962
rect 2712 1930 2748 1962
rect 2780 1930 2816 1962
rect 2848 1930 2884 1962
rect 2916 1930 2952 1962
rect 2984 1930 3020 1962
rect 3052 1930 3088 1962
rect 3120 1930 3156 1962
rect 3188 1930 3224 1962
rect 3256 1930 3292 1962
rect 3324 1930 3360 1962
rect 3392 1930 3428 1962
rect 3460 1930 3496 1962
rect 3528 1930 3564 1962
rect 3596 1930 3632 1962
rect 3664 1930 3700 1962
rect 3732 1930 3768 1962
rect 3800 1930 3836 1962
rect 3868 1930 3904 1962
rect 3936 1930 3972 1962
rect 4004 1930 4040 1962
rect 4072 1930 4108 1962
rect 4140 1930 4176 1962
rect 4208 1930 4244 1962
rect 4276 1930 4312 1962
rect 4344 1930 4380 1962
rect 4412 1930 4448 1962
rect 4480 1930 4516 1962
rect 4548 1930 4584 1962
rect 4616 1930 4652 1962
rect 4684 1930 4720 1962
rect 4752 1930 4788 1962
rect 4820 1930 4856 1962
rect 4888 1930 4924 1962
rect 4956 1930 4992 1962
rect 5024 1930 5060 1962
rect 5092 1930 5128 1962
rect 5160 1930 5196 1962
rect 5228 1930 5264 1962
rect 5296 1930 5332 1962
rect 5364 1930 5400 1962
rect 5432 1930 5468 1962
rect 5500 1930 5536 1962
rect 5568 1930 5604 1962
rect 5636 1930 5672 1962
rect 5704 1930 5740 1962
rect 5772 1930 5808 1962
rect 5840 1930 5876 1962
rect 5908 1930 5944 1962
rect 5976 1930 6012 1962
rect 6044 1930 6080 1962
rect 6112 1930 6148 1962
rect 6180 1930 6216 1962
rect 6248 1930 6284 1962
rect 6316 1930 6352 1962
rect 6384 1930 6420 1962
rect 6452 1930 6488 1962
rect 6520 1930 6556 1962
rect 6588 1930 6624 1962
rect 6656 1930 6692 1962
rect 6724 1930 6760 1962
rect 6792 1930 6828 1962
rect 6860 1930 6896 1962
rect 6928 1930 6964 1962
rect 6996 1930 7032 1962
rect 7064 1930 7100 1962
rect 7132 1930 7168 1962
rect 7200 1930 7236 1962
rect 7268 1930 7304 1962
rect 7336 1930 7372 1962
rect 7404 1930 7440 1962
rect 7472 1930 7508 1962
rect 7540 1930 7576 1962
rect 7608 1930 7644 1962
rect 7676 1930 7712 1962
rect 7744 1930 7780 1962
rect 7812 1930 7848 1962
rect 7880 1930 7916 1962
rect 7948 1930 7984 1962
rect 8016 1930 8052 1962
rect 8084 1930 8120 1962
rect 8152 1930 8188 1962
rect 8220 1930 8256 1962
rect 8288 1930 8324 1962
rect 8356 1930 8392 1962
rect 8424 1930 8460 1962
rect 8492 1930 8528 1962
rect 8560 1930 8596 1962
rect 8628 1930 8664 1962
rect 8696 1930 8732 1962
rect 8764 1930 8800 1962
rect 8832 1930 8868 1962
rect 8900 1930 8936 1962
rect 8968 1930 9004 1962
rect 9036 1930 9072 1962
rect 9104 1930 9140 1962
rect 9172 1930 9208 1962
rect 9240 1930 9276 1962
rect 9308 1930 9344 1962
rect 9376 1930 9412 1962
rect 9444 1930 9480 1962
rect 9512 1930 9548 1962
rect 9580 1930 9616 1962
rect 9648 1930 9684 1962
rect 9716 1930 9752 1962
rect 9784 1930 9820 1962
rect 9852 1930 9888 1962
rect 9920 1930 9956 1962
rect 9988 1930 10024 1962
rect 10056 1930 10092 1962
rect 10124 1930 10160 1962
rect 10192 1930 10228 1962
rect 10260 1930 10296 1962
rect 10328 1930 10364 1962
rect 10396 1930 10432 1962
rect 10464 1930 10500 1962
rect 10532 1930 10568 1962
rect 10600 1930 10636 1962
rect 10668 1930 10704 1962
rect 10736 1930 10772 1962
rect 10804 1930 10840 1962
rect 10872 1930 10908 1962
rect 10940 1930 10976 1962
rect 11008 1930 11044 1962
rect 11076 1930 11112 1962
rect 11144 1930 11180 1962
rect 11212 1930 11248 1962
rect 11280 1930 11316 1962
rect 11348 1930 11384 1962
rect 11416 1930 11452 1962
rect 11484 1930 11520 1962
rect 11552 1930 11588 1962
rect 11620 1930 11656 1962
rect 11688 1930 11724 1962
rect 11756 1930 11792 1962
rect 11824 1930 11860 1962
rect 11892 1930 11928 1962
rect 11960 1930 11996 1962
rect 12028 1930 12064 1962
rect 12096 1930 12132 1962
rect 12164 1930 12200 1962
rect 12232 1930 12268 1962
rect 12300 1930 12336 1962
rect 12368 1930 12404 1962
rect 12436 1930 12472 1962
rect 12504 1930 12540 1962
rect 12572 1930 12608 1962
rect 12640 1930 12676 1962
rect 12708 1930 12744 1962
rect 12776 1930 12812 1962
rect 12844 1930 12880 1962
rect 12912 1930 12948 1962
rect 12980 1930 13016 1962
rect 13048 1930 13084 1962
rect 13116 1930 13152 1962
rect 13184 1930 13220 1962
rect 13252 1930 13288 1962
rect 13320 1930 13356 1962
rect 13388 1930 13424 1962
rect 13456 1930 13492 1962
rect 13524 1930 13560 1962
rect 13592 1930 13628 1962
rect 13660 1930 13696 1962
rect 13728 1930 13764 1962
rect 13796 1930 13832 1962
rect 13864 1930 13900 1962
rect 13932 1930 13968 1962
rect 14000 1930 14036 1962
rect 14068 1930 14104 1962
rect 14136 1930 14172 1962
rect 14204 1930 14240 1962
rect 14272 1930 14308 1962
rect 14340 1930 14376 1962
rect 14408 1930 14444 1962
rect 14476 1930 14512 1962
rect 14544 1930 14580 1962
rect 14612 1930 14648 1962
rect 14680 1930 14716 1962
rect 14748 1930 14784 1962
rect 14816 1930 14852 1962
rect 14884 1930 14920 1962
rect 14952 1930 14988 1962
rect 15020 1930 15056 1962
rect 15088 1930 15124 1962
rect 15156 1930 15192 1962
rect 15224 1930 15260 1962
rect 15292 1930 15328 1962
rect 15360 1930 15396 1962
rect 15428 1930 15464 1962
rect 15496 1930 15532 1962
rect 15564 1930 15600 1962
rect 15632 1930 15668 1962
rect 15700 1930 15736 1962
rect 15768 1930 15804 1962
rect 15836 1930 15872 1962
rect 15904 1930 15940 1962
rect 15972 1930 16000 1962
rect 0 1912 16000 1930
rect 0 1856 68 1912
rect 0 1824 18 1856
rect 50 1824 68 1856
rect 0 1788 68 1824
rect 0 1756 18 1788
rect 50 1756 68 1788
rect 0 1720 68 1756
rect 0 1688 18 1720
rect 50 1688 68 1720
rect 0 1652 68 1688
rect 0 1620 18 1652
rect 50 1620 68 1652
rect 15932 1856 16000 1912
rect 15932 1824 15950 1856
rect 15982 1824 16000 1856
rect 15932 1788 16000 1824
rect 15932 1756 15950 1788
rect 15982 1756 16000 1788
rect 15932 1720 16000 1756
rect 15932 1688 15950 1720
rect 15982 1688 16000 1720
rect 15932 1652 16000 1688
rect 0 1584 68 1620
rect 0 1552 18 1584
rect 50 1552 68 1584
rect 0 1516 68 1552
rect 0 1484 18 1516
rect 50 1484 68 1516
rect 0 1448 68 1484
rect 0 1416 18 1448
rect 50 1416 68 1448
rect 0 1380 68 1416
rect 0 1348 18 1380
rect 50 1348 68 1380
rect 0 1312 68 1348
rect 0 1280 18 1312
rect 50 1280 68 1312
rect 0 1244 68 1280
rect 0 1212 18 1244
rect 50 1212 68 1244
rect 0 1176 68 1212
rect 0 1144 18 1176
rect 50 1144 68 1176
rect 0 1108 68 1144
rect 0 1076 18 1108
rect 50 1076 68 1108
rect 0 1040 68 1076
rect 0 1008 18 1040
rect 50 1008 68 1040
rect 0 972 68 1008
rect 0 940 18 972
rect 50 940 68 972
rect 0 904 68 940
rect 0 872 18 904
rect 50 872 68 904
rect 0 836 68 872
rect 0 804 18 836
rect 50 804 68 836
rect 0 768 68 804
rect 0 736 18 768
rect 50 736 68 768
rect 0 700 68 736
rect 0 668 18 700
rect 50 668 68 700
rect 0 632 68 668
rect 0 600 18 632
rect 50 600 68 632
rect 0 564 68 600
rect 0 532 18 564
rect 50 532 68 564
rect 0 496 68 532
rect 0 464 18 496
rect 50 464 68 496
rect 0 428 68 464
rect 0 396 18 428
rect 50 396 68 428
rect 0 360 68 396
rect 15932 1620 15950 1652
rect 15982 1620 16000 1652
rect 15932 1584 16000 1620
rect 15932 1552 15950 1584
rect 15982 1552 16000 1584
rect 15932 1516 16000 1552
rect 15932 1484 15950 1516
rect 15982 1484 16000 1516
rect 15932 1448 16000 1484
rect 15932 1416 15950 1448
rect 15982 1416 16000 1448
rect 15932 1380 16000 1416
rect 15932 1348 15950 1380
rect 15982 1348 16000 1380
rect 15932 1312 16000 1348
rect 15932 1280 15950 1312
rect 15982 1280 16000 1312
rect 15932 1244 16000 1280
rect 15932 1212 15950 1244
rect 15982 1212 16000 1244
rect 15932 1176 16000 1212
rect 15932 1144 15950 1176
rect 15982 1144 16000 1176
rect 15932 1108 16000 1144
rect 15932 1076 15950 1108
rect 15982 1076 16000 1108
rect 15932 1040 16000 1076
rect 15932 1008 15950 1040
rect 15982 1008 16000 1040
rect 15932 972 16000 1008
rect 15932 940 15950 972
rect 15982 940 16000 972
rect 15932 904 16000 940
rect 15932 872 15950 904
rect 15982 872 16000 904
rect 15932 836 16000 872
rect 15932 804 15950 836
rect 15982 804 16000 836
rect 15932 768 16000 804
rect 15932 736 15950 768
rect 15982 736 16000 768
rect 15932 700 16000 736
rect 15932 668 15950 700
rect 15982 668 16000 700
rect 15932 632 16000 668
rect 15932 600 15950 632
rect 15982 600 16000 632
rect 15932 564 16000 600
rect 15932 532 15950 564
rect 15982 532 16000 564
rect 15932 496 16000 532
rect 15932 464 15950 496
rect 15982 464 16000 496
rect 15932 428 16000 464
rect 15932 396 15950 428
rect 15982 396 16000 428
rect 0 328 18 360
rect 50 328 68 360
rect 0 292 68 328
rect 0 260 18 292
rect 50 260 68 292
rect 0 224 68 260
rect 0 192 18 224
rect 50 192 68 224
rect 0 156 68 192
rect 0 124 18 156
rect 50 124 68 156
rect 0 68 68 124
rect 15932 360 16000 396
rect 15932 328 15950 360
rect 15982 328 16000 360
rect 15932 292 16000 328
rect 15932 260 15950 292
rect 15982 260 16000 292
rect 15932 224 16000 260
rect 15932 192 15950 224
rect 15982 192 16000 224
rect 15932 156 16000 192
rect 15932 124 15950 156
rect 15982 124 16000 156
rect 15932 68 16000 124
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 2 16000 18
rect 2 0 16000 2
<< psubdiffcont >>
rect 402 1580 434 1612
rect 470 1580 502 1612
rect 538 1580 570 1612
rect 606 1580 638 1612
rect 674 1580 706 1612
rect 742 1580 774 1612
rect 810 1580 842 1612
rect 878 1580 910 1612
rect 946 1580 978 1612
rect 1014 1580 1046 1612
rect 1082 1580 1114 1612
rect 1150 1580 1182 1612
rect 1218 1580 1250 1612
rect 1286 1580 1318 1612
rect 1354 1580 1386 1612
rect 1422 1580 1454 1612
rect 1490 1580 1522 1612
rect 1558 1580 1590 1612
rect 1626 1580 1658 1612
rect 1694 1580 1726 1612
rect 1762 1580 1794 1612
rect 1830 1580 1862 1612
rect 1898 1580 1930 1612
rect 1966 1580 1998 1612
rect 2034 1580 2066 1612
rect 2102 1580 2134 1612
rect 2170 1580 2202 1612
rect 2238 1580 2270 1612
rect 2306 1580 2338 1612
rect 2374 1580 2406 1612
rect 2442 1580 2474 1612
rect 2510 1580 2542 1612
rect 2578 1580 2610 1612
rect 2646 1580 2678 1612
rect 2714 1580 2746 1612
rect 2782 1580 2814 1612
rect 2850 1580 2882 1612
rect 2918 1580 2950 1612
rect 2986 1580 3018 1612
rect 3054 1580 3086 1612
rect 3122 1580 3154 1612
rect 3190 1580 3222 1612
rect 3258 1580 3290 1612
rect 3326 1580 3358 1612
rect 3394 1580 3426 1612
rect 3462 1580 3494 1612
rect 3530 1580 3562 1612
rect 3598 1580 3630 1612
rect 3666 1580 3698 1612
rect 3734 1580 3766 1612
rect 3802 1580 3834 1612
rect 3870 1580 3902 1612
rect 3938 1580 3970 1612
rect 4006 1580 4038 1612
rect 4074 1580 4106 1612
rect 4142 1580 4174 1612
rect 4210 1580 4242 1612
rect 4278 1580 4310 1612
rect 4346 1580 4378 1612
rect 4414 1580 4446 1612
rect 4482 1580 4514 1612
rect 4550 1580 4582 1612
rect 4618 1580 4650 1612
rect 4686 1580 4718 1612
rect 4754 1580 4786 1612
rect 4822 1580 4854 1612
rect 4890 1580 4922 1612
rect 4958 1580 4990 1612
rect 5026 1580 5058 1612
rect 5094 1580 5126 1612
rect 5162 1580 5194 1612
rect 5230 1580 5262 1612
rect 5298 1580 5330 1612
rect 5366 1580 5398 1612
rect 5434 1580 5466 1612
rect 5502 1580 5534 1612
rect 5570 1580 5602 1612
rect 5638 1580 5670 1612
rect 5706 1580 5738 1612
rect 5774 1580 5806 1612
rect 5842 1580 5874 1612
rect 5910 1580 5942 1612
rect 5978 1580 6010 1612
rect 6046 1580 6078 1612
rect 6114 1580 6146 1612
rect 6182 1580 6214 1612
rect 6250 1580 6282 1612
rect 6318 1580 6350 1612
rect 6386 1580 6418 1612
rect 6454 1580 6486 1612
rect 6522 1580 6554 1612
rect 6590 1580 6622 1612
rect 6658 1580 6690 1612
rect 6726 1580 6758 1612
rect 6794 1580 6826 1612
rect 6862 1580 6894 1612
rect 6930 1580 6962 1612
rect 6998 1580 7030 1612
rect 7066 1580 7098 1612
rect 7134 1580 7166 1612
rect 7202 1580 7234 1612
rect 7270 1580 7302 1612
rect 7338 1580 7370 1612
rect 7406 1580 7438 1612
rect 7474 1580 7506 1612
rect 7542 1580 7574 1612
rect 7610 1580 7642 1612
rect 7678 1580 7710 1612
rect 7746 1580 7778 1612
rect 7814 1580 7846 1612
rect 7882 1580 7914 1612
rect 7950 1580 7982 1612
rect 8018 1580 8050 1612
rect 8086 1580 8118 1612
rect 8154 1580 8186 1612
rect 8222 1580 8254 1612
rect 8290 1580 8322 1612
rect 8358 1580 8390 1612
rect 8426 1580 8458 1612
rect 8494 1580 8526 1612
rect 8562 1580 8594 1612
rect 8630 1580 8662 1612
rect 8698 1580 8730 1612
rect 8766 1580 8798 1612
rect 8834 1580 8866 1612
rect 8902 1580 8934 1612
rect 8970 1580 9002 1612
rect 9038 1580 9070 1612
rect 9106 1580 9138 1612
rect 9174 1580 9206 1612
rect 9242 1580 9274 1612
rect 9310 1580 9342 1612
rect 9378 1580 9410 1612
rect 9446 1580 9478 1612
rect 9514 1580 9546 1612
rect 9582 1580 9614 1612
rect 9650 1580 9682 1612
rect 9718 1580 9750 1612
rect 9786 1580 9818 1612
rect 9854 1580 9886 1612
rect 9922 1580 9954 1612
rect 9990 1580 10022 1612
rect 10058 1580 10090 1612
rect 10126 1580 10158 1612
rect 10194 1580 10226 1612
rect 10262 1580 10294 1612
rect 10330 1580 10362 1612
rect 10398 1580 10430 1612
rect 10466 1580 10498 1612
rect 10534 1580 10566 1612
rect 10602 1580 10634 1612
rect 10670 1580 10702 1612
rect 10738 1580 10770 1612
rect 10806 1580 10838 1612
rect 10874 1580 10906 1612
rect 10942 1580 10974 1612
rect 11010 1580 11042 1612
rect 11078 1580 11110 1612
rect 11146 1580 11178 1612
rect 11214 1580 11246 1612
rect 11282 1580 11314 1612
rect 11350 1580 11382 1612
rect 11418 1580 11450 1612
rect 11486 1580 11518 1612
rect 11554 1580 11586 1612
rect 11622 1580 11654 1612
rect 11690 1580 11722 1612
rect 11758 1580 11790 1612
rect 11826 1580 11858 1612
rect 11894 1580 11926 1612
rect 11962 1580 11994 1612
rect 12030 1580 12062 1612
rect 12098 1580 12130 1612
rect 12166 1580 12198 1612
rect 12234 1580 12266 1612
rect 12302 1580 12334 1612
rect 12370 1580 12402 1612
rect 12438 1580 12470 1612
rect 12506 1580 12538 1612
rect 12574 1580 12606 1612
rect 12642 1580 12674 1612
rect 12710 1580 12742 1612
rect 12778 1580 12810 1612
rect 12846 1580 12878 1612
rect 12914 1580 12946 1612
rect 12982 1580 13014 1612
rect 13050 1580 13082 1612
rect 13118 1580 13150 1612
rect 13186 1580 13218 1612
rect 13254 1580 13286 1612
rect 13322 1580 13354 1612
rect 13390 1580 13422 1612
rect 13458 1580 13490 1612
rect 13526 1580 13558 1612
rect 13594 1580 13626 1612
rect 13662 1580 13694 1612
rect 13730 1580 13762 1612
rect 13798 1580 13830 1612
rect 13866 1580 13898 1612
rect 13934 1580 13966 1612
rect 14002 1580 14034 1612
rect 14070 1580 14102 1612
rect 14138 1580 14170 1612
rect 14206 1580 14238 1612
rect 14274 1580 14306 1612
rect 14342 1580 14374 1612
rect 14410 1580 14442 1612
rect 14478 1580 14510 1612
rect 14546 1580 14578 1612
rect 14614 1580 14646 1612
rect 14682 1580 14714 1612
rect 14750 1580 14782 1612
rect 14818 1580 14850 1612
rect 14886 1580 14918 1612
rect 14954 1580 14986 1612
rect 15022 1580 15054 1612
rect 15090 1580 15122 1612
rect 15158 1580 15190 1612
rect 15226 1580 15258 1612
rect 15294 1580 15326 1612
rect 15362 1580 15394 1612
rect 15430 1580 15462 1612
rect 15498 1580 15530 1612
rect 15566 1580 15598 1612
rect 378 1494 410 1526
rect 378 1426 410 1458
rect 15590 1494 15622 1526
rect 378 1358 410 1390
rect 378 1290 410 1322
rect 378 1222 410 1254
rect 378 1154 410 1186
rect 378 1086 410 1118
rect 378 1018 410 1050
rect 378 950 410 982
rect 378 882 410 914
rect 378 814 410 846
rect 378 746 410 778
rect 378 678 410 710
rect 378 610 410 642
rect 378 542 410 574
rect 15590 1426 15622 1458
rect 15590 1358 15622 1390
rect 15590 1290 15622 1322
rect 15590 1222 15622 1254
rect 15590 1154 15622 1186
rect 15590 1086 15622 1118
rect 15590 1018 15622 1050
rect 15590 950 15622 982
rect 15590 882 15622 914
rect 15590 814 15622 846
rect 15590 746 15622 778
rect 15590 678 15622 710
rect 15590 610 15622 642
rect 378 474 410 506
rect 15590 542 15622 574
rect 15590 474 15622 506
rect 402 388 434 420
rect 470 388 502 420
rect 538 388 570 420
rect 606 388 638 420
rect 674 388 706 420
rect 742 388 774 420
rect 810 388 842 420
rect 878 388 910 420
rect 946 388 978 420
rect 1014 388 1046 420
rect 1082 388 1114 420
rect 1150 388 1182 420
rect 1218 388 1250 420
rect 1286 388 1318 420
rect 1354 388 1386 420
rect 1422 388 1454 420
rect 1490 388 1522 420
rect 1558 388 1590 420
rect 1626 388 1658 420
rect 1694 388 1726 420
rect 1762 388 1794 420
rect 1830 388 1862 420
rect 1898 388 1930 420
rect 1966 388 1998 420
rect 2034 388 2066 420
rect 2102 388 2134 420
rect 2170 388 2202 420
rect 2238 388 2270 420
rect 2306 388 2338 420
rect 2374 388 2406 420
rect 2442 388 2474 420
rect 2510 388 2542 420
rect 2578 388 2610 420
rect 2646 388 2678 420
rect 2714 388 2746 420
rect 2782 388 2814 420
rect 2850 388 2882 420
rect 2918 388 2950 420
rect 2986 388 3018 420
rect 3054 388 3086 420
rect 3122 388 3154 420
rect 3190 388 3222 420
rect 3258 388 3290 420
rect 3326 388 3358 420
rect 3394 388 3426 420
rect 3462 388 3494 420
rect 3530 388 3562 420
rect 3598 388 3630 420
rect 3666 388 3698 420
rect 3734 388 3766 420
rect 3802 388 3834 420
rect 3870 388 3902 420
rect 3938 388 3970 420
rect 4006 388 4038 420
rect 4074 388 4106 420
rect 4142 388 4174 420
rect 4210 388 4242 420
rect 4278 388 4310 420
rect 4346 388 4378 420
rect 4414 388 4446 420
rect 4482 388 4514 420
rect 4550 388 4582 420
rect 4618 388 4650 420
rect 4686 388 4718 420
rect 4754 388 4786 420
rect 4822 388 4854 420
rect 4890 388 4922 420
rect 4958 388 4990 420
rect 5026 388 5058 420
rect 5094 388 5126 420
rect 5162 388 5194 420
rect 5230 388 5262 420
rect 5298 388 5330 420
rect 5366 388 5398 420
rect 5434 388 5466 420
rect 5502 388 5534 420
rect 5570 388 5602 420
rect 5638 388 5670 420
rect 5706 388 5738 420
rect 5774 388 5806 420
rect 5842 388 5874 420
rect 5910 388 5942 420
rect 5978 388 6010 420
rect 6046 388 6078 420
rect 6114 388 6146 420
rect 6182 388 6214 420
rect 6250 388 6282 420
rect 6318 388 6350 420
rect 6386 388 6418 420
rect 6454 388 6486 420
rect 6522 388 6554 420
rect 6590 388 6622 420
rect 6658 388 6690 420
rect 6726 388 6758 420
rect 6794 388 6826 420
rect 6862 388 6894 420
rect 6930 388 6962 420
rect 6998 388 7030 420
rect 7066 388 7098 420
rect 7134 388 7166 420
rect 7202 388 7234 420
rect 7270 388 7302 420
rect 7338 388 7370 420
rect 7406 388 7438 420
rect 7474 388 7506 420
rect 7542 388 7574 420
rect 7610 388 7642 420
rect 7678 388 7710 420
rect 7746 388 7778 420
rect 7814 388 7846 420
rect 7882 388 7914 420
rect 7950 388 7982 420
rect 8018 388 8050 420
rect 8086 388 8118 420
rect 8154 388 8186 420
rect 8222 388 8254 420
rect 8290 388 8322 420
rect 8358 388 8390 420
rect 8426 388 8458 420
rect 8494 388 8526 420
rect 8562 388 8594 420
rect 8630 388 8662 420
rect 8698 388 8730 420
rect 8766 388 8798 420
rect 8834 388 8866 420
rect 8902 388 8934 420
rect 8970 388 9002 420
rect 9038 388 9070 420
rect 9106 388 9138 420
rect 9174 388 9206 420
rect 9242 388 9274 420
rect 9310 388 9342 420
rect 9378 388 9410 420
rect 9446 388 9478 420
rect 9514 388 9546 420
rect 9582 388 9614 420
rect 9650 388 9682 420
rect 9718 388 9750 420
rect 9786 388 9818 420
rect 9854 388 9886 420
rect 9922 388 9954 420
rect 9990 388 10022 420
rect 10058 388 10090 420
rect 10126 388 10158 420
rect 10194 388 10226 420
rect 10262 388 10294 420
rect 10330 388 10362 420
rect 10398 388 10430 420
rect 10466 388 10498 420
rect 10534 388 10566 420
rect 10602 388 10634 420
rect 10670 388 10702 420
rect 10738 388 10770 420
rect 10806 388 10838 420
rect 10874 388 10906 420
rect 10942 388 10974 420
rect 11010 388 11042 420
rect 11078 388 11110 420
rect 11146 388 11178 420
rect 11214 388 11246 420
rect 11282 388 11314 420
rect 11350 388 11382 420
rect 11418 388 11450 420
rect 11486 388 11518 420
rect 11554 388 11586 420
rect 11622 388 11654 420
rect 11690 388 11722 420
rect 11758 388 11790 420
rect 11826 388 11858 420
rect 11894 388 11926 420
rect 11962 388 11994 420
rect 12030 388 12062 420
rect 12098 388 12130 420
rect 12166 388 12198 420
rect 12234 388 12266 420
rect 12302 388 12334 420
rect 12370 388 12402 420
rect 12438 388 12470 420
rect 12506 388 12538 420
rect 12574 388 12606 420
rect 12642 388 12674 420
rect 12710 388 12742 420
rect 12778 388 12810 420
rect 12846 388 12878 420
rect 12914 388 12946 420
rect 12982 388 13014 420
rect 13050 388 13082 420
rect 13118 388 13150 420
rect 13186 388 13218 420
rect 13254 388 13286 420
rect 13322 388 13354 420
rect 13390 388 13422 420
rect 13458 388 13490 420
rect 13526 388 13558 420
rect 13594 388 13626 420
rect 13662 388 13694 420
rect 13730 388 13762 420
rect 13798 388 13830 420
rect 13866 388 13898 420
rect 13934 388 13966 420
rect 14002 388 14034 420
rect 14070 388 14102 420
rect 14138 388 14170 420
rect 14206 388 14238 420
rect 14274 388 14306 420
rect 14342 388 14374 420
rect 14410 388 14442 420
rect 14478 388 14510 420
rect 14546 388 14578 420
rect 14614 388 14646 420
rect 14682 388 14714 420
rect 14750 388 14782 420
rect 14818 388 14850 420
rect 14886 388 14918 420
rect 14954 388 14986 420
rect 15022 388 15054 420
rect 15090 388 15122 420
rect 15158 388 15190 420
rect 15226 388 15258 420
rect 15294 388 15326 420
rect 15362 388 15394 420
rect 15430 388 15462 420
rect 15498 388 15530 420
rect 15566 388 15598 420
<< nsubdiffcont >>
rect 28 1930 60 1962
rect 96 1930 128 1962
rect 164 1930 196 1962
rect 232 1930 264 1962
rect 300 1930 332 1962
rect 368 1930 400 1962
rect 436 1930 468 1962
rect 504 1930 536 1962
rect 572 1930 604 1962
rect 640 1930 672 1962
rect 708 1930 740 1962
rect 776 1930 808 1962
rect 844 1930 876 1962
rect 912 1930 944 1962
rect 980 1930 1012 1962
rect 1048 1930 1080 1962
rect 1116 1930 1148 1962
rect 1184 1930 1216 1962
rect 1252 1930 1284 1962
rect 1320 1930 1352 1962
rect 1388 1930 1420 1962
rect 1456 1930 1488 1962
rect 1524 1930 1556 1962
rect 1592 1930 1624 1962
rect 1660 1930 1692 1962
rect 1728 1930 1760 1962
rect 1796 1930 1828 1962
rect 1864 1930 1896 1962
rect 1932 1930 1964 1962
rect 2000 1930 2032 1962
rect 2068 1930 2100 1962
rect 2136 1930 2168 1962
rect 2204 1930 2236 1962
rect 2272 1930 2304 1962
rect 2340 1930 2372 1962
rect 2408 1930 2440 1962
rect 2476 1930 2508 1962
rect 2544 1930 2576 1962
rect 2612 1930 2644 1962
rect 2680 1930 2712 1962
rect 2748 1930 2780 1962
rect 2816 1930 2848 1962
rect 2884 1930 2916 1962
rect 2952 1930 2984 1962
rect 3020 1930 3052 1962
rect 3088 1930 3120 1962
rect 3156 1930 3188 1962
rect 3224 1930 3256 1962
rect 3292 1930 3324 1962
rect 3360 1930 3392 1962
rect 3428 1930 3460 1962
rect 3496 1930 3528 1962
rect 3564 1930 3596 1962
rect 3632 1930 3664 1962
rect 3700 1930 3732 1962
rect 3768 1930 3800 1962
rect 3836 1930 3868 1962
rect 3904 1930 3936 1962
rect 3972 1930 4004 1962
rect 4040 1930 4072 1962
rect 4108 1930 4140 1962
rect 4176 1930 4208 1962
rect 4244 1930 4276 1962
rect 4312 1930 4344 1962
rect 4380 1930 4412 1962
rect 4448 1930 4480 1962
rect 4516 1930 4548 1962
rect 4584 1930 4616 1962
rect 4652 1930 4684 1962
rect 4720 1930 4752 1962
rect 4788 1930 4820 1962
rect 4856 1930 4888 1962
rect 4924 1930 4956 1962
rect 4992 1930 5024 1962
rect 5060 1930 5092 1962
rect 5128 1930 5160 1962
rect 5196 1930 5228 1962
rect 5264 1930 5296 1962
rect 5332 1930 5364 1962
rect 5400 1930 5432 1962
rect 5468 1930 5500 1962
rect 5536 1930 5568 1962
rect 5604 1930 5636 1962
rect 5672 1930 5704 1962
rect 5740 1930 5772 1962
rect 5808 1930 5840 1962
rect 5876 1930 5908 1962
rect 5944 1930 5976 1962
rect 6012 1930 6044 1962
rect 6080 1930 6112 1962
rect 6148 1930 6180 1962
rect 6216 1930 6248 1962
rect 6284 1930 6316 1962
rect 6352 1930 6384 1962
rect 6420 1930 6452 1962
rect 6488 1930 6520 1962
rect 6556 1930 6588 1962
rect 6624 1930 6656 1962
rect 6692 1930 6724 1962
rect 6760 1930 6792 1962
rect 6828 1930 6860 1962
rect 6896 1930 6928 1962
rect 6964 1930 6996 1962
rect 7032 1930 7064 1962
rect 7100 1930 7132 1962
rect 7168 1930 7200 1962
rect 7236 1930 7268 1962
rect 7304 1930 7336 1962
rect 7372 1930 7404 1962
rect 7440 1930 7472 1962
rect 7508 1930 7540 1962
rect 7576 1930 7608 1962
rect 7644 1930 7676 1962
rect 7712 1930 7744 1962
rect 7780 1930 7812 1962
rect 7848 1930 7880 1962
rect 7916 1930 7948 1962
rect 7984 1930 8016 1962
rect 8052 1930 8084 1962
rect 8120 1930 8152 1962
rect 8188 1930 8220 1962
rect 8256 1930 8288 1962
rect 8324 1930 8356 1962
rect 8392 1930 8424 1962
rect 8460 1930 8492 1962
rect 8528 1930 8560 1962
rect 8596 1930 8628 1962
rect 8664 1930 8696 1962
rect 8732 1930 8764 1962
rect 8800 1930 8832 1962
rect 8868 1930 8900 1962
rect 8936 1930 8968 1962
rect 9004 1930 9036 1962
rect 9072 1930 9104 1962
rect 9140 1930 9172 1962
rect 9208 1930 9240 1962
rect 9276 1930 9308 1962
rect 9344 1930 9376 1962
rect 9412 1930 9444 1962
rect 9480 1930 9512 1962
rect 9548 1930 9580 1962
rect 9616 1930 9648 1962
rect 9684 1930 9716 1962
rect 9752 1930 9784 1962
rect 9820 1930 9852 1962
rect 9888 1930 9920 1962
rect 9956 1930 9988 1962
rect 10024 1930 10056 1962
rect 10092 1930 10124 1962
rect 10160 1930 10192 1962
rect 10228 1930 10260 1962
rect 10296 1930 10328 1962
rect 10364 1930 10396 1962
rect 10432 1930 10464 1962
rect 10500 1930 10532 1962
rect 10568 1930 10600 1962
rect 10636 1930 10668 1962
rect 10704 1930 10736 1962
rect 10772 1930 10804 1962
rect 10840 1930 10872 1962
rect 10908 1930 10940 1962
rect 10976 1930 11008 1962
rect 11044 1930 11076 1962
rect 11112 1930 11144 1962
rect 11180 1930 11212 1962
rect 11248 1930 11280 1962
rect 11316 1930 11348 1962
rect 11384 1930 11416 1962
rect 11452 1930 11484 1962
rect 11520 1930 11552 1962
rect 11588 1930 11620 1962
rect 11656 1930 11688 1962
rect 11724 1930 11756 1962
rect 11792 1930 11824 1962
rect 11860 1930 11892 1962
rect 11928 1930 11960 1962
rect 11996 1930 12028 1962
rect 12064 1930 12096 1962
rect 12132 1930 12164 1962
rect 12200 1930 12232 1962
rect 12268 1930 12300 1962
rect 12336 1930 12368 1962
rect 12404 1930 12436 1962
rect 12472 1930 12504 1962
rect 12540 1930 12572 1962
rect 12608 1930 12640 1962
rect 12676 1930 12708 1962
rect 12744 1930 12776 1962
rect 12812 1930 12844 1962
rect 12880 1930 12912 1962
rect 12948 1930 12980 1962
rect 13016 1930 13048 1962
rect 13084 1930 13116 1962
rect 13152 1930 13184 1962
rect 13220 1930 13252 1962
rect 13288 1930 13320 1962
rect 13356 1930 13388 1962
rect 13424 1930 13456 1962
rect 13492 1930 13524 1962
rect 13560 1930 13592 1962
rect 13628 1930 13660 1962
rect 13696 1930 13728 1962
rect 13764 1930 13796 1962
rect 13832 1930 13864 1962
rect 13900 1930 13932 1962
rect 13968 1930 14000 1962
rect 14036 1930 14068 1962
rect 14104 1930 14136 1962
rect 14172 1930 14204 1962
rect 14240 1930 14272 1962
rect 14308 1930 14340 1962
rect 14376 1930 14408 1962
rect 14444 1930 14476 1962
rect 14512 1930 14544 1962
rect 14580 1930 14612 1962
rect 14648 1930 14680 1962
rect 14716 1930 14748 1962
rect 14784 1930 14816 1962
rect 14852 1930 14884 1962
rect 14920 1930 14952 1962
rect 14988 1930 15020 1962
rect 15056 1930 15088 1962
rect 15124 1930 15156 1962
rect 15192 1930 15224 1962
rect 15260 1930 15292 1962
rect 15328 1930 15360 1962
rect 15396 1930 15428 1962
rect 15464 1930 15496 1962
rect 15532 1930 15564 1962
rect 15600 1930 15632 1962
rect 15668 1930 15700 1962
rect 15736 1930 15768 1962
rect 15804 1930 15836 1962
rect 15872 1930 15904 1962
rect 15940 1930 15972 1962
rect 18 1824 50 1856
rect 18 1756 50 1788
rect 18 1688 50 1720
rect 18 1620 50 1652
rect 15950 1824 15982 1856
rect 15950 1756 15982 1788
rect 15950 1688 15982 1720
rect 18 1552 50 1584
rect 18 1484 50 1516
rect 18 1416 50 1448
rect 18 1348 50 1380
rect 18 1280 50 1312
rect 18 1212 50 1244
rect 18 1144 50 1176
rect 18 1076 50 1108
rect 18 1008 50 1040
rect 18 940 50 972
rect 18 872 50 904
rect 18 804 50 836
rect 18 736 50 768
rect 18 668 50 700
rect 18 600 50 632
rect 18 532 50 564
rect 18 464 50 496
rect 18 396 50 428
rect 15950 1620 15982 1652
rect 15950 1552 15982 1584
rect 15950 1484 15982 1516
rect 15950 1416 15982 1448
rect 15950 1348 15982 1380
rect 15950 1280 15982 1312
rect 15950 1212 15982 1244
rect 15950 1144 15982 1176
rect 15950 1076 15982 1108
rect 15950 1008 15982 1040
rect 15950 940 15982 972
rect 15950 872 15982 904
rect 15950 804 15982 836
rect 15950 736 15982 768
rect 15950 668 15982 700
rect 15950 600 15982 632
rect 15950 532 15982 564
rect 15950 464 15982 496
rect 15950 396 15982 428
rect 18 328 50 360
rect 18 260 50 292
rect 18 192 50 224
rect 18 124 50 156
rect 15950 328 15982 360
rect 15950 260 15982 292
rect 15950 192 15982 224
rect 15950 124 15982 156
rect 28 18 60 50
rect 96 18 128 50
rect 164 18 196 50
rect 232 18 264 50
rect 300 18 332 50
rect 368 18 400 50
rect 436 18 468 50
rect 504 18 536 50
rect 572 18 604 50
rect 640 18 672 50
rect 708 18 740 50
rect 776 18 808 50
rect 844 18 876 50
rect 912 18 944 50
rect 980 18 1012 50
rect 1048 18 1080 50
rect 1116 18 1148 50
rect 1184 18 1216 50
rect 1252 18 1284 50
rect 1320 18 1352 50
rect 1388 18 1420 50
rect 1456 18 1488 50
rect 1524 18 1556 50
rect 1592 18 1624 50
rect 1660 18 1692 50
rect 1728 18 1760 50
rect 1796 18 1828 50
rect 1864 18 1896 50
rect 1932 18 1964 50
rect 2000 18 2032 50
rect 2068 18 2100 50
rect 2136 18 2168 50
rect 2204 18 2236 50
rect 2272 18 2304 50
rect 2340 18 2372 50
rect 2408 18 2440 50
rect 2476 18 2508 50
rect 2544 18 2576 50
rect 2612 18 2644 50
rect 2680 18 2712 50
rect 2748 18 2780 50
rect 2816 18 2848 50
rect 2884 18 2916 50
rect 2952 18 2984 50
rect 3020 18 3052 50
rect 3088 18 3120 50
rect 3156 18 3188 50
rect 3224 18 3256 50
rect 3292 18 3324 50
rect 3360 18 3392 50
rect 3428 18 3460 50
rect 3496 18 3528 50
rect 3564 18 3596 50
rect 3632 18 3664 50
rect 3700 18 3732 50
rect 3768 18 3800 50
rect 3836 18 3868 50
rect 3904 18 3936 50
rect 3972 18 4004 50
rect 4040 18 4072 50
rect 4108 18 4140 50
rect 4176 18 4208 50
rect 4244 18 4276 50
rect 4312 18 4344 50
rect 4380 18 4412 50
rect 4448 18 4480 50
rect 4516 18 4548 50
rect 4584 18 4616 50
rect 4652 18 4684 50
rect 4720 18 4752 50
rect 4788 18 4820 50
rect 4856 18 4888 50
rect 4924 18 4956 50
rect 4992 18 5024 50
rect 5060 18 5092 50
rect 5128 18 5160 50
rect 5196 18 5228 50
rect 5264 18 5296 50
rect 5332 18 5364 50
rect 5400 18 5432 50
rect 5468 18 5500 50
rect 5536 18 5568 50
rect 5604 18 5636 50
rect 5672 18 5704 50
rect 5740 18 5772 50
rect 5808 18 5840 50
rect 5876 18 5908 50
rect 5944 18 5976 50
rect 6012 18 6044 50
rect 6080 18 6112 50
rect 6148 18 6180 50
rect 6216 18 6248 50
rect 6284 18 6316 50
rect 6352 18 6384 50
rect 6420 18 6452 50
rect 6488 18 6520 50
rect 6556 18 6588 50
rect 6624 18 6656 50
rect 6692 18 6724 50
rect 6760 18 6792 50
rect 6828 18 6860 50
rect 6896 18 6928 50
rect 6964 18 6996 50
rect 7032 18 7064 50
rect 7100 18 7132 50
rect 7168 18 7200 50
rect 7236 18 7268 50
rect 7304 18 7336 50
rect 7372 18 7404 50
rect 7440 18 7472 50
rect 7508 18 7540 50
rect 7576 18 7608 50
rect 7644 18 7676 50
rect 7712 18 7744 50
rect 7780 18 7812 50
rect 7848 18 7880 50
rect 7916 18 7948 50
rect 7984 18 8016 50
rect 8052 18 8084 50
rect 8120 18 8152 50
rect 8188 18 8220 50
rect 8256 18 8288 50
rect 8324 18 8356 50
rect 8392 18 8424 50
rect 8460 18 8492 50
rect 8528 18 8560 50
rect 8596 18 8628 50
rect 8664 18 8696 50
rect 8732 18 8764 50
rect 8800 18 8832 50
rect 8868 18 8900 50
rect 8936 18 8968 50
rect 9004 18 9036 50
rect 9072 18 9104 50
rect 9140 18 9172 50
rect 9208 18 9240 50
rect 9276 18 9308 50
rect 9344 18 9376 50
rect 9412 18 9444 50
rect 9480 18 9512 50
rect 9548 18 9580 50
rect 9616 18 9648 50
rect 9684 18 9716 50
rect 9752 18 9784 50
rect 9820 18 9852 50
rect 9888 18 9920 50
rect 9956 18 9988 50
rect 10024 18 10056 50
rect 10092 18 10124 50
rect 10160 18 10192 50
rect 10228 18 10260 50
rect 10296 18 10328 50
rect 10364 18 10396 50
rect 10432 18 10464 50
rect 10500 18 10532 50
rect 10568 18 10600 50
rect 10636 18 10668 50
rect 10704 18 10736 50
rect 10772 18 10804 50
rect 10840 18 10872 50
rect 10908 18 10940 50
rect 10976 18 11008 50
rect 11044 18 11076 50
rect 11112 18 11144 50
rect 11180 18 11212 50
rect 11248 18 11280 50
rect 11316 18 11348 50
rect 11384 18 11416 50
rect 11452 18 11484 50
rect 11520 18 11552 50
rect 11588 18 11620 50
rect 11656 18 11688 50
rect 11724 18 11756 50
rect 11792 18 11824 50
rect 11860 18 11892 50
rect 11928 18 11960 50
rect 11996 18 12028 50
rect 12064 18 12096 50
rect 12132 18 12164 50
rect 12200 18 12232 50
rect 12268 18 12300 50
rect 12336 18 12368 50
rect 12404 18 12436 50
rect 12472 18 12504 50
rect 12540 18 12572 50
rect 12608 18 12640 50
rect 12676 18 12708 50
rect 12744 18 12776 50
rect 12812 18 12844 50
rect 12880 18 12912 50
rect 12948 18 12980 50
rect 13016 18 13048 50
rect 13084 18 13116 50
rect 13152 18 13184 50
rect 13220 18 13252 50
rect 13288 18 13320 50
rect 13356 18 13388 50
rect 13424 18 13456 50
rect 13492 18 13524 50
rect 13560 18 13592 50
rect 13628 18 13660 50
rect 13696 18 13728 50
rect 13764 18 13796 50
rect 13832 18 13864 50
rect 13900 18 13932 50
rect 13968 18 14000 50
rect 14036 18 14068 50
rect 14104 18 14136 50
rect 14172 18 14204 50
rect 14240 18 14272 50
rect 14308 18 14340 50
rect 14376 18 14408 50
rect 14444 18 14476 50
rect 14512 18 14544 50
rect 14580 18 14612 50
rect 14648 18 14680 50
rect 14716 18 14748 50
rect 14784 18 14816 50
rect 14852 18 14884 50
rect 14920 18 14952 50
rect 14988 18 15020 50
rect 15056 18 15088 50
rect 15124 18 15156 50
rect 15192 18 15224 50
rect 15260 18 15292 50
rect 15328 18 15360 50
rect 15396 18 15428 50
rect 15464 18 15496 50
rect 15532 18 15564 50
rect 15600 18 15632 50
rect 15668 18 15700 50
rect 15736 18 15768 50
rect 15804 18 15836 50
rect 15872 18 15904 50
rect 15940 18 15972 50
<< poly >>
rect 5044 1490 5164 1504
rect 5044 1458 5088 1490
rect 5120 1458 5164 1490
rect 5044 1430 5164 1458
rect 5400 1490 5520 1504
rect 5400 1458 5444 1490
rect 5476 1458 5520 1490
rect 5400 1430 5520 1458
rect 5648 1490 5768 1504
rect 5648 1458 5692 1490
rect 5724 1458 5768 1490
rect 5648 1430 5768 1458
rect 6004 1490 6124 1504
rect 6004 1458 6048 1490
rect 6080 1458 6124 1490
rect 6004 1430 6124 1458
rect 6252 1490 6372 1504
rect 6252 1458 6296 1490
rect 6328 1458 6372 1490
rect 6252 1430 6372 1458
rect 6608 1490 6728 1504
rect 6608 1458 6652 1490
rect 6684 1458 6728 1490
rect 6608 1430 6728 1458
rect 6856 1490 6976 1504
rect 6856 1458 6900 1490
rect 6932 1458 6976 1490
rect 6856 1430 6976 1458
rect 7212 1490 7332 1504
rect 7212 1458 7256 1490
rect 7288 1458 7332 1490
rect 7212 1430 7332 1458
rect 7460 1490 7580 1504
rect 7460 1458 7504 1490
rect 7536 1458 7580 1490
rect 7460 1430 7580 1458
rect 7816 1490 7936 1504
rect 7816 1458 7860 1490
rect 7892 1458 7936 1490
rect 7816 1430 7936 1458
rect 8064 1490 8184 1504
rect 8064 1458 8108 1490
rect 8140 1458 8184 1490
rect 8064 1430 8184 1458
rect 8420 1490 8540 1504
rect 8420 1458 8464 1490
rect 8496 1458 8540 1490
rect 8420 1430 8540 1458
rect 8668 1490 8788 1504
rect 8668 1458 8712 1490
rect 8744 1458 8788 1490
rect 8668 1430 8788 1458
rect 9024 1490 9144 1504
rect 9024 1458 9068 1490
rect 9100 1458 9144 1490
rect 9024 1430 9144 1458
rect 9272 1490 9392 1504
rect 9272 1458 9316 1490
rect 9348 1458 9392 1490
rect 9272 1430 9392 1458
rect 9628 1490 9748 1504
rect 9628 1458 9672 1490
rect 9704 1458 9748 1490
rect 9628 1430 9748 1458
rect 9876 1490 9996 1504
rect 9876 1458 9920 1490
rect 9952 1458 9996 1490
rect 9876 1430 9996 1458
rect 10232 1490 10352 1504
rect 10232 1458 10276 1490
rect 10308 1458 10352 1490
rect 10232 1430 10352 1458
rect 10480 1490 10600 1504
rect 10480 1458 10524 1490
rect 10556 1458 10600 1490
rect 10480 1430 10600 1458
rect 10836 1490 10956 1504
rect 10836 1458 10880 1490
rect 10912 1458 10956 1490
rect 10836 1430 10956 1458
rect 13261 1416 13361 1430
rect 13261 1384 13275 1416
rect 13347 1384 13361 1416
rect 13261 1344 13361 1384
rect 13261 596 13361 636
rect 13261 564 13275 596
rect 13347 564 13361 596
rect 13261 550 13361 564
rect 5044 522 5164 550
rect 5044 490 5088 522
rect 5120 490 5164 522
rect 5044 476 5164 490
rect 5400 522 5520 550
rect 5400 490 5444 522
rect 5476 490 5520 522
rect 5400 476 5520 490
rect 5648 522 5768 550
rect 5648 490 5692 522
rect 5724 490 5768 522
rect 5648 476 5768 490
rect 6004 522 6124 550
rect 6004 490 6048 522
rect 6080 490 6124 522
rect 6004 476 6124 490
rect 6252 522 6372 550
rect 6252 490 6296 522
rect 6328 490 6372 522
rect 6252 476 6372 490
rect 6608 522 6728 550
rect 6608 490 6652 522
rect 6684 490 6728 522
rect 6608 476 6728 490
rect 6856 522 6976 550
rect 6856 490 6900 522
rect 6932 490 6976 522
rect 6856 476 6976 490
rect 7212 522 7332 550
rect 7212 490 7256 522
rect 7288 490 7332 522
rect 7212 476 7332 490
rect 7460 522 7580 550
rect 7460 490 7504 522
rect 7536 490 7580 522
rect 7460 476 7580 490
rect 7816 522 7936 550
rect 7816 490 7860 522
rect 7892 490 7936 522
rect 7816 476 7936 490
rect 8064 522 8184 550
rect 8064 490 8108 522
rect 8140 490 8184 522
rect 8064 476 8184 490
rect 8420 522 8540 550
rect 8420 490 8464 522
rect 8496 490 8540 522
rect 8420 476 8540 490
rect 8668 522 8788 550
rect 8668 490 8712 522
rect 8744 490 8788 522
rect 8668 476 8788 490
rect 9024 522 9144 550
rect 9024 490 9068 522
rect 9100 490 9144 522
rect 9024 476 9144 490
rect 9272 522 9392 550
rect 9272 490 9316 522
rect 9348 490 9392 522
rect 9272 476 9392 490
rect 9628 522 9748 550
rect 9628 490 9672 522
rect 9704 490 9748 522
rect 9628 476 9748 490
rect 9876 522 9996 550
rect 9876 490 9920 522
rect 9952 490 9996 522
rect 9876 476 9996 490
rect 10232 522 10352 550
rect 10232 490 10276 522
rect 10308 490 10352 522
rect 10232 476 10352 490
rect 10480 522 10600 550
rect 10480 490 10524 522
rect 10556 490 10600 522
rect 10480 476 10600 490
rect 10836 522 10956 550
rect 10836 490 10880 522
rect 10912 490 10956 522
rect 10836 476 10956 490
<< polycont >>
rect 5088 1458 5120 1490
rect 5444 1458 5476 1490
rect 5692 1458 5724 1490
rect 6048 1458 6080 1490
rect 6296 1458 6328 1490
rect 6652 1458 6684 1490
rect 6900 1458 6932 1490
rect 7256 1458 7288 1490
rect 7504 1458 7536 1490
rect 7860 1458 7892 1490
rect 8108 1458 8140 1490
rect 8464 1458 8496 1490
rect 8712 1458 8744 1490
rect 9068 1458 9100 1490
rect 9316 1458 9348 1490
rect 9672 1458 9704 1490
rect 9920 1458 9952 1490
rect 10276 1458 10308 1490
rect 10524 1458 10556 1490
rect 10880 1458 10912 1490
rect 13275 1384 13347 1416
rect 13275 564 13347 596
rect 5088 490 5120 522
rect 5444 490 5476 522
rect 5692 490 5724 522
rect 6048 490 6080 522
rect 6296 490 6328 522
rect 6652 490 6684 522
rect 6900 490 6932 522
rect 7256 490 7288 522
rect 7504 490 7536 522
rect 7860 490 7892 522
rect 8108 490 8140 522
rect 8464 490 8496 522
rect 8712 490 8744 522
rect 9068 490 9100 522
rect 9316 490 9348 522
rect 9672 490 9704 522
rect 9920 490 9952 522
rect 10276 490 10308 522
rect 10524 490 10556 522
rect 10880 490 10912 522
<< ppolyres >>
rect 13261 636 13361 1344
<< metal1 >>
rect 0 1979 9416 1980
rect 9587 1979 16000 1980
rect 0 1962 16000 1979
rect 0 1930 28 1962
rect 60 1930 96 1962
rect 128 1930 164 1962
rect 196 1930 232 1962
rect 264 1930 300 1962
rect 332 1930 368 1962
rect 400 1930 436 1962
rect 468 1930 504 1962
rect 536 1930 572 1962
rect 604 1930 640 1962
rect 672 1930 708 1962
rect 740 1930 776 1962
rect 808 1930 844 1962
rect 876 1930 912 1962
rect 944 1930 980 1962
rect 1012 1930 1048 1962
rect 1080 1930 1116 1962
rect 1148 1930 1184 1962
rect 1216 1930 1252 1962
rect 1284 1930 1320 1962
rect 1352 1930 1388 1962
rect 1420 1930 1456 1962
rect 1488 1930 1524 1962
rect 1556 1930 1592 1962
rect 1624 1930 1660 1962
rect 1692 1930 1728 1962
rect 1760 1930 1796 1962
rect 1828 1930 1864 1962
rect 1896 1930 1932 1962
rect 1964 1930 2000 1962
rect 2032 1930 2068 1962
rect 2100 1930 2136 1962
rect 2168 1930 2204 1962
rect 2236 1930 2272 1962
rect 2304 1930 2340 1962
rect 2372 1930 2408 1962
rect 2440 1930 2476 1962
rect 2508 1930 2544 1962
rect 2576 1930 2612 1962
rect 2644 1930 2680 1962
rect 2712 1930 2748 1962
rect 2780 1930 2816 1962
rect 2848 1930 2884 1962
rect 2916 1930 2952 1962
rect 2984 1930 3020 1962
rect 3052 1930 3088 1962
rect 3120 1930 3156 1962
rect 3188 1930 3224 1962
rect 3256 1930 3292 1962
rect 3324 1930 3360 1962
rect 3392 1930 3428 1962
rect 3460 1930 3496 1962
rect 3528 1930 3564 1962
rect 3596 1930 3632 1962
rect 3664 1930 3700 1962
rect 3732 1930 3768 1962
rect 3800 1930 3836 1962
rect 3868 1930 3904 1962
rect 3936 1930 3972 1962
rect 4004 1930 4040 1962
rect 4072 1930 4108 1962
rect 4140 1930 4176 1962
rect 4208 1930 4244 1962
rect 4276 1930 4312 1962
rect 4344 1930 4380 1962
rect 4412 1930 4448 1962
rect 4480 1930 4516 1962
rect 4548 1930 4584 1962
rect 4616 1930 4652 1962
rect 4684 1930 4720 1962
rect 4752 1930 4788 1962
rect 4820 1930 4856 1962
rect 4888 1930 4924 1962
rect 4956 1930 4992 1962
rect 5024 1930 5060 1962
rect 5092 1930 5128 1962
rect 5160 1930 5196 1962
rect 5228 1930 5264 1962
rect 5296 1930 5332 1962
rect 5364 1930 5400 1962
rect 5432 1930 5468 1962
rect 5500 1930 5536 1962
rect 5568 1930 5604 1962
rect 5636 1930 5672 1962
rect 5704 1930 5740 1962
rect 5772 1930 5808 1962
rect 5840 1930 5876 1962
rect 5908 1930 5944 1962
rect 5976 1930 6012 1962
rect 6044 1930 6080 1962
rect 6112 1930 6148 1962
rect 6180 1930 6216 1962
rect 6248 1930 6284 1962
rect 6316 1930 6352 1962
rect 6384 1930 6420 1962
rect 6452 1930 6488 1962
rect 6520 1930 6556 1962
rect 6588 1930 6624 1962
rect 6656 1930 6692 1962
rect 6724 1930 6760 1962
rect 6792 1930 6828 1962
rect 6860 1930 6896 1962
rect 6928 1930 6964 1962
rect 6996 1930 7032 1962
rect 7064 1930 7100 1962
rect 7132 1930 7168 1962
rect 7200 1930 7236 1962
rect 7268 1930 7304 1962
rect 7336 1930 7372 1962
rect 7404 1930 7440 1962
rect 7472 1930 7508 1962
rect 7540 1930 7576 1962
rect 7608 1930 7644 1962
rect 7676 1930 7712 1962
rect 7744 1930 7780 1962
rect 7812 1930 7848 1962
rect 7880 1930 7916 1962
rect 7948 1930 7984 1962
rect 8016 1930 8052 1962
rect 8084 1930 8120 1962
rect 8152 1930 8188 1962
rect 8220 1930 8256 1962
rect 8288 1930 8324 1962
rect 8356 1930 8392 1962
rect 8424 1930 8460 1962
rect 8492 1930 8528 1962
rect 8560 1930 8596 1962
rect 8628 1930 8664 1962
rect 8696 1930 8732 1962
rect 8764 1930 8800 1962
rect 8832 1930 8868 1962
rect 8900 1930 8936 1962
rect 8968 1930 9004 1962
rect 9036 1930 9072 1962
rect 9104 1930 9140 1962
rect 9172 1930 9208 1962
rect 9240 1930 9276 1962
rect 9308 1930 9344 1962
rect 9376 1930 9412 1962
rect 9444 1930 9480 1962
rect 9512 1930 9548 1962
rect 9580 1930 9616 1962
rect 9648 1930 9684 1962
rect 9716 1930 9752 1962
rect 9784 1930 9820 1962
rect 9852 1930 9888 1962
rect 9920 1930 9956 1962
rect 9988 1930 10024 1962
rect 10056 1930 10092 1962
rect 10124 1930 10160 1962
rect 10192 1930 10228 1962
rect 10260 1930 10296 1962
rect 10328 1930 10364 1962
rect 10396 1930 10432 1962
rect 10464 1930 10500 1962
rect 10532 1930 10568 1962
rect 10600 1930 10636 1962
rect 10668 1930 10704 1962
rect 10736 1930 10772 1962
rect 10804 1930 10840 1962
rect 10872 1930 10908 1962
rect 10940 1930 10976 1962
rect 11008 1930 11044 1962
rect 11076 1930 11112 1962
rect 11144 1930 11180 1962
rect 11212 1930 11248 1962
rect 11280 1930 11316 1962
rect 11348 1930 11384 1962
rect 11416 1930 11452 1962
rect 11484 1930 11520 1962
rect 11552 1930 11588 1962
rect 11620 1930 11656 1962
rect 11688 1930 11724 1962
rect 11756 1930 11792 1962
rect 11824 1930 11860 1962
rect 11892 1930 11928 1962
rect 11960 1930 11996 1962
rect 12028 1930 12064 1962
rect 12096 1930 12132 1962
rect 12164 1930 12200 1962
rect 12232 1930 12268 1962
rect 12300 1930 12336 1962
rect 12368 1930 12404 1962
rect 12436 1930 12472 1962
rect 12504 1930 12540 1962
rect 12572 1930 12608 1962
rect 12640 1930 12676 1962
rect 12708 1930 12744 1962
rect 12776 1930 12812 1962
rect 12844 1930 12880 1962
rect 12912 1930 12948 1962
rect 12980 1930 13016 1962
rect 13048 1930 13084 1962
rect 13116 1930 13152 1962
rect 13184 1930 13220 1962
rect 13252 1930 13288 1962
rect 13320 1930 13356 1962
rect 13388 1930 13424 1962
rect 13456 1930 13492 1962
rect 13524 1930 13560 1962
rect 13592 1930 13628 1962
rect 13660 1930 13696 1962
rect 13728 1930 13764 1962
rect 13796 1930 13832 1962
rect 13864 1930 13900 1962
rect 13932 1930 13968 1962
rect 14000 1930 14036 1962
rect 14068 1930 14104 1962
rect 14136 1930 14172 1962
rect 14204 1930 14240 1962
rect 14272 1930 14308 1962
rect 14340 1930 14376 1962
rect 14408 1930 14444 1962
rect 14476 1930 14512 1962
rect 14544 1930 14580 1962
rect 14612 1930 14648 1962
rect 14680 1930 14716 1962
rect 14748 1930 14784 1962
rect 14816 1930 14852 1962
rect 14884 1930 14920 1962
rect 14952 1930 14988 1962
rect 15020 1930 15056 1962
rect 15088 1930 15124 1962
rect 15156 1930 15192 1962
rect 15224 1930 15260 1962
rect 15292 1930 15328 1962
rect 15360 1930 15396 1962
rect 15428 1930 15464 1962
rect 15496 1930 15532 1962
rect 15564 1930 15600 1962
rect 15632 1930 15668 1962
rect 15700 1930 15736 1962
rect 15768 1930 15804 1962
rect 15836 1930 15872 1962
rect 15904 1930 15940 1962
rect 15972 1930 16000 1962
rect 0 1912 16000 1930
rect 0 1856 68 1912
rect 0 1824 18 1856
rect 50 1824 68 1856
rect 0 1788 68 1824
rect 0 1756 18 1788
rect 50 1756 68 1788
rect 0 1720 68 1756
rect 0 1688 18 1720
rect 50 1688 68 1720
rect 0 1652 68 1688
rect 0 1620 18 1652
rect 50 1620 68 1652
rect 15932 1856 16000 1912
rect 15932 1824 15950 1856
rect 15982 1824 16000 1856
rect 15932 1788 16000 1824
rect 15932 1756 15950 1788
rect 15982 1756 16000 1788
rect 15932 1720 16000 1756
rect 15932 1688 15950 1720
rect 15982 1688 16000 1720
rect 15932 1652 16000 1688
rect 0 1584 68 1620
rect 0 1552 18 1584
rect 50 1552 68 1584
rect 0 1516 68 1552
rect 0 1484 18 1516
rect 50 1484 68 1516
rect 0 1448 68 1484
rect 0 1416 18 1448
rect 50 1416 68 1448
rect 0 1380 68 1416
rect 0 1348 18 1380
rect 50 1348 68 1380
rect 0 1312 68 1348
rect 0 1280 18 1312
rect 50 1280 68 1312
rect 0 1244 68 1280
rect 0 1212 18 1244
rect 50 1212 68 1244
rect 0 1176 68 1212
rect 0 1144 18 1176
rect 50 1144 68 1176
rect 0 1108 68 1144
rect 0 1076 18 1108
rect 50 1076 68 1108
rect 0 1040 68 1076
rect 0 1008 18 1040
rect 50 1008 68 1040
rect 0 972 68 1008
rect 0 940 18 972
rect 50 940 68 972
rect 0 904 68 940
rect 0 872 18 904
rect 50 872 68 904
rect 0 836 68 872
rect 0 804 18 836
rect 50 804 68 836
rect 0 768 68 804
rect 0 736 18 768
rect 50 736 68 768
rect 0 700 68 736
rect 0 668 18 700
rect 50 668 68 700
rect 0 632 68 668
rect 0 600 18 632
rect 50 600 68 632
rect 0 564 68 600
rect 0 532 18 564
rect 50 532 68 564
rect 0 496 68 532
rect 0 464 18 496
rect 50 464 68 496
rect 0 428 68 464
rect 0 396 18 428
rect 50 396 68 428
rect 0 360 68 396
rect 360 1612 15640 1630
rect 360 1580 402 1612
rect 434 1580 470 1612
rect 502 1580 538 1612
rect 570 1580 606 1612
rect 638 1580 674 1612
rect 706 1580 742 1612
rect 774 1580 810 1612
rect 842 1580 878 1612
rect 910 1580 946 1612
rect 978 1580 1014 1612
rect 1046 1580 1082 1612
rect 1114 1580 1150 1612
rect 1182 1580 1218 1612
rect 1250 1580 1286 1612
rect 1318 1580 1354 1612
rect 1386 1580 1422 1612
rect 1454 1580 1490 1612
rect 1522 1580 1558 1612
rect 1590 1580 1626 1612
rect 1658 1580 1694 1612
rect 1726 1580 1762 1612
rect 1794 1580 1830 1612
rect 1862 1580 1898 1612
rect 1930 1580 1966 1612
rect 1998 1580 2034 1612
rect 2066 1580 2102 1612
rect 2134 1580 2170 1612
rect 2202 1580 2238 1612
rect 2270 1580 2306 1612
rect 2338 1580 2374 1612
rect 2406 1580 2442 1612
rect 2474 1580 2510 1612
rect 2542 1580 2578 1612
rect 2610 1580 2646 1612
rect 2678 1580 2714 1612
rect 2746 1580 2782 1612
rect 2814 1580 2850 1612
rect 2882 1580 2918 1612
rect 2950 1580 2986 1612
rect 3018 1580 3054 1612
rect 3086 1580 3122 1612
rect 3154 1580 3190 1612
rect 3222 1580 3258 1612
rect 3290 1580 3326 1612
rect 3358 1580 3394 1612
rect 3426 1580 3462 1612
rect 3494 1580 3530 1612
rect 3562 1580 3598 1612
rect 3630 1580 3666 1612
rect 3698 1580 3734 1612
rect 3766 1580 3802 1612
rect 3834 1580 3870 1612
rect 3902 1580 3938 1612
rect 3970 1580 4006 1612
rect 4038 1580 4074 1612
rect 4106 1580 4142 1612
rect 4174 1580 4210 1612
rect 4242 1580 4278 1612
rect 4310 1580 4346 1612
rect 4378 1580 4414 1612
rect 4446 1580 4482 1612
rect 4514 1580 4550 1612
rect 4582 1580 4618 1612
rect 4650 1580 4686 1612
rect 4718 1580 4754 1612
rect 4786 1580 4822 1612
rect 4854 1580 4890 1612
rect 4922 1580 4958 1612
rect 4990 1606 5026 1612
rect 5000 1580 5026 1606
rect 5058 1580 5094 1612
rect 5126 1580 5162 1612
rect 5194 1580 5230 1612
rect 5262 1580 5298 1612
rect 5330 1580 5366 1612
rect 5398 1580 5434 1612
rect 5466 1580 5502 1612
rect 5534 1606 5570 1612
rect 5602 1606 5638 1612
rect 5534 1580 5564 1606
rect 5604 1580 5638 1606
rect 5670 1580 5706 1612
rect 5738 1580 5774 1612
rect 5806 1580 5842 1612
rect 5874 1580 5910 1612
rect 5942 1580 5978 1612
rect 6010 1580 6046 1612
rect 6078 1580 6114 1612
rect 6146 1606 6182 1612
rect 6146 1580 6168 1606
rect 6214 1580 6250 1612
rect 6282 1580 6318 1612
rect 6350 1580 6386 1612
rect 6418 1580 6454 1612
rect 6486 1580 6522 1612
rect 6554 1580 6590 1612
rect 6622 1580 6658 1612
rect 6690 1580 6726 1612
rect 6758 1606 6794 1612
rect 6758 1580 6772 1606
rect 6826 1580 6862 1612
rect 6894 1580 6930 1612
rect 6962 1580 6998 1612
rect 7030 1580 7066 1612
rect 7098 1580 7134 1612
rect 7166 1580 7202 1612
rect 7234 1580 7270 1612
rect 7302 1580 7338 1612
rect 7370 1606 7406 1612
rect 7370 1580 7376 1606
rect 7438 1580 7474 1612
rect 7506 1580 7542 1612
rect 7574 1580 7610 1612
rect 7642 1580 7678 1612
rect 7710 1580 7746 1612
rect 7778 1580 7814 1612
rect 7846 1580 7882 1612
rect 7914 1580 7950 1612
rect 7982 1606 8018 1612
rect 8050 1580 8086 1612
rect 8118 1580 8154 1612
rect 8186 1580 8222 1612
rect 8254 1580 8290 1612
rect 8322 1580 8358 1612
rect 8390 1580 8426 1612
rect 8458 1580 8494 1612
rect 8526 1580 8562 1612
rect 8594 1606 8630 1612
rect 8624 1580 8630 1606
rect 8662 1580 8698 1612
rect 8730 1580 8766 1612
rect 8798 1580 8834 1612
rect 8866 1580 8902 1612
rect 8934 1580 8970 1612
rect 9002 1580 9038 1612
rect 9070 1580 9106 1612
rect 9138 1580 9174 1612
rect 9206 1606 9242 1612
rect 9228 1580 9242 1606
rect 9274 1580 9310 1612
rect 9342 1580 9378 1612
rect 9410 1580 9446 1612
rect 9478 1580 9514 1612
rect 9546 1580 9582 1612
rect 9614 1580 9650 1612
rect 9682 1580 9718 1612
rect 9750 1580 9786 1612
rect 9818 1606 9854 1612
rect 9832 1580 9854 1606
rect 9886 1580 9922 1612
rect 9954 1580 9990 1612
rect 10022 1580 10058 1612
rect 10090 1580 10126 1612
rect 10158 1580 10194 1612
rect 10226 1580 10262 1612
rect 10294 1580 10330 1612
rect 10362 1606 10398 1612
rect 10430 1606 10466 1612
rect 10362 1580 10396 1606
rect 10436 1580 10466 1606
rect 10498 1580 10534 1612
rect 10566 1580 10602 1612
rect 10634 1580 10670 1612
rect 10702 1580 10738 1612
rect 10770 1580 10806 1612
rect 10838 1580 10874 1612
rect 10906 1580 10942 1612
rect 10974 1606 11010 1612
rect 10974 1580 11000 1606
rect 11042 1580 11078 1612
rect 11110 1580 11146 1612
rect 11178 1580 11214 1612
rect 11246 1580 11282 1612
rect 11314 1580 11350 1612
rect 11382 1580 11418 1612
rect 11450 1580 11486 1612
rect 11518 1580 11554 1612
rect 11586 1580 11622 1612
rect 11654 1580 11690 1612
rect 11722 1580 11758 1612
rect 11790 1580 11826 1612
rect 11858 1580 11894 1612
rect 11926 1580 11962 1612
rect 11994 1580 12030 1612
rect 12062 1580 12098 1612
rect 12130 1580 12166 1612
rect 12198 1580 12234 1612
rect 12266 1580 12302 1612
rect 12334 1580 12370 1612
rect 12402 1580 12438 1612
rect 12470 1580 12506 1612
rect 12538 1580 12574 1612
rect 12606 1580 12642 1612
rect 12674 1580 12710 1612
rect 12742 1580 12778 1612
rect 12810 1580 12846 1612
rect 12878 1580 12914 1612
rect 12946 1580 12982 1612
rect 13014 1580 13050 1612
rect 13082 1580 13118 1612
rect 13150 1580 13186 1612
rect 13218 1580 13254 1612
rect 13286 1580 13322 1612
rect 13354 1580 13390 1612
rect 13422 1580 13458 1612
rect 13490 1580 13526 1612
rect 13558 1580 13594 1612
rect 13626 1580 13662 1612
rect 13694 1580 13730 1612
rect 13762 1580 13798 1612
rect 13830 1580 13866 1612
rect 13898 1580 13934 1612
rect 13966 1580 14002 1612
rect 14034 1580 14070 1612
rect 14102 1580 14138 1612
rect 14170 1580 14206 1612
rect 14238 1580 14274 1612
rect 14306 1580 14342 1612
rect 14374 1580 14410 1612
rect 14442 1580 14478 1612
rect 14510 1580 14546 1612
rect 14578 1580 14614 1612
rect 14646 1580 14682 1612
rect 14714 1580 14750 1612
rect 14782 1580 14818 1612
rect 14850 1580 14886 1612
rect 14918 1580 14954 1612
rect 14986 1580 15022 1612
rect 15054 1580 15090 1612
rect 15122 1580 15158 1612
rect 15190 1580 15226 1612
rect 15258 1580 15294 1612
rect 15326 1580 15362 1612
rect 15394 1580 15430 1612
rect 15462 1580 15498 1612
rect 15530 1580 15566 1612
rect 15598 1580 15640 1612
rect 360 1566 4960 1580
rect 5000 1566 5564 1580
rect 5604 1566 6168 1580
rect 6208 1566 6772 1580
rect 6812 1566 7376 1580
rect 7416 1566 7980 1580
rect 8020 1566 8584 1580
rect 8624 1566 9188 1580
rect 9228 1566 9792 1580
rect 9832 1566 10396 1580
rect 10436 1566 11000 1580
rect 11040 1566 15640 1580
rect 360 1562 15640 1566
rect 360 1526 428 1562
rect 4959 1552 5001 1562
rect 5563 1552 5605 1562
rect 6167 1552 6209 1562
rect 6771 1552 6813 1562
rect 7375 1552 7417 1562
rect 7979 1552 8021 1562
rect 8583 1552 8625 1562
rect 9187 1552 9229 1562
rect 9791 1552 9833 1562
rect 10395 1552 10437 1562
rect 10999 1552 11041 1562
rect 360 1494 378 1526
rect 410 1494 428 1526
rect 15572 1526 15640 1562
rect 360 1458 428 1494
rect 360 1426 378 1458
rect 410 1426 428 1458
rect 5088 1490 13327 1506
rect 5120 1474 5444 1490
rect 360 1390 428 1426
rect 360 1358 378 1390
rect 410 1358 428 1390
rect 360 1322 428 1358
rect 360 1290 378 1322
rect 410 1290 428 1322
rect 360 1254 428 1290
rect 360 1222 378 1254
rect 410 1222 428 1254
rect 360 1186 428 1222
rect 360 1154 378 1186
rect 410 1154 428 1186
rect 360 1118 428 1154
rect 360 1086 378 1118
rect 410 1086 428 1118
rect 360 1050 428 1086
rect 360 1018 378 1050
rect 410 1018 428 1050
rect 360 982 428 1018
rect 360 950 378 982
rect 410 950 428 982
rect 360 914 428 950
rect 360 882 378 914
rect 410 882 428 914
rect 360 846 428 882
rect 360 814 378 846
rect 410 814 428 846
rect 360 778 428 814
rect 360 746 378 778
rect 410 746 428 778
rect 360 710 428 746
rect 360 678 378 710
rect 410 678 428 710
rect 360 642 428 678
rect 360 610 378 642
rect 410 610 428 642
rect 360 574 428 610
rect 360 542 378 574
rect 410 542 428 574
rect 4959 1420 5001 1430
rect 4959 560 4960 1420
rect 5000 560 5001 1420
rect 4959 550 5001 560
rect 360 506 428 542
rect 360 474 378 506
rect 410 474 428 506
rect 5088 522 5120 1458
rect 5476 1474 5692 1490
rect 5220 1420 5344 1430
rect 5220 560 5221 1420
rect 5343 560 5344 1420
rect 5220 550 5344 560
rect 5088 474 5120 490
rect 5444 522 5476 1458
rect 5724 1474 6048 1490
rect 5563 1420 5605 1430
rect 5563 560 5564 1420
rect 5604 560 5605 1420
rect 5563 550 5605 560
rect 5444 474 5476 490
rect 5692 522 5724 1458
rect 6080 1474 6296 1490
rect 5824 1420 5948 1430
rect 5824 560 5825 1420
rect 5947 560 5948 1420
rect 5824 550 5948 560
rect 5692 474 5724 490
rect 6048 522 6080 1458
rect 6328 1474 6652 1490
rect 6167 1420 6209 1430
rect 6167 560 6168 1420
rect 6208 560 6209 1420
rect 6167 550 6209 560
rect 6048 474 6080 490
rect 6296 522 6328 1458
rect 6684 1474 6900 1490
rect 6428 1420 6552 1430
rect 6428 560 6429 1420
rect 6551 560 6552 1420
rect 6428 550 6552 560
rect 6296 474 6328 490
rect 6652 522 6684 1458
rect 6932 1474 7256 1490
rect 6771 1420 6813 1430
rect 6771 560 6772 1420
rect 6812 560 6813 1420
rect 6771 550 6813 560
rect 6652 474 6684 490
rect 6900 522 6932 1458
rect 7288 1474 7504 1490
rect 7032 1420 7156 1430
rect 7032 560 7033 1420
rect 7155 560 7156 1420
rect 7032 550 7156 560
rect 6900 474 6932 490
rect 7256 522 7288 1458
rect 7536 1474 7860 1490
rect 7375 1420 7417 1430
rect 7375 560 7376 1420
rect 7416 560 7417 1420
rect 7375 550 7417 560
rect 7256 474 7288 490
rect 7504 522 7536 1458
rect 7892 1474 8108 1490
rect 7636 1420 7760 1430
rect 7636 560 7637 1420
rect 7759 560 7760 1420
rect 7636 550 7760 560
rect 7504 474 7536 490
rect 7860 522 7892 1458
rect 8140 1474 8464 1490
rect 7979 1420 8021 1430
rect 7979 560 7980 1420
rect 8020 560 8021 1420
rect 7979 550 8021 560
rect 7860 474 7892 490
rect 8108 522 8140 1458
rect 8496 1474 8712 1490
rect 8240 1420 8364 1430
rect 8240 560 8241 1420
rect 8363 560 8364 1420
rect 8240 550 8364 560
rect 8108 474 8140 490
rect 8464 522 8496 1458
rect 8744 1474 9068 1490
rect 8583 1420 8625 1430
rect 8583 560 8584 1420
rect 8624 560 8625 1420
rect 8583 550 8625 560
rect 8464 474 8496 490
rect 8712 522 8744 1458
rect 9100 1474 9316 1490
rect 8844 1420 8968 1430
rect 8844 560 8845 1420
rect 8967 560 8968 1420
rect 8844 550 8968 560
rect 8712 474 8744 490
rect 9068 522 9100 1458
rect 9348 1474 9672 1490
rect 9187 1420 9229 1430
rect 9187 560 9188 1420
rect 9228 560 9229 1420
rect 9187 550 9229 560
rect 9068 474 9100 490
rect 9316 522 9348 1458
rect 9704 1474 9920 1490
rect 9448 1420 9572 1430
rect 9448 560 9449 1420
rect 9571 560 9572 1420
rect 9448 550 9572 560
rect 9316 474 9348 490
rect 9672 522 9704 1458
rect 9952 1474 10276 1490
rect 9791 1420 9833 1430
rect 9791 560 9792 1420
rect 9832 560 9833 1420
rect 9791 550 9833 560
rect 9672 474 9704 490
rect 9920 522 9952 1458
rect 10308 1474 10524 1490
rect 10052 1420 10176 1430
rect 10052 560 10053 1420
rect 10175 560 10176 1420
rect 10052 550 10176 560
rect 9920 474 9952 490
rect 10276 522 10308 1458
rect 10556 1474 10880 1490
rect 10395 1420 10437 1430
rect 10395 560 10396 1420
rect 10436 560 10437 1420
rect 10395 550 10437 560
rect 10276 474 10308 490
rect 10524 522 10556 1458
rect 10912 1474 13327 1490
rect 10656 1420 10780 1430
rect 10656 560 10657 1420
rect 10779 560 10780 1420
rect 10656 550 10780 560
rect 10524 474 10556 490
rect 10880 522 10912 1458
rect 13295 1430 13327 1474
rect 15572 1494 15590 1526
rect 15622 1494 15640 1526
rect 15572 1458 15640 1494
rect 10999 1420 11041 1430
rect 10999 560 11000 1420
rect 11040 560 11041 1420
rect 13265 1416 13357 1430
rect 13265 1384 13275 1416
rect 13347 1384 13357 1416
rect 13265 1370 13357 1384
rect 15572 1426 15590 1458
rect 15622 1426 15640 1458
rect 15572 1390 15640 1426
rect 13295 1368 13327 1370
rect 15572 1358 15590 1390
rect 15622 1358 15640 1390
rect 15572 1322 15640 1358
rect 15572 1290 15590 1322
rect 15622 1290 15640 1322
rect 15572 1254 15640 1290
rect 15572 1222 15590 1254
rect 15622 1222 15640 1254
rect 15572 1186 15640 1222
rect 15572 1154 15590 1186
rect 15622 1154 15640 1186
rect 15572 1118 15640 1154
rect 15572 1086 15590 1118
rect 15622 1086 15640 1118
rect 15572 1050 15640 1086
rect 15572 1018 15590 1050
rect 15622 1018 15640 1050
rect 15572 982 15640 1018
rect 15572 950 15590 982
rect 15622 950 15640 982
rect 15572 914 15640 950
rect 15572 882 15590 914
rect 15622 882 15640 914
rect 15572 846 15640 882
rect 15572 814 15590 846
rect 15622 814 15640 846
rect 15572 778 15640 814
rect 15572 746 15590 778
rect 15622 746 15640 778
rect 15572 710 15640 746
rect 15572 678 15590 710
rect 15622 678 15640 710
rect 15572 642 15640 678
rect 15572 610 15590 642
rect 15622 610 15640 642
rect 10999 550 11041 560
rect 13249 599 13373 608
rect 13249 559 13250 599
rect 13372 559 13373 599
rect 13249 550 13373 559
rect 15572 574 15640 610
rect 10880 474 10912 490
rect 15572 542 15590 574
rect 15622 542 15640 574
rect 15572 506 15640 542
rect 15572 474 15590 506
rect 15622 474 15640 506
rect 360 438 428 474
rect 15572 438 15640 474
rect 360 420 15640 438
rect 360 388 402 420
rect 434 388 470 420
rect 502 388 538 420
rect 570 388 606 420
rect 638 388 674 420
rect 706 388 742 420
rect 774 388 810 420
rect 842 388 878 420
rect 910 388 946 420
rect 978 388 1014 420
rect 1046 388 1082 420
rect 1114 388 1150 420
rect 1182 388 1218 420
rect 1250 388 1286 420
rect 1318 388 1354 420
rect 1386 388 1422 420
rect 1454 388 1490 420
rect 1522 388 1558 420
rect 1590 388 1626 420
rect 1658 388 1694 420
rect 1726 388 1762 420
rect 1794 388 1830 420
rect 1862 388 1898 420
rect 1930 388 1966 420
rect 1998 388 2034 420
rect 2066 388 2102 420
rect 2134 388 2170 420
rect 2202 388 2238 420
rect 2270 388 2306 420
rect 2338 388 2374 420
rect 2406 388 2442 420
rect 2474 388 2510 420
rect 2542 388 2578 420
rect 2610 388 2646 420
rect 2678 388 2714 420
rect 2746 388 2782 420
rect 2814 388 2850 420
rect 2882 388 2918 420
rect 2950 388 2986 420
rect 3018 388 3054 420
rect 3086 388 3122 420
rect 3154 388 3190 420
rect 3222 388 3258 420
rect 3290 388 3326 420
rect 3358 388 3394 420
rect 3426 388 3462 420
rect 3494 388 3530 420
rect 3562 388 3598 420
rect 3630 388 3666 420
rect 3698 388 3734 420
rect 3766 388 3802 420
rect 3834 388 3870 420
rect 3902 388 3938 420
rect 3970 388 4006 420
rect 4038 388 4074 420
rect 4106 388 4142 420
rect 4174 388 4210 420
rect 4242 388 4278 420
rect 4310 388 4346 420
rect 4378 388 4414 420
rect 4446 388 4482 420
rect 4514 388 4550 420
rect 4582 388 4618 420
rect 4650 388 4686 420
rect 4718 388 4754 420
rect 4786 388 4822 420
rect 4854 388 4890 420
rect 4922 388 4958 420
rect 4990 414 5026 420
rect 5000 388 5026 414
rect 5058 388 5094 420
rect 5126 388 5162 420
rect 5194 388 5230 420
rect 5262 388 5298 420
rect 5330 388 5366 420
rect 5398 388 5434 420
rect 5466 388 5502 420
rect 5534 414 5570 420
rect 5602 414 5638 420
rect 5534 388 5564 414
rect 5604 388 5638 414
rect 5670 388 5706 420
rect 5738 388 5774 420
rect 5806 388 5842 420
rect 5874 388 5910 420
rect 5942 388 5978 420
rect 6010 388 6046 420
rect 6078 388 6114 420
rect 6146 414 6182 420
rect 6146 388 6168 414
rect 6214 388 6250 420
rect 6282 388 6318 420
rect 6350 388 6386 420
rect 6418 388 6454 420
rect 6486 388 6522 420
rect 6554 388 6590 420
rect 6622 388 6658 420
rect 6690 388 6726 420
rect 6758 414 6794 420
rect 6758 388 6772 414
rect 6826 388 6862 420
rect 6894 388 6930 420
rect 6962 388 6998 420
rect 7030 388 7066 420
rect 7098 388 7134 420
rect 7166 388 7202 420
rect 7234 388 7270 420
rect 7302 388 7338 420
rect 7370 414 7406 420
rect 7370 388 7376 414
rect 7438 388 7474 420
rect 7506 388 7542 420
rect 7574 388 7610 420
rect 7642 388 7678 420
rect 7710 388 7746 420
rect 7778 388 7814 420
rect 7846 388 7882 420
rect 7914 388 7950 420
rect 7982 414 8018 420
rect 8050 388 8086 420
rect 8118 388 8154 420
rect 8186 388 8222 420
rect 8254 388 8290 420
rect 8322 388 8358 420
rect 8390 388 8426 420
rect 8458 388 8494 420
rect 8526 388 8562 420
rect 8594 414 8630 420
rect 8624 388 8630 414
rect 8662 388 8698 420
rect 8730 388 8766 420
rect 8798 388 8834 420
rect 8866 388 8902 420
rect 8934 388 8970 420
rect 9002 388 9038 420
rect 9070 388 9106 420
rect 9138 388 9174 420
rect 9206 414 9242 420
rect 9228 388 9242 414
rect 9274 388 9310 420
rect 9342 388 9378 420
rect 9410 388 9446 420
rect 9478 388 9514 420
rect 9546 388 9582 420
rect 9614 388 9650 420
rect 9682 388 9718 420
rect 9750 388 9786 420
rect 9818 414 9854 420
rect 9832 388 9854 414
rect 9886 388 9922 420
rect 9954 388 9990 420
rect 10022 388 10058 420
rect 10090 388 10126 420
rect 10158 388 10194 420
rect 10226 388 10262 420
rect 10294 388 10330 420
rect 10362 414 10398 420
rect 10430 414 10466 420
rect 10362 388 10396 414
rect 10436 388 10466 414
rect 10498 388 10534 420
rect 10566 388 10602 420
rect 10634 388 10670 420
rect 10702 388 10738 420
rect 10770 388 10806 420
rect 10838 388 10874 420
rect 10906 388 10942 420
rect 10974 414 11010 420
rect 10974 388 11000 414
rect 11042 388 11078 420
rect 11110 388 11146 420
rect 11178 388 11214 420
rect 11246 388 11282 420
rect 11314 388 11350 420
rect 11382 388 11418 420
rect 11450 388 11486 420
rect 11518 388 11554 420
rect 11586 388 11622 420
rect 11654 388 11690 420
rect 11722 388 11758 420
rect 11790 388 11826 420
rect 11858 388 11894 420
rect 11926 388 11962 420
rect 11994 388 12030 420
rect 12062 388 12098 420
rect 12130 388 12166 420
rect 12198 388 12234 420
rect 12266 388 12302 420
rect 12334 388 12370 420
rect 12402 388 12438 420
rect 12470 388 12506 420
rect 12538 388 12574 420
rect 12606 388 12642 420
rect 12674 388 12710 420
rect 12742 388 12778 420
rect 12810 388 12846 420
rect 12878 388 12914 420
rect 12946 388 12982 420
rect 13014 388 13050 420
rect 13082 388 13118 420
rect 13150 388 13186 420
rect 13218 414 13254 420
rect 13286 414 13322 420
rect 13354 414 13390 420
rect 13218 388 13250 414
rect 13372 388 13390 414
rect 13422 388 13458 420
rect 13490 388 13526 420
rect 13558 388 13594 420
rect 13626 388 13662 420
rect 13694 388 13730 420
rect 13762 388 13798 420
rect 13830 388 13866 420
rect 13898 388 13934 420
rect 13966 388 14002 420
rect 14034 388 14070 420
rect 14102 388 14138 420
rect 14170 388 14206 420
rect 14238 388 14274 420
rect 14306 388 14342 420
rect 14374 388 14410 420
rect 14442 388 14478 420
rect 14510 388 14546 420
rect 14578 388 14614 420
rect 14646 388 14682 420
rect 14714 388 14750 420
rect 14782 388 14818 420
rect 14850 388 14886 420
rect 14918 388 14954 420
rect 14986 388 15022 420
rect 15054 388 15090 420
rect 15122 388 15158 420
rect 15190 388 15226 420
rect 15258 388 15294 420
rect 15326 388 15362 420
rect 15394 388 15430 420
rect 15462 388 15498 420
rect 15530 388 15566 420
rect 15598 388 15640 420
rect 360 374 4960 388
rect 5000 374 5564 388
rect 5604 374 6168 388
rect 6208 374 6772 388
rect 6812 374 7376 388
rect 7416 374 7980 388
rect 8020 374 8584 388
rect 8624 374 9188 388
rect 9228 374 9792 388
rect 9832 374 10396 388
rect 10436 374 11000 388
rect 11040 374 13250 388
rect 13372 374 15640 388
rect 360 370 15640 374
rect 15932 1620 15950 1652
rect 15982 1620 16000 1652
rect 15932 1584 16000 1620
rect 15932 1552 15950 1584
rect 15982 1552 16000 1584
rect 15932 1516 16000 1552
rect 15932 1484 15950 1516
rect 15982 1484 16000 1516
rect 15932 1448 16000 1484
rect 15932 1416 15950 1448
rect 15982 1416 16000 1448
rect 15932 1380 16000 1416
rect 15932 1348 15950 1380
rect 15982 1348 16000 1380
rect 15932 1312 16000 1348
rect 15932 1280 15950 1312
rect 15982 1280 16000 1312
rect 15932 1244 16000 1280
rect 15932 1212 15950 1244
rect 15982 1212 16000 1244
rect 15932 1176 16000 1212
rect 15932 1144 15950 1176
rect 15982 1144 16000 1176
rect 15932 1108 16000 1144
rect 15932 1076 15950 1108
rect 15982 1076 16000 1108
rect 15932 1040 16000 1076
rect 15932 1008 15950 1040
rect 15982 1008 16000 1040
rect 15932 972 16000 1008
rect 15932 940 15950 972
rect 15982 940 16000 972
rect 15932 904 16000 940
rect 15932 872 15950 904
rect 15982 872 16000 904
rect 15932 836 16000 872
rect 15932 804 15950 836
rect 15982 804 16000 836
rect 15932 768 16000 804
rect 15932 736 15950 768
rect 15982 736 16000 768
rect 15932 700 16000 736
rect 15932 668 15950 700
rect 15982 668 16000 700
rect 15932 632 16000 668
rect 15932 600 15950 632
rect 15982 600 16000 632
rect 15932 564 16000 600
rect 15932 532 15950 564
rect 15982 532 16000 564
rect 15932 496 16000 532
rect 15932 464 15950 496
rect 15982 464 16000 496
rect 15932 428 16000 464
rect 15932 396 15950 428
rect 15982 396 16000 428
rect 4959 360 5001 370
rect 5563 360 5605 370
rect 6167 360 6209 370
rect 6771 360 6813 370
rect 7375 360 7417 370
rect 7979 360 8021 370
rect 8583 360 8625 370
rect 9187 360 9229 370
rect 9791 360 9833 370
rect 10395 360 10437 370
rect 10999 360 11041 370
rect 13249 365 13373 370
rect 15932 360 16000 396
rect 0 328 18 360
rect 50 328 68 360
rect 0 292 68 328
rect 0 260 18 292
rect 50 260 68 292
rect 0 224 68 260
rect 0 192 18 224
rect 50 192 68 224
rect 0 156 68 192
rect 0 124 18 156
rect 50 124 68 156
rect 0 68 68 124
rect 15932 328 15950 360
rect 15982 328 16000 360
rect 15932 292 16000 328
rect 15932 260 15950 292
rect 15982 260 16000 292
rect 15932 224 16000 260
rect 15932 192 15950 224
rect 15982 192 16000 224
rect 15932 156 16000 192
rect 15932 124 15950 156
rect 15982 124 16000 156
rect 15932 68 16000 124
rect 0 50 16000 68
rect 0 18 28 50
rect 60 18 96 50
rect 128 18 164 50
rect 196 18 232 50
rect 264 18 300 50
rect 332 18 368 50
rect 400 18 436 50
rect 468 18 504 50
rect 536 18 572 50
rect 604 18 640 50
rect 672 18 708 50
rect 740 18 776 50
rect 808 18 844 50
rect 876 18 912 50
rect 944 18 980 50
rect 1012 18 1048 50
rect 1080 18 1116 50
rect 1148 18 1184 50
rect 1216 18 1252 50
rect 1284 18 1320 50
rect 1352 18 1388 50
rect 1420 18 1456 50
rect 1488 18 1524 50
rect 1556 18 1592 50
rect 1624 18 1660 50
rect 1692 18 1728 50
rect 1760 18 1796 50
rect 1828 18 1864 50
rect 1896 18 1932 50
rect 1964 18 2000 50
rect 2032 18 2068 50
rect 2100 18 2136 50
rect 2168 18 2204 50
rect 2236 18 2272 50
rect 2304 18 2340 50
rect 2372 18 2408 50
rect 2440 18 2476 50
rect 2508 18 2544 50
rect 2576 18 2612 50
rect 2644 18 2680 50
rect 2712 18 2748 50
rect 2780 18 2816 50
rect 2848 18 2884 50
rect 2916 18 2952 50
rect 2984 18 3020 50
rect 3052 18 3088 50
rect 3120 18 3156 50
rect 3188 18 3224 50
rect 3256 18 3292 50
rect 3324 18 3360 50
rect 3392 18 3428 50
rect 3460 18 3496 50
rect 3528 18 3564 50
rect 3596 18 3632 50
rect 3664 18 3700 50
rect 3732 18 3768 50
rect 3800 18 3836 50
rect 3868 18 3904 50
rect 3936 18 3972 50
rect 4004 18 4040 50
rect 4072 18 4108 50
rect 4140 18 4176 50
rect 4208 18 4244 50
rect 4276 18 4312 50
rect 4344 18 4380 50
rect 4412 18 4448 50
rect 4480 18 4516 50
rect 4548 18 4584 50
rect 4616 18 4652 50
rect 4684 18 4720 50
rect 4752 18 4788 50
rect 4820 18 4856 50
rect 4888 18 4924 50
rect 4956 18 4992 50
rect 5024 18 5060 50
rect 5092 18 5128 50
rect 5160 18 5196 50
rect 5228 18 5264 50
rect 5296 18 5332 50
rect 5364 18 5400 50
rect 5432 18 5468 50
rect 5500 18 5536 50
rect 5568 18 5604 50
rect 5636 18 5672 50
rect 5704 18 5740 50
rect 5772 18 5808 50
rect 5840 18 5876 50
rect 5908 18 5944 50
rect 5976 18 6012 50
rect 6044 18 6080 50
rect 6112 18 6148 50
rect 6180 18 6216 50
rect 6248 18 6284 50
rect 6316 18 6352 50
rect 6384 18 6420 50
rect 6452 18 6488 50
rect 6520 18 6556 50
rect 6588 18 6624 50
rect 6656 18 6692 50
rect 6724 18 6760 50
rect 6792 18 6828 50
rect 6860 18 6896 50
rect 6928 18 6964 50
rect 6996 18 7032 50
rect 7064 18 7100 50
rect 7132 18 7168 50
rect 7200 18 7236 50
rect 7268 18 7304 50
rect 7336 18 7372 50
rect 7404 18 7440 50
rect 7472 18 7508 50
rect 7540 18 7576 50
rect 7608 18 7644 50
rect 7676 18 7712 50
rect 7744 18 7780 50
rect 7812 18 7848 50
rect 7880 18 7916 50
rect 7948 18 7984 50
rect 8016 18 8052 50
rect 8084 18 8120 50
rect 8152 18 8188 50
rect 8220 18 8256 50
rect 8288 18 8324 50
rect 8356 18 8392 50
rect 8424 18 8460 50
rect 8492 18 8528 50
rect 8560 18 8596 50
rect 8628 18 8664 50
rect 8696 18 8732 50
rect 8764 18 8800 50
rect 8832 18 8868 50
rect 8900 18 8936 50
rect 8968 18 9004 50
rect 9036 18 9072 50
rect 9104 18 9140 50
rect 9172 18 9208 50
rect 9240 18 9276 50
rect 9308 18 9344 50
rect 9376 18 9412 50
rect 9444 18 9480 50
rect 9512 18 9548 50
rect 9580 18 9616 50
rect 9648 18 9684 50
rect 9716 18 9752 50
rect 9784 18 9820 50
rect 9852 18 9888 50
rect 9920 18 9956 50
rect 9988 18 10024 50
rect 10056 18 10092 50
rect 10124 18 10160 50
rect 10192 18 10228 50
rect 10260 18 10296 50
rect 10328 18 10364 50
rect 10396 18 10432 50
rect 10464 18 10500 50
rect 10532 18 10568 50
rect 10600 18 10636 50
rect 10668 18 10704 50
rect 10736 18 10772 50
rect 10804 18 10840 50
rect 10872 18 10908 50
rect 10940 18 10976 50
rect 11008 18 11044 50
rect 11076 18 11112 50
rect 11144 18 11180 50
rect 11212 18 11248 50
rect 11280 18 11316 50
rect 11348 18 11384 50
rect 11416 18 11452 50
rect 11484 18 11520 50
rect 11552 18 11588 50
rect 11620 18 11656 50
rect 11688 18 11724 50
rect 11756 18 11792 50
rect 11824 18 11860 50
rect 11892 18 11928 50
rect 11960 18 11996 50
rect 12028 18 12064 50
rect 12096 18 12132 50
rect 12164 18 12200 50
rect 12232 18 12268 50
rect 12300 18 12336 50
rect 12368 18 12404 50
rect 12436 18 12472 50
rect 12504 18 12540 50
rect 12572 18 12608 50
rect 12640 18 12676 50
rect 12708 18 12744 50
rect 12776 18 12812 50
rect 12844 18 12880 50
rect 12912 18 12948 50
rect 12980 18 13016 50
rect 13048 18 13084 50
rect 13116 18 13152 50
rect 13184 18 13220 50
rect 13252 18 13288 50
rect 13320 18 13356 50
rect 13388 18 13424 50
rect 13456 18 13492 50
rect 13524 18 13560 50
rect 13592 18 13628 50
rect 13660 18 13696 50
rect 13728 18 13764 50
rect 13796 18 13832 50
rect 13864 18 13900 50
rect 13932 18 13968 50
rect 14000 18 14036 50
rect 14068 18 14104 50
rect 14136 18 14172 50
rect 14204 18 14240 50
rect 14272 18 14308 50
rect 14340 18 14376 50
rect 14408 18 14444 50
rect 14476 18 14512 50
rect 14544 18 14580 50
rect 14612 18 14648 50
rect 14680 18 14716 50
rect 14748 18 14784 50
rect 14816 18 14852 50
rect 14884 18 14920 50
rect 14952 18 14988 50
rect 15020 18 15056 50
rect 15088 18 15124 50
rect 15156 18 15192 50
rect 15224 18 15260 50
rect 15292 18 15328 50
rect 15360 18 15396 50
rect 15428 18 15464 50
rect 15496 18 15532 50
rect 15564 18 15600 50
rect 15632 18 15668 50
rect 15700 18 15736 50
rect 15768 18 15804 50
rect 15836 18 15872 50
rect 15904 18 15940 50
rect 15972 18 16000 50
rect 0 2 16000 18
rect 2 0 16000 2
<< via1 >>
rect 4960 1580 4990 1606
rect 4990 1580 5000 1606
rect 5564 1580 5570 1606
rect 5570 1580 5602 1606
rect 5602 1580 5604 1606
rect 6168 1580 6182 1606
rect 6182 1580 6208 1606
rect 6772 1580 6794 1606
rect 6794 1580 6812 1606
rect 7376 1580 7406 1606
rect 7406 1580 7416 1606
rect 7980 1580 7982 1606
rect 7982 1580 8018 1606
rect 8018 1580 8020 1606
rect 8584 1580 8594 1606
rect 8594 1580 8624 1606
rect 9188 1580 9206 1606
rect 9206 1580 9228 1606
rect 9792 1580 9818 1606
rect 9818 1580 9832 1606
rect 10396 1580 10398 1606
rect 10398 1580 10430 1606
rect 10430 1580 10436 1606
rect 11000 1580 11010 1606
rect 11010 1580 11040 1606
rect 4960 1566 5000 1580
rect 5564 1566 5604 1580
rect 6168 1566 6208 1580
rect 6772 1566 6812 1580
rect 7376 1566 7416 1580
rect 7980 1566 8020 1580
rect 8584 1566 8624 1580
rect 9188 1566 9228 1580
rect 9792 1566 9832 1580
rect 10396 1566 10436 1580
rect 11000 1566 11040 1580
rect 4960 1414 5000 1420
rect 4960 1382 4964 1414
rect 4964 1382 4996 1414
rect 4996 1382 5000 1414
rect 4960 1346 5000 1382
rect 4960 1314 4964 1346
rect 4964 1314 4996 1346
rect 4996 1314 5000 1346
rect 4960 1278 5000 1314
rect 4960 1246 4964 1278
rect 4964 1246 4996 1278
rect 4996 1246 5000 1278
rect 4960 1210 5000 1246
rect 4960 1178 4964 1210
rect 4964 1178 4996 1210
rect 4996 1178 5000 1210
rect 4960 1142 5000 1178
rect 4960 1110 4964 1142
rect 4964 1110 4996 1142
rect 4996 1110 5000 1142
rect 4960 1074 5000 1110
rect 4960 1042 4964 1074
rect 4964 1042 4996 1074
rect 4996 1042 5000 1074
rect 4960 1006 5000 1042
rect 4960 974 4964 1006
rect 4964 974 4996 1006
rect 4996 974 5000 1006
rect 4960 938 5000 974
rect 4960 906 4964 938
rect 4964 906 4996 938
rect 4996 906 5000 938
rect 4960 870 5000 906
rect 4960 838 4964 870
rect 4964 838 4996 870
rect 4996 838 5000 870
rect 4960 802 5000 838
rect 4960 770 4964 802
rect 4964 770 4996 802
rect 4996 770 5000 802
rect 4960 734 5000 770
rect 4960 702 4964 734
rect 4964 702 4996 734
rect 4996 702 5000 734
rect 4960 666 5000 702
rect 4960 634 4964 666
rect 4964 634 4996 666
rect 4996 634 5000 666
rect 4960 598 5000 634
rect 4960 566 4964 598
rect 4964 566 4996 598
rect 4996 566 5000 598
rect 4960 560 5000 566
rect 5221 1414 5343 1420
rect 5221 1382 5266 1414
rect 5266 1382 5298 1414
rect 5298 1382 5343 1414
rect 5221 1346 5343 1382
rect 5221 1314 5266 1346
rect 5266 1314 5298 1346
rect 5298 1314 5343 1346
rect 5221 1278 5343 1314
rect 5221 1246 5266 1278
rect 5266 1246 5298 1278
rect 5298 1246 5343 1278
rect 5221 1210 5343 1246
rect 5221 1178 5266 1210
rect 5266 1178 5298 1210
rect 5298 1178 5343 1210
rect 5221 1142 5343 1178
rect 5221 1110 5266 1142
rect 5266 1110 5298 1142
rect 5298 1110 5343 1142
rect 5221 1074 5343 1110
rect 5221 1042 5266 1074
rect 5266 1042 5298 1074
rect 5298 1042 5343 1074
rect 5221 1006 5343 1042
rect 5221 974 5266 1006
rect 5266 974 5298 1006
rect 5298 974 5343 1006
rect 5221 938 5343 974
rect 5221 906 5266 938
rect 5266 906 5298 938
rect 5298 906 5343 938
rect 5221 870 5343 906
rect 5221 838 5266 870
rect 5266 838 5298 870
rect 5298 838 5343 870
rect 5221 802 5343 838
rect 5221 770 5266 802
rect 5266 770 5298 802
rect 5298 770 5343 802
rect 5221 734 5343 770
rect 5221 702 5266 734
rect 5266 702 5298 734
rect 5298 702 5343 734
rect 5221 666 5343 702
rect 5221 634 5266 666
rect 5266 634 5298 666
rect 5298 634 5343 666
rect 5221 598 5343 634
rect 5221 566 5266 598
rect 5266 566 5298 598
rect 5298 566 5343 598
rect 5221 560 5343 566
rect 5564 1414 5604 1420
rect 5564 1382 5568 1414
rect 5568 1382 5600 1414
rect 5600 1382 5604 1414
rect 5564 1346 5604 1382
rect 5564 1314 5568 1346
rect 5568 1314 5600 1346
rect 5600 1314 5604 1346
rect 5564 1278 5604 1314
rect 5564 1246 5568 1278
rect 5568 1246 5600 1278
rect 5600 1246 5604 1278
rect 5564 1210 5604 1246
rect 5564 1178 5568 1210
rect 5568 1178 5600 1210
rect 5600 1178 5604 1210
rect 5564 1142 5604 1178
rect 5564 1110 5568 1142
rect 5568 1110 5600 1142
rect 5600 1110 5604 1142
rect 5564 1074 5604 1110
rect 5564 1042 5568 1074
rect 5568 1042 5600 1074
rect 5600 1042 5604 1074
rect 5564 1006 5604 1042
rect 5564 974 5568 1006
rect 5568 974 5600 1006
rect 5600 974 5604 1006
rect 5564 938 5604 974
rect 5564 906 5568 938
rect 5568 906 5600 938
rect 5600 906 5604 938
rect 5564 870 5604 906
rect 5564 838 5568 870
rect 5568 838 5600 870
rect 5600 838 5604 870
rect 5564 802 5604 838
rect 5564 770 5568 802
rect 5568 770 5600 802
rect 5600 770 5604 802
rect 5564 734 5604 770
rect 5564 702 5568 734
rect 5568 702 5600 734
rect 5600 702 5604 734
rect 5564 666 5604 702
rect 5564 634 5568 666
rect 5568 634 5600 666
rect 5600 634 5604 666
rect 5564 598 5604 634
rect 5564 566 5568 598
rect 5568 566 5600 598
rect 5600 566 5604 598
rect 5564 560 5604 566
rect 5825 1414 5947 1420
rect 5825 1382 5870 1414
rect 5870 1382 5902 1414
rect 5902 1382 5947 1414
rect 5825 1346 5947 1382
rect 5825 1314 5870 1346
rect 5870 1314 5902 1346
rect 5902 1314 5947 1346
rect 5825 1278 5947 1314
rect 5825 1246 5870 1278
rect 5870 1246 5902 1278
rect 5902 1246 5947 1278
rect 5825 1210 5947 1246
rect 5825 1178 5870 1210
rect 5870 1178 5902 1210
rect 5902 1178 5947 1210
rect 5825 1142 5947 1178
rect 5825 1110 5870 1142
rect 5870 1110 5902 1142
rect 5902 1110 5947 1142
rect 5825 1074 5947 1110
rect 5825 1042 5870 1074
rect 5870 1042 5902 1074
rect 5902 1042 5947 1074
rect 5825 1006 5947 1042
rect 5825 974 5870 1006
rect 5870 974 5902 1006
rect 5902 974 5947 1006
rect 5825 938 5947 974
rect 5825 906 5870 938
rect 5870 906 5902 938
rect 5902 906 5947 938
rect 5825 870 5947 906
rect 5825 838 5870 870
rect 5870 838 5902 870
rect 5902 838 5947 870
rect 5825 802 5947 838
rect 5825 770 5870 802
rect 5870 770 5902 802
rect 5902 770 5947 802
rect 5825 734 5947 770
rect 5825 702 5870 734
rect 5870 702 5902 734
rect 5902 702 5947 734
rect 5825 666 5947 702
rect 5825 634 5870 666
rect 5870 634 5902 666
rect 5902 634 5947 666
rect 5825 598 5947 634
rect 5825 566 5870 598
rect 5870 566 5902 598
rect 5902 566 5947 598
rect 5825 560 5947 566
rect 6168 1414 6208 1420
rect 6168 1382 6172 1414
rect 6172 1382 6204 1414
rect 6204 1382 6208 1414
rect 6168 1346 6208 1382
rect 6168 1314 6172 1346
rect 6172 1314 6204 1346
rect 6204 1314 6208 1346
rect 6168 1278 6208 1314
rect 6168 1246 6172 1278
rect 6172 1246 6204 1278
rect 6204 1246 6208 1278
rect 6168 1210 6208 1246
rect 6168 1178 6172 1210
rect 6172 1178 6204 1210
rect 6204 1178 6208 1210
rect 6168 1142 6208 1178
rect 6168 1110 6172 1142
rect 6172 1110 6204 1142
rect 6204 1110 6208 1142
rect 6168 1074 6208 1110
rect 6168 1042 6172 1074
rect 6172 1042 6204 1074
rect 6204 1042 6208 1074
rect 6168 1006 6208 1042
rect 6168 974 6172 1006
rect 6172 974 6204 1006
rect 6204 974 6208 1006
rect 6168 938 6208 974
rect 6168 906 6172 938
rect 6172 906 6204 938
rect 6204 906 6208 938
rect 6168 870 6208 906
rect 6168 838 6172 870
rect 6172 838 6204 870
rect 6204 838 6208 870
rect 6168 802 6208 838
rect 6168 770 6172 802
rect 6172 770 6204 802
rect 6204 770 6208 802
rect 6168 734 6208 770
rect 6168 702 6172 734
rect 6172 702 6204 734
rect 6204 702 6208 734
rect 6168 666 6208 702
rect 6168 634 6172 666
rect 6172 634 6204 666
rect 6204 634 6208 666
rect 6168 598 6208 634
rect 6168 566 6172 598
rect 6172 566 6204 598
rect 6204 566 6208 598
rect 6168 560 6208 566
rect 6429 1414 6551 1420
rect 6429 1382 6474 1414
rect 6474 1382 6506 1414
rect 6506 1382 6551 1414
rect 6429 1346 6551 1382
rect 6429 1314 6474 1346
rect 6474 1314 6506 1346
rect 6506 1314 6551 1346
rect 6429 1278 6551 1314
rect 6429 1246 6474 1278
rect 6474 1246 6506 1278
rect 6506 1246 6551 1278
rect 6429 1210 6551 1246
rect 6429 1178 6474 1210
rect 6474 1178 6506 1210
rect 6506 1178 6551 1210
rect 6429 1142 6551 1178
rect 6429 1110 6474 1142
rect 6474 1110 6506 1142
rect 6506 1110 6551 1142
rect 6429 1074 6551 1110
rect 6429 1042 6474 1074
rect 6474 1042 6506 1074
rect 6506 1042 6551 1074
rect 6429 1006 6551 1042
rect 6429 974 6474 1006
rect 6474 974 6506 1006
rect 6506 974 6551 1006
rect 6429 938 6551 974
rect 6429 906 6474 938
rect 6474 906 6506 938
rect 6506 906 6551 938
rect 6429 870 6551 906
rect 6429 838 6474 870
rect 6474 838 6506 870
rect 6506 838 6551 870
rect 6429 802 6551 838
rect 6429 770 6474 802
rect 6474 770 6506 802
rect 6506 770 6551 802
rect 6429 734 6551 770
rect 6429 702 6474 734
rect 6474 702 6506 734
rect 6506 702 6551 734
rect 6429 666 6551 702
rect 6429 634 6474 666
rect 6474 634 6506 666
rect 6506 634 6551 666
rect 6429 598 6551 634
rect 6429 566 6474 598
rect 6474 566 6506 598
rect 6506 566 6551 598
rect 6429 560 6551 566
rect 6772 1414 6812 1420
rect 6772 1382 6776 1414
rect 6776 1382 6808 1414
rect 6808 1382 6812 1414
rect 6772 1346 6812 1382
rect 6772 1314 6776 1346
rect 6776 1314 6808 1346
rect 6808 1314 6812 1346
rect 6772 1278 6812 1314
rect 6772 1246 6776 1278
rect 6776 1246 6808 1278
rect 6808 1246 6812 1278
rect 6772 1210 6812 1246
rect 6772 1178 6776 1210
rect 6776 1178 6808 1210
rect 6808 1178 6812 1210
rect 6772 1142 6812 1178
rect 6772 1110 6776 1142
rect 6776 1110 6808 1142
rect 6808 1110 6812 1142
rect 6772 1074 6812 1110
rect 6772 1042 6776 1074
rect 6776 1042 6808 1074
rect 6808 1042 6812 1074
rect 6772 1006 6812 1042
rect 6772 974 6776 1006
rect 6776 974 6808 1006
rect 6808 974 6812 1006
rect 6772 938 6812 974
rect 6772 906 6776 938
rect 6776 906 6808 938
rect 6808 906 6812 938
rect 6772 870 6812 906
rect 6772 838 6776 870
rect 6776 838 6808 870
rect 6808 838 6812 870
rect 6772 802 6812 838
rect 6772 770 6776 802
rect 6776 770 6808 802
rect 6808 770 6812 802
rect 6772 734 6812 770
rect 6772 702 6776 734
rect 6776 702 6808 734
rect 6808 702 6812 734
rect 6772 666 6812 702
rect 6772 634 6776 666
rect 6776 634 6808 666
rect 6808 634 6812 666
rect 6772 598 6812 634
rect 6772 566 6776 598
rect 6776 566 6808 598
rect 6808 566 6812 598
rect 6772 560 6812 566
rect 7033 1414 7155 1420
rect 7033 1382 7078 1414
rect 7078 1382 7110 1414
rect 7110 1382 7155 1414
rect 7033 1346 7155 1382
rect 7033 1314 7078 1346
rect 7078 1314 7110 1346
rect 7110 1314 7155 1346
rect 7033 1278 7155 1314
rect 7033 1246 7078 1278
rect 7078 1246 7110 1278
rect 7110 1246 7155 1278
rect 7033 1210 7155 1246
rect 7033 1178 7078 1210
rect 7078 1178 7110 1210
rect 7110 1178 7155 1210
rect 7033 1142 7155 1178
rect 7033 1110 7078 1142
rect 7078 1110 7110 1142
rect 7110 1110 7155 1142
rect 7033 1074 7155 1110
rect 7033 1042 7078 1074
rect 7078 1042 7110 1074
rect 7110 1042 7155 1074
rect 7033 1006 7155 1042
rect 7033 974 7078 1006
rect 7078 974 7110 1006
rect 7110 974 7155 1006
rect 7033 938 7155 974
rect 7033 906 7078 938
rect 7078 906 7110 938
rect 7110 906 7155 938
rect 7033 870 7155 906
rect 7033 838 7078 870
rect 7078 838 7110 870
rect 7110 838 7155 870
rect 7033 802 7155 838
rect 7033 770 7078 802
rect 7078 770 7110 802
rect 7110 770 7155 802
rect 7033 734 7155 770
rect 7033 702 7078 734
rect 7078 702 7110 734
rect 7110 702 7155 734
rect 7033 666 7155 702
rect 7033 634 7078 666
rect 7078 634 7110 666
rect 7110 634 7155 666
rect 7033 598 7155 634
rect 7033 566 7078 598
rect 7078 566 7110 598
rect 7110 566 7155 598
rect 7033 560 7155 566
rect 7376 1414 7416 1420
rect 7376 1382 7380 1414
rect 7380 1382 7412 1414
rect 7412 1382 7416 1414
rect 7376 1346 7416 1382
rect 7376 1314 7380 1346
rect 7380 1314 7412 1346
rect 7412 1314 7416 1346
rect 7376 1278 7416 1314
rect 7376 1246 7380 1278
rect 7380 1246 7412 1278
rect 7412 1246 7416 1278
rect 7376 1210 7416 1246
rect 7376 1178 7380 1210
rect 7380 1178 7412 1210
rect 7412 1178 7416 1210
rect 7376 1142 7416 1178
rect 7376 1110 7380 1142
rect 7380 1110 7412 1142
rect 7412 1110 7416 1142
rect 7376 1074 7416 1110
rect 7376 1042 7380 1074
rect 7380 1042 7412 1074
rect 7412 1042 7416 1074
rect 7376 1006 7416 1042
rect 7376 974 7380 1006
rect 7380 974 7412 1006
rect 7412 974 7416 1006
rect 7376 938 7416 974
rect 7376 906 7380 938
rect 7380 906 7412 938
rect 7412 906 7416 938
rect 7376 870 7416 906
rect 7376 838 7380 870
rect 7380 838 7412 870
rect 7412 838 7416 870
rect 7376 802 7416 838
rect 7376 770 7380 802
rect 7380 770 7412 802
rect 7412 770 7416 802
rect 7376 734 7416 770
rect 7376 702 7380 734
rect 7380 702 7412 734
rect 7412 702 7416 734
rect 7376 666 7416 702
rect 7376 634 7380 666
rect 7380 634 7412 666
rect 7412 634 7416 666
rect 7376 598 7416 634
rect 7376 566 7380 598
rect 7380 566 7412 598
rect 7412 566 7416 598
rect 7376 560 7416 566
rect 7637 1414 7759 1420
rect 7637 1382 7682 1414
rect 7682 1382 7714 1414
rect 7714 1382 7759 1414
rect 7637 1346 7759 1382
rect 7637 1314 7682 1346
rect 7682 1314 7714 1346
rect 7714 1314 7759 1346
rect 7637 1278 7759 1314
rect 7637 1246 7682 1278
rect 7682 1246 7714 1278
rect 7714 1246 7759 1278
rect 7637 1210 7759 1246
rect 7637 1178 7682 1210
rect 7682 1178 7714 1210
rect 7714 1178 7759 1210
rect 7637 1142 7759 1178
rect 7637 1110 7682 1142
rect 7682 1110 7714 1142
rect 7714 1110 7759 1142
rect 7637 1074 7759 1110
rect 7637 1042 7682 1074
rect 7682 1042 7714 1074
rect 7714 1042 7759 1074
rect 7637 1006 7759 1042
rect 7637 974 7682 1006
rect 7682 974 7714 1006
rect 7714 974 7759 1006
rect 7637 938 7759 974
rect 7637 906 7682 938
rect 7682 906 7714 938
rect 7714 906 7759 938
rect 7637 870 7759 906
rect 7637 838 7682 870
rect 7682 838 7714 870
rect 7714 838 7759 870
rect 7637 802 7759 838
rect 7637 770 7682 802
rect 7682 770 7714 802
rect 7714 770 7759 802
rect 7637 734 7759 770
rect 7637 702 7682 734
rect 7682 702 7714 734
rect 7714 702 7759 734
rect 7637 666 7759 702
rect 7637 634 7682 666
rect 7682 634 7714 666
rect 7714 634 7759 666
rect 7637 598 7759 634
rect 7637 566 7682 598
rect 7682 566 7714 598
rect 7714 566 7759 598
rect 7637 560 7759 566
rect 7980 1414 8020 1420
rect 7980 1382 7984 1414
rect 7984 1382 8016 1414
rect 8016 1382 8020 1414
rect 7980 1346 8020 1382
rect 7980 1314 7984 1346
rect 7984 1314 8016 1346
rect 8016 1314 8020 1346
rect 7980 1278 8020 1314
rect 7980 1246 7984 1278
rect 7984 1246 8016 1278
rect 8016 1246 8020 1278
rect 7980 1210 8020 1246
rect 7980 1178 7984 1210
rect 7984 1178 8016 1210
rect 8016 1178 8020 1210
rect 7980 1142 8020 1178
rect 7980 1110 7984 1142
rect 7984 1110 8016 1142
rect 8016 1110 8020 1142
rect 7980 1074 8020 1110
rect 7980 1042 7984 1074
rect 7984 1042 8016 1074
rect 8016 1042 8020 1074
rect 7980 1006 8020 1042
rect 7980 974 7984 1006
rect 7984 974 8016 1006
rect 8016 974 8020 1006
rect 7980 938 8020 974
rect 7980 906 7984 938
rect 7984 906 8016 938
rect 8016 906 8020 938
rect 7980 870 8020 906
rect 7980 838 7984 870
rect 7984 838 8016 870
rect 8016 838 8020 870
rect 7980 802 8020 838
rect 7980 770 7984 802
rect 7984 770 8016 802
rect 8016 770 8020 802
rect 7980 734 8020 770
rect 7980 702 7984 734
rect 7984 702 8016 734
rect 8016 702 8020 734
rect 7980 666 8020 702
rect 7980 634 7984 666
rect 7984 634 8016 666
rect 8016 634 8020 666
rect 7980 598 8020 634
rect 7980 566 7984 598
rect 7984 566 8016 598
rect 8016 566 8020 598
rect 7980 560 8020 566
rect 8241 1414 8363 1420
rect 8241 1382 8286 1414
rect 8286 1382 8318 1414
rect 8318 1382 8363 1414
rect 8241 1346 8363 1382
rect 8241 1314 8286 1346
rect 8286 1314 8318 1346
rect 8318 1314 8363 1346
rect 8241 1278 8363 1314
rect 8241 1246 8286 1278
rect 8286 1246 8318 1278
rect 8318 1246 8363 1278
rect 8241 1210 8363 1246
rect 8241 1178 8286 1210
rect 8286 1178 8318 1210
rect 8318 1178 8363 1210
rect 8241 1142 8363 1178
rect 8241 1110 8286 1142
rect 8286 1110 8318 1142
rect 8318 1110 8363 1142
rect 8241 1074 8363 1110
rect 8241 1042 8286 1074
rect 8286 1042 8318 1074
rect 8318 1042 8363 1074
rect 8241 1006 8363 1042
rect 8241 974 8286 1006
rect 8286 974 8318 1006
rect 8318 974 8363 1006
rect 8241 938 8363 974
rect 8241 906 8286 938
rect 8286 906 8318 938
rect 8318 906 8363 938
rect 8241 870 8363 906
rect 8241 838 8286 870
rect 8286 838 8318 870
rect 8318 838 8363 870
rect 8241 802 8363 838
rect 8241 770 8286 802
rect 8286 770 8318 802
rect 8318 770 8363 802
rect 8241 734 8363 770
rect 8241 702 8286 734
rect 8286 702 8318 734
rect 8318 702 8363 734
rect 8241 666 8363 702
rect 8241 634 8286 666
rect 8286 634 8318 666
rect 8318 634 8363 666
rect 8241 598 8363 634
rect 8241 566 8286 598
rect 8286 566 8318 598
rect 8318 566 8363 598
rect 8241 560 8363 566
rect 8584 1414 8624 1420
rect 8584 1382 8588 1414
rect 8588 1382 8620 1414
rect 8620 1382 8624 1414
rect 8584 1346 8624 1382
rect 8584 1314 8588 1346
rect 8588 1314 8620 1346
rect 8620 1314 8624 1346
rect 8584 1278 8624 1314
rect 8584 1246 8588 1278
rect 8588 1246 8620 1278
rect 8620 1246 8624 1278
rect 8584 1210 8624 1246
rect 8584 1178 8588 1210
rect 8588 1178 8620 1210
rect 8620 1178 8624 1210
rect 8584 1142 8624 1178
rect 8584 1110 8588 1142
rect 8588 1110 8620 1142
rect 8620 1110 8624 1142
rect 8584 1074 8624 1110
rect 8584 1042 8588 1074
rect 8588 1042 8620 1074
rect 8620 1042 8624 1074
rect 8584 1006 8624 1042
rect 8584 974 8588 1006
rect 8588 974 8620 1006
rect 8620 974 8624 1006
rect 8584 938 8624 974
rect 8584 906 8588 938
rect 8588 906 8620 938
rect 8620 906 8624 938
rect 8584 870 8624 906
rect 8584 838 8588 870
rect 8588 838 8620 870
rect 8620 838 8624 870
rect 8584 802 8624 838
rect 8584 770 8588 802
rect 8588 770 8620 802
rect 8620 770 8624 802
rect 8584 734 8624 770
rect 8584 702 8588 734
rect 8588 702 8620 734
rect 8620 702 8624 734
rect 8584 666 8624 702
rect 8584 634 8588 666
rect 8588 634 8620 666
rect 8620 634 8624 666
rect 8584 598 8624 634
rect 8584 566 8588 598
rect 8588 566 8620 598
rect 8620 566 8624 598
rect 8584 560 8624 566
rect 8845 1414 8967 1420
rect 8845 1382 8890 1414
rect 8890 1382 8922 1414
rect 8922 1382 8967 1414
rect 8845 1346 8967 1382
rect 8845 1314 8890 1346
rect 8890 1314 8922 1346
rect 8922 1314 8967 1346
rect 8845 1278 8967 1314
rect 8845 1246 8890 1278
rect 8890 1246 8922 1278
rect 8922 1246 8967 1278
rect 8845 1210 8967 1246
rect 8845 1178 8890 1210
rect 8890 1178 8922 1210
rect 8922 1178 8967 1210
rect 8845 1142 8967 1178
rect 8845 1110 8890 1142
rect 8890 1110 8922 1142
rect 8922 1110 8967 1142
rect 8845 1074 8967 1110
rect 8845 1042 8890 1074
rect 8890 1042 8922 1074
rect 8922 1042 8967 1074
rect 8845 1006 8967 1042
rect 8845 974 8890 1006
rect 8890 974 8922 1006
rect 8922 974 8967 1006
rect 8845 938 8967 974
rect 8845 906 8890 938
rect 8890 906 8922 938
rect 8922 906 8967 938
rect 8845 870 8967 906
rect 8845 838 8890 870
rect 8890 838 8922 870
rect 8922 838 8967 870
rect 8845 802 8967 838
rect 8845 770 8890 802
rect 8890 770 8922 802
rect 8922 770 8967 802
rect 8845 734 8967 770
rect 8845 702 8890 734
rect 8890 702 8922 734
rect 8922 702 8967 734
rect 8845 666 8967 702
rect 8845 634 8890 666
rect 8890 634 8922 666
rect 8922 634 8967 666
rect 8845 598 8967 634
rect 8845 566 8890 598
rect 8890 566 8922 598
rect 8922 566 8967 598
rect 8845 560 8967 566
rect 9188 1414 9228 1420
rect 9188 1382 9192 1414
rect 9192 1382 9224 1414
rect 9224 1382 9228 1414
rect 9188 1346 9228 1382
rect 9188 1314 9192 1346
rect 9192 1314 9224 1346
rect 9224 1314 9228 1346
rect 9188 1278 9228 1314
rect 9188 1246 9192 1278
rect 9192 1246 9224 1278
rect 9224 1246 9228 1278
rect 9188 1210 9228 1246
rect 9188 1178 9192 1210
rect 9192 1178 9224 1210
rect 9224 1178 9228 1210
rect 9188 1142 9228 1178
rect 9188 1110 9192 1142
rect 9192 1110 9224 1142
rect 9224 1110 9228 1142
rect 9188 1074 9228 1110
rect 9188 1042 9192 1074
rect 9192 1042 9224 1074
rect 9224 1042 9228 1074
rect 9188 1006 9228 1042
rect 9188 974 9192 1006
rect 9192 974 9224 1006
rect 9224 974 9228 1006
rect 9188 938 9228 974
rect 9188 906 9192 938
rect 9192 906 9224 938
rect 9224 906 9228 938
rect 9188 870 9228 906
rect 9188 838 9192 870
rect 9192 838 9224 870
rect 9224 838 9228 870
rect 9188 802 9228 838
rect 9188 770 9192 802
rect 9192 770 9224 802
rect 9224 770 9228 802
rect 9188 734 9228 770
rect 9188 702 9192 734
rect 9192 702 9224 734
rect 9224 702 9228 734
rect 9188 666 9228 702
rect 9188 634 9192 666
rect 9192 634 9224 666
rect 9224 634 9228 666
rect 9188 598 9228 634
rect 9188 566 9192 598
rect 9192 566 9224 598
rect 9224 566 9228 598
rect 9188 560 9228 566
rect 9449 1414 9571 1420
rect 9449 1382 9494 1414
rect 9494 1382 9526 1414
rect 9526 1382 9571 1414
rect 9449 1346 9571 1382
rect 9449 1314 9494 1346
rect 9494 1314 9526 1346
rect 9526 1314 9571 1346
rect 9449 1278 9571 1314
rect 9449 1246 9494 1278
rect 9494 1246 9526 1278
rect 9526 1246 9571 1278
rect 9449 1210 9571 1246
rect 9449 1178 9494 1210
rect 9494 1178 9526 1210
rect 9526 1178 9571 1210
rect 9449 1142 9571 1178
rect 9449 1110 9494 1142
rect 9494 1110 9526 1142
rect 9526 1110 9571 1142
rect 9449 1074 9571 1110
rect 9449 1042 9494 1074
rect 9494 1042 9526 1074
rect 9526 1042 9571 1074
rect 9449 1006 9571 1042
rect 9449 974 9494 1006
rect 9494 974 9526 1006
rect 9526 974 9571 1006
rect 9449 938 9571 974
rect 9449 906 9494 938
rect 9494 906 9526 938
rect 9526 906 9571 938
rect 9449 870 9571 906
rect 9449 838 9494 870
rect 9494 838 9526 870
rect 9526 838 9571 870
rect 9449 802 9571 838
rect 9449 770 9494 802
rect 9494 770 9526 802
rect 9526 770 9571 802
rect 9449 734 9571 770
rect 9449 702 9494 734
rect 9494 702 9526 734
rect 9526 702 9571 734
rect 9449 666 9571 702
rect 9449 634 9494 666
rect 9494 634 9526 666
rect 9526 634 9571 666
rect 9449 598 9571 634
rect 9449 566 9494 598
rect 9494 566 9526 598
rect 9526 566 9571 598
rect 9449 560 9571 566
rect 9792 1414 9832 1420
rect 9792 1382 9796 1414
rect 9796 1382 9828 1414
rect 9828 1382 9832 1414
rect 9792 1346 9832 1382
rect 9792 1314 9796 1346
rect 9796 1314 9828 1346
rect 9828 1314 9832 1346
rect 9792 1278 9832 1314
rect 9792 1246 9796 1278
rect 9796 1246 9828 1278
rect 9828 1246 9832 1278
rect 9792 1210 9832 1246
rect 9792 1178 9796 1210
rect 9796 1178 9828 1210
rect 9828 1178 9832 1210
rect 9792 1142 9832 1178
rect 9792 1110 9796 1142
rect 9796 1110 9828 1142
rect 9828 1110 9832 1142
rect 9792 1074 9832 1110
rect 9792 1042 9796 1074
rect 9796 1042 9828 1074
rect 9828 1042 9832 1074
rect 9792 1006 9832 1042
rect 9792 974 9796 1006
rect 9796 974 9828 1006
rect 9828 974 9832 1006
rect 9792 938 9832 974
rect 9792 906 9796 938
rect 9796 906 9828 938
rect 9828 906 9832 938
rect 9792 870 9832 906
rect 9792 838 9796 870
rect 9796 838 9828 870
rect 9828 838 9832 870
rect 9792 802 9832 838
rect 9792 770 9796 802
rect 9796 770 9828 802
rect 9828 770 9832 802
rect 9792 734 9832 770
rect 9792 702 9796 734
rect 9796 702 9828 734
rect 9828 702 9832 734
rect 9792 666 9832 702
rect 9792 634 9796 666
rect 9796 634 9828 666
rect 9828 634 9832 666
rect 9792 598 9832 634
rect 9792 566 9796 598
rect 9796 566 9828 598
rect 9828 566 9832 598
rect 9792 560 9832 566
rect 10053 1414 10175 1420
rect 10053 1382 10098 1414
rect 10098 1382 10130 1414
rect 10130 1382 10175 1414
rect 10053 1346 10175 1382
rect 10053 1314 10098 1346
rect 10098 1314 10130 1346
rect 10130 1314 10175 1346
rect 10053 1278 10175 1314
rect 10053 1246 10098 1278
rect 10098 1246 10130 1278
rect 10130 1246 10175 1278
rect 10053 1210 10175 1246
rect 10053 1178 10098 1210
rect 10098 1178 10130 1210
rect 10130 1178 10175 1210
rect 10053 1142 10175 1178
rect 10053 1110 10098 1142
rect 10098 1110 10130 1142
rect 10130 1110 10175 1142
rect 10053 1074 10175 1110
rect 10053 1042 10098 1074
rect 10098 1042 10130 1074
rect 10130 1042 10175 1074
rect 10053 1006 10175 1042
rect 10053 974 10098 1006
rect 10098 974 10130 1006
rect 10130 974 10175 1006
rect 10053 938 10175 974
rect 10053 906 10098 938
rect 10098 906 10130 938
rect 10130 906 10175 938
rect 10053 870 10175 906
rect 10053 838 10098 870
rect 10098 838 10130 870
rect 10130 838 10175 870
rect 10053 802 10175 838
rect 10053 770 10098 802
rect 10098 770 10130 802
rect 10130 770 10175 802
rect 10053 734 10175 770
rect 10053 702 10098 734
rect 10098 702 10130 734
rect 10130 702 10175 734
rect 10053 666 10175 702
rect 10053 634 10098 666
rect 10098 634 10130 666
rect 10130 634 10175 666
rect 10053 598 10175 634
rect 10053 566 10098 598
rect 10098 566 10130 598
rect 10130 566 10175 598
rect 10053 560 10175 566
rect 10396 1414 10436 1420
rect 10396 1382 10400 1414
rect 10400 1382 10432 1414
rect 10432 1382 10436 1414
rect 10396 1346 10436 1382
rect 10396 1314 10400 1346
rect 10400 1314 10432 1346
rect 10432 1314 10436 1346
rect 10396 1278 10436 1314
rect 10396 1246 10400 1278
rect 10400 1246 10432 1278
rect 10432 1246 10436 1278
rect 10396 1210 10436 1246
rect 10396 1178 10400 1210
rect 10400 1178 10432 1210
rect 10432 1178 10436 1210
rect 10396 1142 10436 1178
rect 10396 1110 10400 1142
rect 10400 1110 10432 1142
rect 10432 1110 10436 1142
rect 10396 1074 10436 1110
rect 10396 1042 10400 1074
rect 10400 1042 10432 1074
rect 10432 1042 10436 1074
rect 10396 1006 10436 1042
rect 10396 974 10400 1006
rect 10400 974 10432 1006
rect 10432 974 10436 1006
rect 10396 938 10436 974
rect 10396 906 10400 938
rect 10400 906 10432 938
rect 10432 906 10436 938
rect 10396 870 10436 906
rect 10396 838 10400 870
rect 10400 838 10432 870
rect 10432 838 10436 870
rect 10396 802 10436 838
rect 10396 770 10400 802
rect 10400 770 10432 802
rect 10432 770 10436 802
rect 10396 734 10436 770
rect 10396 702 10400 734
rect 10400 702 10432 734
rect 10432 702 10436 734
rect 10396 666 10436 702
rect 10396 634 10400 666
rect 10400 634 10432 666
rect 10432 634 10436 666
rect 10396 598 10436 634
rect 10396 566 10400 598
rect 10400 566 10432 598
rect 10432 566 10436 598
rect 10396 560 10436 566
rect 10657 1414 10779 1420
rect 10657 1382 10702 1414
rect 10702 1382 10734 1414
rect 10734 1382 10779 1414
rect 10657 1346 10779 1382
rect 10657 1314 10702 1346
rect 10702 1314 10734 1346
rect 10734 1314 10779 1346
rect 10657 1278 10779 1314
rect 10657 1246 10702 1278
rect 10702 1246 10734 1278
rect 10734 1246 10779 1278
rect 10657 1210 10779 1246
rect 10657 1178 10702 1210
rect 10702 1178 10734 1210
rect 10734 1178 10779 1210
rect 10657 1142 10779 1178
rect 10657 1110 10702 1142
rect 10702 1110 10734 1142
rect 10734 1110 10779 1142
rect 10657 1074 10779 1110
rect 10657 1042 10702 1074
rect 10702 1042 10734 1074
rect 10734 1042 10779 1074
rect 10657 1006 10779 1042
rect 10657 974 10702 1006
rect 10702 974 10734 1006
rect 10734 974 10779 1006
rect 10657 938 10779 974
rect 10657 906 10702 938
rect 10702 906 10734 938
rect 10734 906 10779 938
rect 10657 870 10779 906
rect 10657 838 10702 870
rect 10702 838 10734 870
rect 10734 838 10779 870
rect 10657 802 10779 838
rect 10657 770 10702 802
rect 10702 770 10734 802
rect 10734 770 10779 802
rect 10657 734 10779 770
rect 10657 702 10702 734
rect 10702 702 10734 734
rect 10734 702 10779 734
rect 10657 666 10779 702
rect 10657 634 10702 666
rect 10702 634 10734 666
rect 10734 634 10779 666
rect 10657 598 10779 634
rect 10657 566 10702 598
rect 10702 566 10734 598
rect 10734 566 10779 598
rect 10657 560 10779 566
rect 11000 1414 11040 1420
rect 11000 1382 11004 1414
rect 11004 1382 11036 1414
rect 11036 1382 11040 1414
rect 11000 1346 11040 1382
rect 11000 1314 11004 1346
rect 11004 1314 11036 1346
rect 11036 1314 11040 1346
rect 11000 1278 11040 1314
rect 11000 1246 11004 1278
rect 11004 1246 11036 1278
rect 11036 1246 11040 1278
rect 11000 1210 11040 1246
rect 11000 1178 11004 1210
rect 11004 1178 11036 1210
rect 11036 1178 11040 1210
rect 11000 1142 11040 1178
rect 11000 1110 11004 1142
rect 11004 1110 11036 1142
rect 11036 1110 11040 1142
rect 11000 1074 11040 1110
rect 11000 1042 11004 1074
rect 11004 1042 11036 1074
rect 11036 1042 11040 1074
rect 11000 1006 11040 1042
rect 11000 974 11004 1006
rect 11004 974 11036 1006
rect 11036 974 11040 1006
rect 11000 938 11040 974
rect 11000 906 11004 938
rect 11004 906 11036 938
rect 11036 906 11040 938
rect 11000 870 11040 906
rect 11000 838 11004 870
rect 11004 838 11036 870
rect 11036 838 11040 870
rect 11000 802 11040 838
rect 11000 770 11004 802
rect 11004 770 11036 802
rect 11036 770 11040 802
rect 11000 734 11040 770
rect 11000 702 11004 734
rect 11004 702 11036 734
rect 11036 702 11040 734
rect 11000 666 11040 702
rect 11000 634 11004 666
rect 11004 634 11036 666
rect 11036 634 11040 666
rect 11000 598 11040 634
rect 11000 566 11004 598
rect 11004 566 11036 598
rect 11036 566 11040 598
rect 11000 560 11040 566
rect 13250 596 13372 599
rect 13250 564 13275 596
rect 13275 564 13347 596
rect 13347 564 13372 596
rect 13250 559 13372 564
rect 4960 388 4990 414
rect 4990 388 5000 414
rect 5564 388 5570 414
rect 5570 388 5602 414
rect 5602 388 5604 414
rect 6168 388 6182 414
rect 6182 388 6208 414
rect 6772 388 6794 414
rect 6794 388 6812 414
rect 7376 388 7406 414
rect 7406 388 7416 414
rect 7980 388 7982 414
rect 7982 388 8018 414
rect 8018 388 8020 414
rect 8584 388 8594 414
rect 8594 388 8624 414
rect 9188 388 9206 414
rect 9206 388 9228 414
rect 9792 388 9818 414
rect 9818 388 9832 414
rect 10396 388 10398 414
rect 10398 388 10430 414
rect 10430 388 10436 414
rect 11000 388 11010 414
rect 11010 388 11040 414
rect 13250 388 13254 414
rect 13254 388 13286 414
rect 13286 388 13322 414
rect 13322 388 13354 414
rect 13354 388 13372 414
rect 4960 374 5000 388
rect 5564 374 5604 388
rect 6168 374 6208 388
rect 6772 374 6812 388
rect 7376 374 7416 388
rect 7980 374 8020 388
rect 8584 374 8624 388
rect 9188 374 9228 388
rect 9792 374 9832 388
rect 10396 374 10436 388
rect 11000 374 11040 388
rect 13250 374 13372 388
<< metal2 >>
rect 9449 2064 9570 2086
rect 4960 1953 5000 1980
rect 4960 0 5000 27
rect 5056 -96 5146 2064
rect 5221 1420 5343 2064
rect 5221 -96 5343 560
rect 5406 -96 5496 2064
rect 5564 1953 5604 1980
rect 5564 0 5604 27
rect 5656 -96 5746 2064
rect 5825 1420 5947 2064
rect 5825 -96 5947 560
rect 6016 -96 6106 2064
rect 6168 1953 6208 1980
rect 6168 0 6208 27
rect 6266 -96 6356 2064
rect 6429 1420 6551 2064
rect 6429 -96 6551 560
rect 6616 -96 6706 2064
rect 6772 1953 6812 1980
rect 6772 0 6812 27
rect 6866 -96 6956 2064
rect 7033 1420 7155 2064
rect 7033 -96 7155 560
rect 7226 -96 7316 2064
rect 7376 1953 7416 1980
rect 7376 0 7416 27
rect 7476 -96 7566 2064
rect 7637 1420 7759 2064
rect 7637 -96 7759 560
rect 7826 -96 7916 2064
rect 7980 1953 8020 1980
rect 7980 0 8020 27
rect 8076 -96 8166 2064
rect 8241 1420 8363 2064
rect 8241 -96 8363 560
rect 8426 -96 8516 2064
rect 8584 1953 8624 1980
rect 8584 0 8624 27
rect 8676 -96 8766 2064
rect 8845 1420 8967 2064
rect 8845 -96 8967 560
rect 9036 -96 9126 2064
rect 9188 1953 9228 1980
rect 9188 0 9228 27
rect 9286 -96 9376 2064
rect 9440 1702 9578 2064
rect 9449 1420 9571 1702
rect 9449 -96 9571 560
rect 9636 -96 9726 2064
rect 9792 1953 9832 1980
rect 9792 0 9832 27
rect 9886 -96 9976 2064
rect 10053 1420 10175 2064
rect 10053 -96 10175 560
rect 10246 -96 10336 2064
rect 10396 1953 10436 1980
rect 10396 0 10436 27
rect 10496 -96 10586 2064
rect 10656 1980 10776 2074
rect 10656 1420 10779 1980
rect 10656 560 10657 1420
rect 10656 551 10779 560
rect 10656 -96 10776 551
rect 10846 -96 10936 2074
rect 11000 1953 11040 1980
rect 13250 599 13372 609
rect 13250 414 13372 559
rect 13250 365 13372 374
rect 11000 0 11040 27
<< via2 >>
rect 4960 1606 5000 1953
rect 4960 1566 5000 1606
rect 4960 1420 5000 1566
rect 4960 560 5000 1420
rect 4960 414 5000 560
rect 4960 374 5000 414
rect 4960 27 5000 374
rect 5564 1606 5604 1953
rect 5564 1566 5604 1606
rect 5564 1420 5604 1566
rect 5564 560 5604 1420
rect 5564 414 5604 560
rect 5564 374 5604 414
rect 5564 27 5604 374
rect 6168 1606 6208 1953
rect 6168 1566 6208 1606
rect 6168 1420 6208 1566
rect 6168 560 6208 1420
rect 6168 414 6208 560
rect 6168 374 6208 414
rect 6168 27 6208 374
rect 6772 1606 6812 1953
rect 6772 1566 6812 1606
rect 6772 1420 6812 1566
rect 6772 560 6812 1420
rect 6772 414 6812 560
rect 6772 374 6812 414
rect 6772 27 6812 374
rect 7376 1606 7416 1953
rect 7376 1566 7416 1606
rect 7376 1420 7416 1566
rect 7376 560 7416 1420
rect 7376 414 7416 560
rect 7376 374 7416 414
rect 7376 27 7416 374
rect 7980 1606 8020 1953
rect 7980 1566 8020 1606
rect 7980 1420 8020 1566
rect 7980 560 8020 1420
rect 7980 414 8020 560
rect 7980 374 8020 414
rect 7980 27 8020 374
rect 8584 1606 8624 1953
rect 8584 1566 8624 1606
rect 8584 1420 8624 1566
rect 8584 560 8624 1420
rect 8584 414 8624 560
rect 8584 374 8624 414
rect 8584 27 8624 374
rect 9188 1606 9228 1953
rect 9188 1566 9228 1606
rect 9188 1420 9228 1566
rect 9188 560 9228 1420
rect 9188 414 9228 560
rect 9188 374 9228 414
rect 9188 27 9228 374
rect 9792 1606 9832 1953
rect 9792 1566 9832 1606
rect 9792 1420 9832 1566
rect 9792 560 9832 1420
rect 9792 414 9832 560
rect 9792 374 9832 414
rect 9792 27 9832 374
rect 10396 1606 10436 1953
rect 10396 1566 10436 1606
rect 10396 1420 10436 1566
rect 10396 560 10436 1420
rect 10396 414 10436 560
rect 10396 374 10436 414
rect 10396 27 10436 374
rect 11000 1606 11040 1953
rect 11000 1566 11040 1606
rect 11000 1420 11040 1566
rect 11000 560 11040 1420
rect 11000 414 11040 560
rect 11000 374 11040 414
rect 11000 27 11040 374
<< metal3 >>
rect 4960 1953 5000 1962
rect 4960 18 5000 27
rect 5056 -96 5146 2064
rect 5406 -96 5496 2064
rect 5564 1953 5604 1962
rect 5564 18 5604 27
rect 5656 -96 5746 2064
rect 6016 -96 6106 2064
rect 6168 1953 6208 1962
rect 6168 18 6208 27
rect 6266 -96 6356 2064
rect 6616 -96 6706 2064
rect 6772 1953 6812 1962
rect 6772 18 6812 27
rect 6866 -96 6956 2064
rect 7226 -96 7316 2064
rect 7376 1953 7416 1962
rect 7376 18 7416 27
rect 7476 -96 7566 2064
rect 7826 -96 7916 2064
rect 7980 1953 8020 1962
rect 7980 18 8020 27
rect 8076 -96 8166 2064
rect 8426 -96 8516 2064
rect 8584 1953 8624 1962
rect 8584 18 8624 27
rect 8676 -96 8766 2064
rect 9036 -96 9126 2064
rect 9188 1953 9228 1962
rect 9188 18 9228 27
rect 9286 -96 9376 2064
rect 9636 -96 9726 2064
rect 9792 1953 9832 1962
rect 9792 18 9832 27
rect 9886 -96 9976 2064
rect 10246 -96 10336 2064
rect 10396 1953 10436 1962
rect 10396 18 10436 27
rect 10496 -96 10586 2064
rect 10846 -96 10936 2074
rect 11000 1953 11040 1962
rect 11000 18 11040 27
<< labels >>
flabel metal2 s 10657 551 10779 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 10053 551 10175 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 9449 551 9571 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 8845 551 8967 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 8241 551 8363 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 7637 551 7759 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 6429 551 6551 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel metal2 s 7033 551 7155 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
rlabel metal2 s 5221 551 5343 1980 4 pad
port 2 nsew
flabel metal2 s 5825 551 5947 1980 0 FreeSans 800 0 0 0 pad
port 2 nsew
flabel comment s 13311 990 13311 990 0 FreeSans 734 90 0 0 rppd r=1.959k
rlabel comment s 394 404 394 404 4 sub!
flabel metal1 s 12449 370 12548 420 0 FreeSans 51 0 0 0 iovss
port 4 nsew
<< end >>
