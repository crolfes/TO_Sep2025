magic
tech ihp-sg13g2
magscale 1 2
timestamp 1756361942
<< metal1 >>
rect 7400 2740 7740 2800
rect 7400 -3060 7420 2740
rect 7460 -3060 7740 2740
rect 7400 -3080 7740 -3060
<< via1 >>
rect 40 40 80 2720
rect 420 500 560 2360
rect 5400 1720 6420 1940
rect 5400 820 6420 1040
rect 400 400 2600 500
rect 920 -420 6600 -380
rect 420 -2640 560 -700
rect 5400 -1380 6420 -1160
rect 5400 -2280 6420 -2060
rect 7420 -3060 7460 2740
<< metal2 >>
rect -351 2720 200 2800
rect -351 40 40 2720
rect 80 40 200 2720
rect 300 2360 600 2800
rect 6600 2740 7480 2760
rect 6600 2400 7420 2740
rect 300 2300 420 2360
rect 360 500 420 2300
rect 560 600 600 2360
rect 5000 2380 7420 2400
rect 5000 2370 7120 2380
rect 5200 2220 7120 2370
rect 7280 2220 7420 2380
rect 5200 2200 7420 2220
rect 5000 600 5200 2170
rect 5380 1940 6440 1960
rect 5380 1720 5400 1940
rect 6420 1720 6440 1940
rect 5380 1700 6440 1720
rect 5380 1040 6440 1060
rect 5380 820 5400 1040
rect 6420 820 6440 1040
rect 5380 800 6440 820
rect 6600 600 7420 2200
rect 560 500 2700 600
rect 5000 500 7420 600
rect 360 400 400 500
rect 2600 400 2700 500
rect 360 300 2700 400
rect -351 -160 200 40
rect -351 -460 600 -160
rect 2400 -200 2700 300
rect 4991 400 7420 500
rect 4991 291 7100 400
rect 6600 200 7100 291
rect -351 -461 -48 -460
rect 300 -700 600 -460
rect 900 -380 6600 -200
rect 900 -420 920 -380
rect 900 -480 6600 -420
rect 7000 -600 7100 200
rect 6600 -700 7100 -600
rect 300 -760 420 -700
rect 360 -2640 420 -760
rect 560 -2640 600 -700
rect 360 -2680 600 -2640
rect 5000 -800 7100 -700
rect 7200 -800 7420 400
rect 5000 -1000 7420 -800
rect 5000 -2600 5200 -1000
rect 5380 -1160 6440 -1140
rect 5380 -1380 5400 -1160
rect 6420 -1380 6440 -1160
rect 5380 -1400 6440 -1380
rect 5380 -2060 6440 -2040
rect 5380 -2280 5400 -2060
rect 6420 -2280 6440 -2060
rect 5380 -2300 6440 -2280
rect 6600 -2600 7420 -1000
rect 5000 -2800 7420 -2600
rect 6600 -3060 7420 -2800
rect 7460 -3060 7480 2740
rect 6600 -3100 7480 -3060
<< via2 >>
rect 5000 2170 5200 2370
rect 7120 2220 7280 2380
rect 5400 1720 6420 1940
rect 5400 820 6420 1040
rect 7100 -800 7200 400
rect 5400 -1380 6420 -1160
rect 5400 -2280 6420 -2060
<< metal3 >>
rect 4991 2400 7042 2409
rect 7100 2400 7300 2800
rect 4991 2380 7300 2400
rect 4991 2370 7120 2380
rect 4991 2170 5000 2370
rect 5200 2220 7120 2370
rect 7280 2220 7300 2380
rect 5200 2200 7300 2220
rect 5200 2191 7042 2200
rect 5200 2170 5209 2191
rect 4991 509 5209 2170
rect 7500 1960 7700 2800
rect 5380 1940 7700 1960
rect 5380 1720 5400 1940
rect 6420 1720 7700 1940
rect 5380 1700 7700 1720
rect 7500 1060 7700 1700
rect 5380 1040 7700 1060
rect 5380 820 5400 1040
rect 6420 820 7700 1040
rect 5380 800 7700 820
rect 4991 400 7260 509
rect 4991 291 7100 400
rect 7042 -691 7100 291
rect 4891 -800 7100 -691
rect 7200 -800 7260 400
rect 4891 -909 7260 -800
rect 4893 -2692 5108 -909
rect 7500 -1140 7700 800
rect 5380 -1160 7700 -1140
rect 5380 -1380 5400 -1160
rect 6420 -1380 7700 -1160
rect 5380 -1400 7700 -1380
rect 7500 -2040 7700 -1400
rect 5380 -2060 7700 -2040
rect 5380 -2280 5400 -2060
rect 6420 -2280 7700 -2060
rect 5380 -2300 7700 -2280
rect 4893 -2700 7800 -2692
rect 7900 -2700 8100 2800
rect 4893 -2900 8100 -2700
use sg13g2_DCNDiode  sg13g2_DCNDiode_0
timestamp 1756300284
transform 1 0 358 0 1 -2744
box -456 -456 7068 2508
use sg13g2_DCPDiode  sg13g2_DCPDiode_0
timestamp 1756304713
transform 1 0 358 0 1 358
box -358 -358 6970 2410
<< labels >>
rlabel metal2 -200 2800 -200 2800 1 VSS
port 1 n
rlabel metal2 400 2800 400 2800 1 VDD
port 2 n
rlabel metal3 7200 2800 7200 2800 1 guard
port 3 n
rlabel metal3 7600 2800 7600 2800 1 pad
port 4 n
<< end >>
